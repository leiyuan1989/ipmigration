* 
* No part of this file can be released without the consent of SMIC.
*
* Note: SMIC recommends that users set VNTOL=1E-9 at .option for more smooth convergence.
******************************************************************************************
* 0.11um Mixed Signal 1P8M with MIM Salicide 1.2V/3.3V RF SPICE Model (for HSPICE only)  *
******************************************************************************************
*
* Release version    : 1.14
*
* Release date       : 31/03/2016
*
* Simulation tool    : Synopsys Star-HSPICE version H-2013.03
*
*
*  MIM Capacitor   :
*
*        *------------------------------------------------------------------------------------------------------* 
*        | 1fF/um^2 subckt   |  mim1_rf       |  mim1_shield_rf       | mim1_shield_rf_3t                       |
*        *------------------------------------------------------------------------------------------------------*
*        | 1.5fF/um^2 subckt |  mim15_rf      |  mim15_shield_rf      | mim15_rf_3t       | mim15_shield_rf_3t  |
*        *------------------------------------------------------------------------------------------------------*
*        | 2fF/um^2 subckt   |  mim2_rf_2mask |  mim2_shield_rf_2mask | mim2_shield_rf_2mask_3t                 |
*        *------------------------------------------------------------------------------------------------------*
*        | 3fF/um^2 subckt   |  mim3_rf                                                                         |
*        *------------------------------------------------------------------------------------------------------*
*******************************
* 0.11um 1fF/um^2 MIM Capacitor
*******************************
* 1=port1, 2=port2
.subckt mim1_rf 1 2 lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param
*** mismatch paramters
*+sigma_mis_mim_rf    = agauss(0,1,1)
+ac0 = 0.0384    cc0 = 1.2717  
+ar_c0 = 'lr*wr*mr*1e12*0.81'
+geo_fac='1/sqrt(ar_c0)'
+dmim1_mis_rf      = 'ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a = 0.971
+cvc1  = 8.03e-6            cvc2 = 3.74e-6  ctc1 = 4.088E-05 
+c0    = 'c0_a*ar_c0'
+tcoef(temper) = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((0.1709-5.88E-06*lr*wr*1E12*0.81)*1E-9*(0.0095*pwr(lr*wr*0.81,-0.1852)), 1E-13)'
+Cf_rf     = 'c0*1E-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'              
+Rs_rf     = 'max(189.3258/(lr*wr*1E12*0.81)*(0.9985*exp(547415735.7484*lr*wr*0.81)), 1E-6)'
+Rsub1_rf  = 'max(3.0E+04-2.0*lr*wr*1E12*0.81, 1E-3)'
+Csub1_rf  = 'max((0.08*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox1_rf   = 'max((2.5E-03*lr*wr*1E12*0.81)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max(4.88E+03-6.495E-3*lr*wr*1E12*0.81, 1E-3)'
+Csub2_rf  = 'max((0.1*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox2_rf   = 'max((6.38E-03*lr*wr*1E12*0.81)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls     1 11  Ls_rf m=mr
Cf    22  2  'Cf_rf*(1+dmim1_rf)*(1+dmim1_mis_rf)*tcoef(temper)*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))'
Rs    11 22  Rs_rf m=mr
Rsub1 10  0  Rsub1_rf m=mr
Csub1 10  0  Csub1_rf m=mr
Cox1   1 10  Cox1_rf m=mr
Rsub2 20  0  Rsub2_rf m=mr
Csub2 20  0  Csub2_rf m=mr
Cox2   2 20  Cox2_rf m=mr
.ends mim1_rf
**************************************************************
* 0.11um 1fF/um^2 MIM Capacitor with shielding layer
**************************************************************
* 1=port1, 2=port2
.subckt mim1_shield_rf 1 2 lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param
*** mismatch paramters
*+sigma_mis_mim_rf    = agauss(0,1,1)
+ac0 = 0.0384    cc0 = 1.2717  
+ar_c0 = 'lr*wr*mr*1e12*0.81'
+geo_fac='1/sqrt(ar_c0)'
+dmim1_mis_rf      = 'ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a = 0.971
+cvc1  = 8.03e-6            cvc2 = 3.74e-6  ctc1 = 4.088E-05 
+c0    = 'c0_a*ar_c0'
+tcoef(temper) = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((0.1709-5.88E-06*lr*wr*1E12*0.81)*1E-9*(0.0095*pwr(lr*wr*0.81,-0.1852)), 1E-13)'
+Cf_rf     = 'c0*1E-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'              
+Rs_rf     = 'max(189.3258/(lr*wr*1E12*0.81)*(0.9985*exp(547415735.7484*lr*wr*0.81))*(1.9845*pwr(lr*wr*0.81,0.02675)), 1E-6)'
+Rsub1_rf  = 'max(3.0E+04-2.0*lr*wr*1E12*0.81, 1E-3)'
+Csub1_rf  = 'max((0.08*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox1_rf   = 'max((2.5E-03*lr*wr*1E12*0.81)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max((4.88E+03-6.495E-3*lr*wr*1E12*0.81)/(875777*pwr(lr*wr*0.81,0.38965)), 1E-3)'
+Csub2_rf  = 'max((0.1*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox2_rf   = 'max((6.38E-03*lr*wr*1E12*0.81)*1E-15+(0.08505*lr*wr*1e12+0.9)*1e-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls     1 11  Ls_rf m=mr
Cf    22  2  'Cf_rf*(1+dmim1_shield_rf)*(1+dmim1_mis_rf)*tcoef(temper)*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))'
Rs    11 22  Rs_rf m=mr
Rsub1 10  0  Rsub1_rf m=mr
Csub1 10  0  Csub1_rf m=mr
Cox1   1 10  Cox1_rf m=mr
Rsub2 20  0  Rsub2_rf m=mr
Csub2 20  0  Csub2_rf m=mr
Cox2   2 20  Cox2_rf m=mr
.ends mim1_shield_rf
**************************************************************
* 0.11um 1fF/um^2 MIM Capacitor with shielding layer (3-terminal)
**************************************************************
* 1=port1, 2=port2
.subckt mim1_shield_rf_3t 1 2 p lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param
*** mismatch paramters
*+sigma_mis_mim_rf    = agauss(0,1,1)
+ac0 = 0.0384    cc0 = 1.2717  
+ar_c0 = 'lr*wr*mr*1e12*0.81'
+geo_fac='1/sqrt(ar_c0)'
+dmim1_mis_rf      = 'ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a = 0.971
+cvc1  = 8.03e-6            cvc2 = 3.74e-6  ctc1 = 4.088E-05 
+c0    = 'c0_a*ar_c0'
+tcoef(temper) = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((0.1709-5.88E-06*lr*wr*1E12*0.81)*1E-9*(0.0095*pwr(lr*wr*0.81,-0.1852)), 1E-13)'
+Cf_rf     = 'c0*1E-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'              
+Rs_rf     = 'max(189.3258/(lr*wr*1E12*0.81)*(0.9985*exp(547415735.7484*lr*wr*0.81))*(1.9845*pwr(lr*wr*0.81,0.02675)), 1E-6)'
+Rsub1_rf  = 'max(3.0E+04-2.0*lr*wr*1E12*0.81, 1E-3)'
+Csub1_rf  = 'max((0.08*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox1_rf   = 'max((2.5E-03*lr*wr*1E12*0.81)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max((4.88E+03-6.495E-3*lr*wr*1E12*0.81)/(875777*pwr(lr*wr*0.81,0.38965)), 1E-3)'
+Csub2_rf  = 'max((0.1*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox2_rf   = 'max((6.38E-03*lr*wr*1E12*0.81)*1E-15+(0.08505*lr*wr*1e12+0.9)*1e-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls     1 11  Ls_rf m=mr
Cf    22  2  'Cf_rf*(1+dmim1_shield_rf)*(1+dmim1_mis_rf)*tcoef(temper)*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))'
Rs    11 22  Rs_rf m=mr
Rsub1 10  p  Rsub1_rf m=mr
Csub1 10  p  Csub1_rf m=mr
Cox1   1 10  Cox1_rf m=mr
Rsub2 20  p  Rsub2_rf m=mr
Csub2 20  p  Csub2_rf m=mr
Cox2   2 20  Cox2_rf m=mr
.ends mim1_shield_rf_3t
*********************************
* 0.11um 1.5fF/um^2 MIM Capacitor
*********************************
* 1=port1, 2=port2
.subckt mim15_rf 1 2 lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param
*** mismatch paramters  
*+sigma_mis_mim_rf    = agauss(0,1,1)
+ac0 = 2.2793E-02    cc0 = 1.1757 
+ar_c0 = 'lr*wr*mr*1e12*0.81'
+geo_fac='1/sqrt(ar_c0)'
+dmim15_mis_rf      = 'ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a      = 1.449      ctc1 = 3.758E-05       
+cvc1      = 9.68e-6                    cvc2 = 6.72e-6          
+c0        = 'c0_a*ar_c0'
+tcoef     = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((0.1709-5.88E-06*lr*wr*1E12*0.81)*1E-9, 1E-13)'
+Cf_rf     = 'c0*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'
+Rs_rf     = 'max(189.3258/(lr*wr*1E12*0.81), 1E-6)'
+Rsub1_rf  = 'max(3.0E+04-2.0*lr*wr*1E12*0.81, 1E-3)'
+Csub1_rf  = 'max((0.08*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox1_rf   = 'max((0.08*pwr(wr*lr*0.81*1e12,0.5)+0.02)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max(4.88E+03-6.495E-3*lr*wr*1E12*0.81, 1E-3)'
+Csub2_rf  = 'max((0.1*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox2_rf   = 'max((0.2*pwr(wr*lr*0.81*1e12,0.5)+0.46)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls     1 11  Ls_rf m=mr
Cf    22  2  'Cf_rf*(1+dmim15_rf)*(1+dmim15_mis_rf)*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))'
Rs    11 22  Rs_rf m=mr
Rsub1 10  0  Rsub1_rf  m=mr
Csub1 10  0  Csub1_rf m=mr
Cox1   1 10  Cox1_rf   m=mr
Rsub2 20  0  Rsub2_rf  m=mr
Csub2 20  0  Csub2_rf  m=mr
Cox2   2 20  Cox2_rf m=mr
.ends mim15_rf
****************************************************
* 0.11um 1.5fF/um^2 MIM Capacitor (3-terminal)
****************************************************
* 1=port1, 2=port2
.subckt mim15_rf_3t 1 2 p lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param
*** mismatch paramters  
*+sigma_mis_mim_rf    = agauss(0,1,1)
+ac0 = 2.2793E-02    cc0 = 1.1757 
+ar_c0 = 'lr*wr*mr*1e12*0.81'
+geo_fac='1/sqrt(ar_c0)'
+dmim15_mis_rf      = 'ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a      = 1.449      ctc1 = 3.758E-05       
+cvc1      = 9.68e-6                    cvc2 = 6.72e-6          
+c0        = 'c0_a*ar_c0'
+tcoef     = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((0.1709-5.88E-06*lr*wr*1E12*0.81)*1E-9, 1E-13)'
+Cf_rf     = 'c0*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'
+Rs_rf     = 'max(189.3258/(lr*wr*1E12*0.81), 1E-6)'
+Rsub1_rf  = 'max(3.0E+04-2.0*lr*wr*1E12*0.81, 1E-3)'
+Csub1_rf  = 'max((0.08*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox1_rf   = 'max((0.08*pwr(wr*lr*0.81*1e12,0.5)+0.02)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'
+Rsub2_rf  = 'max(4.88E+03-6.495E-3*lr*wr*1E12*0.81, 1E-3)'
+Csub2_rf  = 'max((0.1*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox2_rf   = 'max((0.2*pwr(wr*lr*0.81*1e12,0.5)+0.46)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls     1 11  Ls_rf m=mr
Cf    22  2  'Cf_rf*(1+dmim15_rf)*(1+dmim15_mis_rf)*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))'
Rs    11 22  Rs_rf m=mr
Rsub1 10  p  Rsub1_rf m=mr
Csub1 10  p  Csub1_rf m=mr
Cox1   1 10  Cox1_rf m=mr
Rsub2 20  p  Rsub2_rf m=mr
Csub2 20  p  Csub2_rf m=mr
Cox2   2 20  Cox2_rf m=mr
.ends mim15_rf_3t
**************************************************************
* 0.11um 1.5fF/um^2 MIM Capacitor with shielding layer
**************************************************************
* 1=port1, 2=port2
.subckt mim15_shield_rf 1 2 lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param
*** mismatch paramters  
*+sigma_mis_mim_rf    = agauss(0,1,1)
+ac0 = 2.2793E-02    cc0 = 1.1757 
+ar_c0 = 'lr*wr*mr*1e12*0.81' 
+geo_fac='1/sqrt(ar_c0)'
+dmim15_mis_rf      = 'ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a      = 1.449      ctc1 = 3.758E-05       
+cvc1      = 9.68e-6                    cvc2 = 6.72e-6          
+c0        = 'c0_a*ar_c0'
+tcoef     = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((0.1709-5.88E-06*lr*wr*1E12*0.81)*1E-9, 1E-13)'
+Cf_rf     = 'c0*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'              
+Rs_rf     = 'max(189.3258/(lr*wr*1E12*0.81)*(1.9845*pwr(lr*wr*0.81,0.02675)), 1E-6)'
+Rsub1_rf  = 'max(3.0E+04-2.0*lr*wr*1E12*0.81, 1E-3)'
+Csub1_rf  = 'max((0.08*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox1_rf   = 'max((0.08*pwr(wr*lr*0.81*1e12,0.5)+0.02)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max((4.88E+03-6.495E-3*lr*wr*1E12*0.81)/(613044*pwr(lr*wr*0.81,0.38965)), 1E-3)'
+Csub2_rf  = 'max((0.1*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox2_rf   = 'max((6.38E-03*lr*wr*1E12*0.81)*1E-15+(0.08505*lr*wr*1e12+0.9)*1e-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls     1 11  Ls_rf m=mr
Cf    22  2  'Cf_rf*(1+dmim15_shield_rf)*(1+dmim15_mis_rf)*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))'
Rs    11 22  Rs_rf m=mr
Rsub1 10  0  Rsub1_rf m=mr
Csub1 10  0  Csub1_rf m=mr
Cox1   1 10  Cox1_rf m=mr
Rsub2 20  0  Rsub2_rf m=mr
Csub2 20  0  Csub2_rf m=mr
Cox2   2 20  Cox2_rf m=mr
.ends mim15_shield_rf m=mr
***************************************************************************
* 0.11um 1.5fF/um^2 MIM Capacitor with shielding layer (3-terminal)
***************************************************************************
* 1=port1, 2=port2
.subckt mim15_shield_rf_3t 1 2 p lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param
*** mismatch paramters  
*+sigma_mis_mim_rf    = agauss(0,1,1)
+ac0 = 2.2793E-02    cc0 = 1.1757 
+ar_c0 = 'lr*wr*mr*1e12*0.81' 
+geo_fac='1/sqrt(ar_c0)'
+dmim15_mis_rf      = 'ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a      = 1.449      ctc1 = 3.758E-05       
+cvc1      = 9.68e-6                    cvc2 = 6.72e-6          
+c0        = 'c0_a*ar_c0'
+tcoef     = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((0.1709-5.88E-06*lr*wr*1E12*0.81)*1E-9, 1E-13)'
+Cf_rf     = 'c0*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'              
+Rs_rf     = 'max(189.3258/(lr*wr*1E12*0.81)*(1.9845*pwr(lr*wr*0.81,0.02675)), 1E-6)'
+Rsub1_rf  = 'max(3.0E+04-2.0*lr*wr*1E12*0.81, 1E-3)'
+Csub1_rf  = 'max((0.08*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox1_rf   = 'max((0.08*pwr(wr*lr*0.81*1e12,0.5)+0.02)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max((4.88E+03-6.495E-3*lr*wr*1E12*0.81)/(613044*pwr(lr*wr*0.81,0.38965)), 1E-3)'
+Csub2_rf  = 'max((0.1*lr*1E6*0.9)*1E-15, 1E-18)'  
+Cox2_rf   = 'max((6.38E-03*lr*wr*1E12*0.81)*1E-15+(0.08505*lr*wr*1e12+0.9)*1e-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls     1 11  Ls_rf m=mr
Cf    22  2  'Cf_rf*(1+dmim15_shield_rf)*(1+dmim15_mis_rf)*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))'
Rs    11 22  Rs_rf m=mr
Rsub1 10  p  Rsub1_rf m=mr
Csub1 10  p  Csub1_rf m=mr
Cox1   1 10  Cox1_rf m=mr
Rsub2 20  p  Rsub2_rf m=mr
Csub2 20  p  Csub2_rf m=mr
Cox2   2 20  Cox2_rf m=mr
.ends mim15_shield_rf_3t 
*******************************
* 0.11um 2fF/um^2 MIM Capacitor
*******************************
* 1=port1, 2=port2
.subckt mim2_rf_2mask 1 2 lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param 
*** mismatch paramters
+ac0 = 0.132900035    cc0 = 0.000206611
*+sigma_mis_mim_rf    = agauss(0,1,1)
+dmim2_2mask_mis_rf = '(ac0/c0+cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a = 2.1 
+cvc1 = -6.119607E-05 cvc2 = 2.660293E-05  ctc1 = 3.25876E-05  
+ar_c0 = 'lr*wr*mr*1e12*0.81'  
+c0    = 'c0_a*ar_c0'
+tcoef = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((2.09*pwr(lr*wr*1e12*0.81,-1.35)+4.1e-6*lr*wr*1e12*0.81+0.0061)*1e-9,1e-15)'
+Cf_rf     = 'c0*(1+DMIM2_RF_2mask)*(1+dmim2_2mask_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'              
+Rs_rf     = 'max(43.7*pwr(lr*wr*1e12*0.81,-0.83)+0.00035*lr*wr*1e12*0.81,1e-6)'
+Rsub1_rf  = 'max(31950*pwr(lr*wr*1e12*0.81,-0.021), 1E-3)'
+Csub1_rf  = 'max((0.08*sqrt(lr*wr*1e12*0.81))*1E-15, 1E-18)'  
+Cox1_rf   = 'max((2.5E-03*lr*wr*1e12*0.81)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max(4929.7*pwr(lr*wr*1e12*0.81,-0.0946), 1E-3)'
+Csub2_rf  = 'max((0.1*sqrt(lr*wr*1e12*0.81))*1E-15, 1E-18)'  
+Cox2_rf   = 'max((6.38E-03*lr*wr*1e12*0.81)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls 1 11    Ls_rf m=mr
Cf 22 2    'Cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))'                                       
Rs 11 22   Rs_rf m=mr
Rsub1 10 0 Rsub1_rf m=mr
Csub1 10 0 Csub1_rf m=mr
Cox1 1 10  Cox1_rf m=mr
Rsub2 20 0 Rsub2_rf m=mr
Csub2 20 0 Csub2_rf m=mr
Cox2 2 20  Cox2_rf m=mr
.ends mim2_rf_2mask
****************************************************
* 0.11um 2fF/um^2 MIM Capacitor with shielding layer 
****************************************************
* 1=port1, 2=port2
.subckt mim2_shield_rf_2mask 1 2 lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param 
*** mismatch paramters
+ac0 = 0.132900035    cc0 = 0.000206611
*+sigma_mis_mim_rf    = agauss(0,1,1)
+dmim2_2mask_mis_rf = '(ac0/c0+cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a = 2.1 
+cvc1 = -6.119607E-05 cvc2 = 2.660293E-05  ctc1 = 3.25876E-05  
+ar_c0 = 'lr*wr*mr*1e12*0.81'  
+c0    = 'c0_a*ar_c0'
+tcoef = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((1.23*pwr(lr*wr*1e12*0.81,-1.25)+4.1e-6*lr*wr*1e12*0.81+0.0061)*1e-9,1e-15)'
+Cf_rf     = 'c0*(1+DMIM2_shield_RF_2mask)*(1+dmim2_2mask_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'              
+Rs_rf     = 'max(43.7*pwr(lr*wr*1e12*0.81,-0.83)+0.00019*lr*wr*1e12*0.81,1e-6)'
+Rsub1_rf  = 'max(31950*pwr(lr*wr*1e12*0.81,-0.021), 1E-3)'
+Csub1_rf  = 'max((0.08*sqrt(lr*wr*1e12*0.81))*1E-15, 1E-18)'  
+Cox1_rf   = 'max((2.5E-03*lr*wr*1e12*0.81)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max(19.557*pwr(lr*wr*1e12*0.81,-0.3473), 1E-3)'
+Csub2_rf  = 'max((0.1*sqrt(lr*wr*1e12*0.81))*1E-15, 1E-18)'  
+Cox2_rf   = 'max((2.9453*pwr(lr*wr*1e12*0.81,0.87)+20.224)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls 1 11    Ls_rf m=mr
Cf 22 2    'Cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))' 
Rs 11 22   Rs_rf    m=mr
Rsub1 10 0 Rsub1_rf m=mr
Csub1 10 0 Csub1_rf m=mr
Cox1 1 10  Cox1_rf m=mr
Rsub2 20 0 Rsub2_rf m=mr
Csub2 20 0 Csub2_rf m=mr
Cox2 2 20  Cox2_rf m=mr
.ends mim2_shield_rf_2mask
****************************************************
* 0.11um 2fF/um^2 MIM Capacitor with shielding layer (3-terminal)
****************************************************
* 1=port1, 2=port2
.subckt mim2_shield_rf_2mask_3t 1 2 p lr=l wr=w mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param 
*** mismatch paramters
+ac0 = 0.132900035    cc0 = 0.000206611
*+sigma_mis_mim_rf    = agauss(0,1,1)
+dmim2_2mask_mis_rf = '(ac0/c0+cc0)*sigma_mis_mim_rf*mismod_mim_rf'
***
+c0_a = 2.1 
+cvc1 = -6.119607E-05 cvc2 = 2.660293E-05  ctc1 = 3.25876E-05  
+ar_c0 = 'lr*wr*mr*1e12*0.81'  
+c0    = 'c0_a*ar_c0'
+tcoef = '1.0+ctc1*(temper-25.0)'
+Ls_rf     = 'max((1.23*pwr(lr*wr*1e12*0.81,-1.25)+4.1e-6*lr*wr*1e12*0.81+0.0061)*1e-9,1e-15)'
+Cf_rf     = 'c0*(1+DMIM2_shield_RF_2mask)*(1+dmim2_2mask_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))'              
+Rs_rf     = 'max(43.7*pwr(lr*wr*1e12*0.81,-0.83)+0.00019*lr*wr*1e12*0.81,1e-6)'
+Rsub1_rf  = 'max(31950*pwr(lr*wr*1e12*0.81,-0.021), 1E-3)'
+Csub1_rf  = 'max((0.08*sqrt(lr*wr*1e12*0.81))*1E-15, 1E-18)'  
+Cox1_rf   = 'max((2.5E-03*lr*wr*1e12*0.81)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max(19.557*pwr(lr*wr*1e12*0.81,-0.3473), 1E-3)'
+Csub2_rf  = 'max((0.1*sqrt(lr*wr*1e12*0.81))*1E-15, 1E-18)'  
+Cox2_rf   = 'max((2.9453*pwr(lr*wr*1e12*0.81,0.87)+20.224)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)'
* equivalent circuit
Ls 1 11    Ls_rf m=mr
Cf 22 2    'Cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))' 
Rs 11 22   Rs_rf    m=mr
Rsub1 10 p Rsub1_rf m=mr
Csub1 10 p Csub1_rf m=mr
Cox1 1 10  Cox1_rf m=mr
Rsub2 20 p Rsub2_rf m=mr
Csub2 20 p Csub2_rf m=mr
Cox2 2 20  Cox2_rf m=mr
.ends mim2_shield_rf_2mask_3t
****************************************************
* 0.11um 3fF/um^2 stacked MIM Capacitor 
****************************************************
.subckt mim3_rf 1 2 wr=w lr=l mr=m mismod_mim_rf=0 xm=8
* mim capacitor scalable model parameters
.param
*** mismatch paramters
*+sigma_mis_mim_rf    = agauss(0,1,1)
+ac0 = 0.3305    cc0 = 0.000152
+dmim3_mis_rf      = '(ac0/c0+cc0)*sigma_mis_mim_rf*mismod_mim_rf'
*** low frequency capacitor    
+c0_a = 3.01368807   c0_p = 0.44926463
+cvc1 = 2.37303251E-06  cvc2 = 8.08656805E-06  ctc1 = 3.92547475E-05  ctc2=1.26746609E-07
*
+ar_c0 = 'lr*wr*mr*1e12*0.81'  
+pe_c0 = '2*(lr+wr)*mr*1e6*0.9' 
+c0    = 'c0_a*ar_c0+c0_p*pe_c0'
+tcoef(temper) = '1.0+ctc1*(temper-25.0)+ctc2*(temper-25.0)*(temper-25.0)'
***
+Ls_rf     = 'max((1.13*pwr(lr*wr*1e12*0.81,-1.4)+0.005)*1E-9, 1E-12)'
+Cf_rf     = 'max(c0*(1+dmim3_rf)*(1+dmim3_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8))),1e-18)'
+Rs_rf     = 'max(65*pwr(lr*wr*1e12*0.81,-1)+0.53, 1E-6)'
+Rsub1_rf  = 'max(1887.8*pwr(lr*wr*1e12*0.81,-0.3764), 1E-3)'
+Csub1_rf  = 'max(73.335*pwr(lr*wr*1e12*0.81,-0.6825)*1E-15, 1E-18)'  
+Cox1_rf   = 'max((0.0172*lr*wr*1e12*0.81+0.2275)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)'            
+Rsub2_rf  = 'max(1000, 1E-3)'
+Csub2_rf  = 'max(1*1E-15, 1E-18)'  
+Cox2_rf   = 'max(0.0098*2*(lr+wr)*1E6*0.9*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)' 
* equivalent circuit
Ls 1 11    Ls_rf m=mr
*Cf 22 2    'Cf_rf*tcoef(temper)*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))'
Cf 22 2    'c0*1e-15'
Rs 11 22   Rs_rf m=mr
Rsub1 10 0 Rsub1_rf m=mr
Csub1 10 0 Csub1_rf m=mr
Cox1 1 10  Cox1_rf m=mr
Rsub2 20 0 Rsub2_rf m=mr
Csub2 20 0 Csub2_rf m=mr
Cox2 2 20  Cox2_rf m=mr
.ends mim3_rf
