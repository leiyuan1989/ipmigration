* 
* No part of this file can be released without the consent of SMIC.
*
************************************************************************************************************
* SMIC 0.11um Mixed Signal 1P6M(1P5M, 1P7M, 1P8M) 1.2V/3.3V SPICE model (for HSPICE only) * 
************************************************************************************************************
*
* Release version    : 1.14
*
* Release date       : 03/28/2016
*
* Simulation tool    : Synopsys Star-HSPICE version I-2013.12
*
*  Inductor   :
* *  *------------------------*-----------------------------------------------------------------------------------------------------*
*    |  Turn, Radius & Width  |T=1~3 step 0.5,W=5~13.5um,R=1.7071*W+16.378~120um;T=3.5~5.0 step 0.5,W=5~8um,R=1.7071*W+16.378~120um |
* *  *------------------------*-----------------------------------------------------------------------------------------------------*
*    |        Model Name      |     diff_ind_3t_rf_pgs_psub_n                             							|   
* *  *------------------------*-----------------------------------------------------------------------------------------------------*
.subckt diff_ind_3t_rf_pgs_psub_n PLUS MINUS CT PSUB r=6e-05 w=8e-06 n=3
.param radius_='0.00833333*(r/1e-06-0)' w_='0.0666667*(w/1e-06-0)'
.param T51='(1-abs(sgn(n-(1.5))))'
.param T52='(min(sgn(radius_-(0.416958))+1,1))'
.param T53='(min(sgn(w_+7.291667e-01*radius_-(0.904432))+1,1))'
.param T54='(min(sgn(w_-(0.6004))+1,1))'
.param T55='(min(sgn(radius_-(0.416375))+1,1))'
.param T56='(min(sgn(radius_-(0.708625))+1,1))'
.param T57='(min(sgn(w_+7.291667e-01*radius_-(0.903207))+1,1))'
.param T58='(min(sgn(w_-(0.5996))+1,1))'
.param T59='(min(sgn(radius_-(0.708042))+1,1))'
.param T60='(1-abs(sgn(n-(1))))'
.param T61='(1-abs(sgn(n-(2.5))))'
.param T62='(1-abs(sgn(n-(2))))'
.param T63='(1-abs(sgn(n-(3.5))))'
.param T64='(1-abs(sgn(n-(3))))'
.param T65='(1-abs(sgn(n-(4.5))))'
.param T66='(1-abs(sgn(n-(4))))'
.param T67='(1-abs(sgn(n-(5))))'
.param S0='T51*(1-T52)*(1-T53)'
.param noS0='(1-S0)'
.param S1='T51*(1-T54)*T55*(1-T56)*noS0'
.param noS1='(1-S1)*noS0'
.param S2='T51*T57*T58*(1-T56)*noS1'
.param noS2='(1-S2)*noS1'
.param S3='T51*(1-T54)*T59*noS2'
.param noS3='(1-S3)*noS2'
.param S4='T51*T59*T58*noS3'
.param noS4='(1-S4)*noS3'
.param S5='T60*(1-T52)*(1-T53)*noS4'
.param noS5='(1-S5)*noS4'
.param S6='T60*(1-T54)*T55*(1-T56)*noS5'
.param noS6='(1-S6)*noS5'
.param S7='T60*T57*T58*(1-T56)*noS6'
.param noS7='(1-S7)*noS6'
.param S8='T60*(1-T54)*T59*noS7'
.param noS8='(1-S8)*noS7'
.param S9='T60*T59*T58*noS8'
.param noS9='(1-S9)*noS8'
.param S10='T61*(1-T52)*(1-T53)*noS9'
.param noS10='(1-S10)*noS9'
.param S11='T61*(1-T54)*T55*(1-T56)*noS10'
.param noS11='(1-S11)*noS10'
.param S12='T61*T57*T58*(1-T56)*noS11'
.param noS12='(1-S12)*noS11'
.param S13='T61*(1-T54)*T59*noS12'
.param noS13='(1-S13)*noS12'
.param S14='T61*T59*T58*noS13'
.param noS14='(1-S14)*noS13'
.param S15='T62*(1-T52)*(1-T53)*noS14'
.param noS15='(1-S15)*noS14'
.param S16='T62*(1-T54)*T55*(1-T56)*noS15'
.param noS16='(1-S16)*noS15'
.param S17='T62*T57*T58*(1-T56)*noS16'
.param noS17='(1-S17)*noS16'
.param S18='T62*(1-T54)*T59*noS17'
.param noS18='(1-S18)*noS17'
.param S19='T62*T59*T58*noS18'
.param noS19='(1-S19)*noS18'
.param S20='T63*(1-T52)*noS19'
.param noS20='(1-S20)*noS19'
.param S21='T63*T55*(1-T56)*noS20'
.param noS21='(1-S21)*noS20'
.param S22='T63*T59*noS21'
.param noS22='(1-S22)*noS21'
.param S23='T64*(1-T52)*(1-T53)*noS22'
.param noS23='(1-S23)*noS22'
.param S24='T64*(1-T54)*T55*(1-T56)*noS23'
.param noS24='(1-S24)*noS23'
.param S25='T64*T57*T58*(1-T56)*noS24'
.param noS25='(1-S25)*noS24'
.param S26='T64*(1-T54)*T59*noS25'
.param noS26='(1-S26)*noS25'
.param S27='T64*T59*T58*noS26'
.param noS27='(1-S27)*noS26'
.param S28='T65*(1-T52)*noS27'
.param noS28='(1-S28)*noS27'
.param S29='T65*T55*(1-T56)*noS28'
.param noS29='(1-S29)*noS28'
.param S30='T65*T59*noS29'
.param noS30='(1-S30)*noS29'
.param S31='T66*(1-T52)*noS30'
.param noS31='(1-S31)*noS30'
.param S32='T66*T55*(1-T56)*noS31'
.param noS32='(1-S32)*noS31'
.param S33='T66*T59*noS32'
.param noS33='(1-S33)*noS32'
.param S34='T67*(1-T52)*noS33'
.param noS34='(1-S34)*noS33'
.param S35='T67*T55*(1-T56)*noS34'
.param noS35='(1-S35)*noS34'
.param S36='T67*T59*noS35'
.param noS36='(1-S36)*noS35'
.param V0_part1='3.492189e+01*S0+1.498634e+01*S1+7.682315e-03*S2+(-1.481196e+00)*S3+2.424670e-02*S4+(-1.024208e-02)*S5+(-1.049143e-02)*S6+2.511711e-03*S7+1.801603e-02*S8+(-1.952706e-02)*S9'
.param V0_part2='V0_part1+(-2.620626e-01)*S10+(-2.422198e-02)*S11+7.593669e-03*S12+2.439187e-02*S13+7.290052e-03*S14+(-1.043667e-02)*S15+(-1.866355e-02)*S16+3.350052e-02*S17+(-8.080399e-03)*S18+1.835389e-01*S19'
.param V0_part3='V0_part2+2.181355e+00*S20+(-3.940592e-01)*S21+2.601884e+01*S22+1.957269e+00*S23+1.061720e-02*S24+4.349154e-02*S25+7.125702e-02*S26+1.894228e-02*S27+(-2.993132e-02)*S28+6.788739e+00*S29'
.param V0='V0_part3+(-4.252155e-02)*S30+5.791451e-01*S31+(-5.808421e-02)*S32+(-8.848007e-02)*S33+4.862153e-01*S34+(-4.010336e-01)*S35+2.682741e-02*S36'
.param V1_part1='4.283626e+01*S0+1.581738e+02*S1+4.399911e-01*S2+1.733295e+02*S3+4.685443e-01*S4+3.302335e-01*S5+3.092447e-01*S6+2.912526e-01*S7+2.989596e-01*S8+2.274747e-01*S9'
.param V1_part2='V1_part1+6.010528e+01*S10+1.106671e+00*S11+9.335041e-01*S12+1.091900e+00*S13+1.045815e+00*S14+6.027723e-01*S15+6.623428e-01*S16+2.667990e+01*S17+6.873701e-01*S18+9.337371e+01*S19'
.param V1_part3='V1_part2+1.050482e+02*S20+1.182353e+02*S21+3.403802e+02*S22+6.107540e+01*S23+1.271372e+00*S24+1.128561e+00*S25+1.353456e+00*S26+1.274330e+00*S27+2.585359e+00*S28+1.928785e+02*S29'
.param V1='V1_part3+3.053140e+00*S30+1.556151e+02*S31+2.218325e+00*S32+2.407477e+00*S33+1.370795e+02*S34+2.398841e+02*S35+3.480377e+00*S36'
.param V2_part1='4.801245e+01*S0+1.638839e+02*S1+(-3.672766e-02)*S2+(-1.554958e+01)*S3+(-8.261173e-02)*S4+(-1.818375e-02)*S5+(-3.250482e-02)*S6+(-1.984307e-02)*S7+(-6.211951e-02)*S8+(-1.346350e-02)*S9'
.param V2_part2='V2_part1+(-9.825263e+00)*S10+(-8.918201e-02)*S11+(-2.160178e-02)*S12+(-1.702241e-01)*S13+(-1.249757e-01)*S14+(-3.073835e-02)*S15+(-6.514747e-02)*S16+(-1.728750e+00)*S17+(-1.401968e-01)*S18+(-1.095303e+01)*S19'
.param V2_part3='V2_part2+(-3.354981e+01)*S20+(-8.227739e+00)*S21+(-3.513983e+02)*S22+(-1.996565e+01)*S23+(-1.396479e-01)*S24+(-4.679902e-02)*S25+(-2.222580e-01)*S26+(-1.557216e-01)*S27+1.411389e-01*S28+(-7.697922e+01)*S29'
.param V2='V2_part3+(-3.763692e-01)*S30+(-4.505495e+01)*S31+(-9.589477e-02)*S32+(-3.125850e-01)*S33+(-3.834353e+01)*S34+(-5.490739e+01)*S35+(-5.795492e-01)*S36'
.param V3_part1='2.327377e+03*S0+1.000000e+04*S1+(-8.559012e-02)*S2+2.138974e+03*S3+(-1.855182e-01)*S4+(-1.289876e-01)*S5+(-3.091244e-01)*S6+(-7.619948e-02)*S7+(-3.131067e-01)*S8+(-1.445760e-01)*S9'
.param V3_part2='V3_part1+(-8.494814e+00)*S10+(-3.495595e-01)*S11+(-1.342189e-01)*S12+(-6.170792e-01)*S13+(-3.035582e-01)*S14+(-1.321953e-01)*S15+(-2.746532e-01)*S16+8.067932e+01*S17+(-4.673918e-01)*S18+1.562098e+02*S19'
.param V3_part3='V3_part2+(-1.023105e+03)*S20+2.507655e+02*S21+(-5.808970e+03)*S22+(-6.904830e+02)*S23+(-4.151939e-01)*S24+(-1.120239e-01)*S25+(-6.504459e-01)*S26+(-3.431432e-01)*S27+(-2.196918e-01)*S28+(-1.278556e+03)*S29'
.param V3='V3_part3+(-1.264217e+00)*S30+(-1.295981e+03)*S31+(-6.065976e-01)*S32+(-1.149697e+00)*S33+(-1.093782e+03)*S34+(-8.594428e+02)*S35+(-1.325990e+00)*S36'
.param V4_part1='2.375940e+03*S0+5.909311e+02*S1+3.353615e-01*S2+(-1.833309e+02)*S3+3.199457e-01*S4+1.764118e-01*S5+1.587815e+00*S6+2.167554e-01*S7+(-7.186602e-01)*S8+2.251099e-01*S9'
.param V4_part2='V4_part1+7.557774e+02*S10+9.594171e-01*S11+5.414884e-01*S12+9.505521e-01*S13+5.400986e-01*S14+7.575932e-01*S15+7.010288e-01*S16+5.101988e+01*S17+6.924701e-01*S18+1.395495e+02*S19'
.param V4_part3='V4_part2+2.156607e+03*S20+4.637788e+02*S21+4.327634e+03*S22+1.179979e+03*S23+1.089390e+00*S24+5.673073e-01*S25+1.037683e+00*S26+6.219731e-01*S27+1.881512e+00*S28+1.831622e+03*S29'
.param V4='V4_part3+1.888878e+00*S30+2.748083e+03*S31+1.597399e+00*S32+1.696741e+00*S33+2.304682e+03*S34+1.732534e+03*S35+2.015920e+00*S36'
.param V5_part1='3.532870e+02*S0+2.057697e+02*S1+1.491421e-01*S2+1.666441e+03*S3+2.366327e-01*S4+1.802261e-01*S5+3.555697e-02*S6+7.885749e-02*S7+1.126420e+00*S8+1.297746e-01*S9'
.param V5_part2='V5_part1+1.872154e+02*S10+2.732231e-01*S11+2.661071e-01*S12+4.029103e-01*S13+4.032899e-01*S14+1.180434e-01*S15+1.957133e-01*S16+1.204702e+02*S17+2.943498e-01*S18+6.277762e+02*S19'
.param V5_part3='V5_part2+4.313371e+02*S20+3.863492e+02*S21+2.225099e+03*S22+3.414972e+02*S23+3.174280e-01*S24+2.885576e-01*S25+4.528886e-01*S26+4.541426e-01*S27+3.234155e-01*S28+8.030358e+02*S29'
.param V5='V5_part3+7.781171e-01*S30+5.463263e+02*S31+4.434254e-01*S32+6.490428e-01*S33+4.652185e+02*S34+7.853602e+02*S35+8.367272e-01*S36'
.param V6_part1='1.483120e+01*S0+2.672647e+01*S1+7.319749e-03*S2+1.699497e+00*S3+(-2.240943e-02)*S4+1.732036e-02*S5+8.606841e-02*S6+0.000000e+00*S7+2.746039e-01*S8+2.930952e-02*S9'
.param V6_part2='V6_part1+6.196135e-01*S10+0.000000e+00*S11+(-2.581440e-02)*S12+(-7.259091e-02)*S13+(-1.941969e-02)*S14+0.000000e+00*S15+0.000000e+00*S16+5.102252e-01*S17+(-3.596031e-02)*S18+6.202202e+00*S19'
.param V6_part3='V6_part2+1.249121e+00*S20+(-1.260548e+00)*S21+(-1.393818e+01)*S22+3.428114e+00*S23+(-2.603205e-02)*S24+(-3.715578e-02)*S25+(-1.115860e-01)*S26+(-1.596824e-02)*S27+0.000000e+00*S28+3.784328e+00*S29'
.param V6='V6_part3+(-6.901881e-02)*S30+2.992865e+00*S31+0.000000e+00*S32+(-1.244395e-02)*S33+3.787482e+00*S34+1.282741e+01*S35+(-1.155982e-01)*S36'
.param V7_part1='9.257384e+00*S0+7.383394e+01*S1+2.974102e-02*S2+4.001306e+01*S3+6.190221e-02*S4+(-7.580406e-02)*S5+(-1.187791e-02)*S6+0.000000e+00*S7+(-1.506513e-01)*S8+9.355381e-02*S9'
.param V7_part2='V7_part1+1.460842e+01*S10+0.000000e+00*S11+6.814036e-02*S12+1.302196e-01*S13+6.025649e-02*S14+0.000000e+00*S15+0.000000e+00*S16+1.803998e+00*S17+5.633675e-02*S18+7.966547e+00*S19'
.param V7_part3='V7_part2+2.159551e+01*S20+1.136919e+01*S21+7.555822e+01*S22+1.100384e+01*S23+1.534491e-01*S24+1.523951e-01*S25+1.995494e-01*S26+1.423537e-01*S27+0.000000e+00*S28+3.496965e+01*S29'
.param V7='V7_part3+1.312035e-01*S30+3.061024e+01*S31+0.000000e+00*S32+4.622166e-02*S33+2.489361e+01*S34+2.205030e+01*S35+2.167665e-01*S36'
.param V8_part1='(-1.407021e+01)*S0+9.647000e+00*S1+7.651212e-03*S2+(-3.212230e-01)*S3+2.127174e-02*S4+1.352886e-04*S5+1.335118e-01*S6+0.000000e+00*S7+(-3.023261e-02)*S8+(-2.961875e-02)*S9'
.param V8_part2='V8_part1+(-2.343889e+00)*S10+0.000000e+00*S11+1.381542e-02*S12+(-3.120560e-02)*S13+2.496862e-02*S14+0.000000e+00*S15+0.000000e+00*S16+(-5.411856e-01)*S17+2.286663e-02*S18+(-5.908294e+00)*S19'
.param V8_part3='V8_part2+(-7.624145e+00)*S20+1.610484e+01*S21+(-4.737496e+01)*S22+(-6.397763e+00)*S23+4.737288e-02*S24+3.880565e-02*S25+(-1.624425e-02)*S26+3.428403e-02*S27+0.000000e+00*S28+(-1.087315e+01)*S29'
.param V8='V8_part3+(-5.110135e-02)*S30+(-1.345875e+01)*S31+0.000000e+00*S32+(-6.143377e-02)*S33+(-1.090480e+01)*S34+9.764329e-01*S35+3.873357e-02*S36'
.param V9_part1='0.000000e+00*S0+0.000000e+00*S1+(-2.425587e-03)*S2+0.000000e+00*S3+7.845951e-04*S4+(-3.831011e-02)*S5+6.054148e+00*S6+(-2.086892e-02)*S7+6.460101e+00*S8+(-2.286587e-02)*S9'
.param V9_part2='V9_part1+0.000000e+00*S10+6.681321e-02*S11+1.367791e-01*S12+6.699186e-02*S13+1.325310e-01*S14+(-1.876271e-02)*S15+(-2.469308e-02)*S16+0.000000e+00*S17+(-2.199189e-02)*S18+7.568486e+01*S19'
.param V9_part3='V9_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+4.048596e+01*S23+6.120767e-02*S24+7.460591e-02*S25+(-8.262422e-03)*S26+1.010589e-01*S27+1.880529e-01*S28+0.000000e+00*S29'
.param V9='V9_part3+1.841110e-01*S30+0.000000e+00*S31+7.165103e-02*S32+8.537364e-02*S33+0.000000e+00*S34+0.000000e+00*S35+1.413876e-01*S36'
.param V10_part1='0.000000e+00*S0+0.000000e+00*S1+1.490644e-02*S2+0.000000e+00*S3+2.225082e-02*S4+1.386896e-01*S5+(-3.168552e-01)*S6+(-5.095974e-03)*S7+(-6.857669e+00)*S8+(-6.440807e-04)*S9'
.param V10_part2='V10_part1+0.000000e+00*S10+3.503042e-02*S11+(-7.428659e-04)*S12+3.203221e-02*S13+1.316413e-02*S14+2.012345e-03*S15+2.633691e-02*S16+0.000000e+00*S17+1.978454e-02*S18+1.235518e+02*S19'
.param V10_part3='V10_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+(-5.123389e+01)*S23+4.413756e-02*S24+6.792172e-02*S25+7.653472e-02*S26+2.243909e-02*S27+9.444277e-02*S28+0.000000e+00*S29'
.param V10='V10_part3+3.190893e-02*S30+0.000000e+00*S31+4.745712e-02*S32+(-5.557110e-03)*S33+0.000000e+00*S34+0.000000e+00*S35+8.719907e-02*S36'
.param V11_part1='0.000000e+00*S0+0.000000e+00*S1+5.201878e-02*S2+0.000000e+00*S3+4.579999e-02*S4+7.601775e-03*S5+1.853511e-01*S6+6.331094e-02*S7+3.193963e+00*S8+6.161649e-02*S9'
.param V11_part2='V11_part1+0.000000e+00*S10+8.798116e-02*S11+6.149647e-02*S12+8.579121e-02*S13+5.641461e-02*S14+6.490333e-02*S15+6.306387e-02*S16+0.000000e+00*S17+6.206904e-02*S18+(-5.143032e+01)*S19'
.param V11_part3='V11_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+2.986609e+01*S23+8.929915e-02*S24+8.686272e-02*S25+1.030668e-01*S26+8.033623e-02*S27+1.021925e-01*S28+0.000000e+00*S29'
.param V11='V11_part3+1.036557e-01*S30+0.000000e+00*S31+8.460913e-02*S32+9.191755e-02*S33+0.000000e+00*S34+0.000000e+00*S35+1.032483e-01*S36'
.param V12_part1='(-1.547436e-03)*S0+3.483073e-03*S1+7.311562e+00*S2+5.059811e-03*S3+(-1.153938e+01)*S4+(-1.439174e-02)*S5+1.232271e-02*S6+6.996528e-02*S7+(-1.224737e-02)*S8+6.698200e-01*S9'
.param V12_part2='V12_part1+1.008465e-02*S10+6.376081e+00*S11+(-3.330483e+00)*S12+3.366684e+01*S13+5.245836e+00*S14+(-1.540133e+01)*S15+(-2.266094e+01)*S16+5.591986e-03*S17+(-1.126024e+01)*S18+(-3.486667e-02)*S19'
.param V12_part3='V12_part2+1.687755e-03*S20+7.379325e-03*S21+(-1.499264e-02)*S22+(-2.900244e-02)*S23+2.436838e+00*S24+6.066456e-01*S25+1.954778e+01*S26+4.262654e+00*S27+2.827834e+00*S28+(-9.598500e-02)*S29'
.param V12='V12_part3+4.885824e+01*S30+(-3.574099e-02)*S31+1.730601e+01*S32+(-7.821387e+00)*S33+(-3.332529e-02)*S34+1.953620e-02*S35+(-1.250170e-01)*S36'
.param V13_part1='4.722017e-01*S0+4.426868e-01*S1+2.313341e+01*S2+5.060677e-01*S3+2.504321e+02*S4+3.906250e-01*S5+3.245473e-01*S6+1.480806e+00*S7+3.532690e-01*S8+7.916999e-02*S9'
.param V13_part2='V13_part1+9.380649e-01*S10+7.038939e+01*S11+6.809913e+01*S12+5.286129e+01*S13+7.722867e+01*S14+1.879016e+02*S15+1.647047e+02*S16+5.610253e-01*S17+2.566462e+02*S18+6.859099e-01*S19'
.param V13_part3='V13_part2+1.646309e+00*S20+1.820255e+00*S21+2.008392e+00*S22+1.172803e+00*S23+6.850587e+01*S24+3.117518e+01*S25+3.714373e+01*S26+5.460962e+01*S27+1.357694e+02*S28+2.792664e+00*S29'
.param V13='V13_part3+5.516973e+02*S30+2.006786e+00*S31+2.430408e+02*S32+4.258481e+02*S33+2.881633e+00*S34+3.129545e+00*S35+6.026809e+02*S36'
.param V14_part1='(-1.768555e-02)*S0+(-6.061043e-02)*S1+(-6.562645e+00)*S2+(-1.170983e-01)*S3+(-5.169041e+01)*S4+(-1.429076e-02)*S5+(-5.675304e-02)*S6+(-2.484306e-01)*S7+(-4.777792e-02)*S8+(-5.917471e-02)*S9'
.param V14_part2='V14_part1+(-6.640791e-02)*S10+(-3.764296e+01)*S11+(-1.160959e+01)*S12+4.180840e+01*S13+(-3.297971e+01)*S14+(-2.421116e+01)*S15+(-1.387397e+01)*S16+(-3.731885e-02)*S17+(-5.160067e+01)*S18+(-7.009159e-02)*S19'
.param V14_part3='V14_part2+(-2.118289e-02)*S20+(-1.332026e-01)*S21+(-3.167635e-01)*S22+2.968973e-03*S23+(-3.161679e+01)*S24+(-5.949352e+00)*S25+4.115001e+01*S26+(-2.263831e+01)*S27+(-4.254578e+01)*S28+2.859600e-02*S29'
.param V14='V14_part3+(-6.088873e+02)*S30+5.757648e-02*S31+(-1.396133e+02)*S32+(-3.394597e+02)*S33+1.328776e-01*S34+(-8.182911e-02)*S35+(-5.328776e+02)*S36'
.param V15_part1='(-1.213710e-01)*S0+(-2.270748e-01)*S1+3.222086e+02*S2+(-3.679758e-01)*S3+8.692029e+01*S4+(-2.330815e-01)*S5+(-3.009752e-01)*S6+(-1.825580e+01)*S7+(-3.698413e-01)*S8+6.033068e-01*S9'
.param V15_part2='V15_part1+(-1.185175e-01)*S10+(-9.420818e+02)*S11+(-5.382300e+02)*S12+1.096670e+03*S13+(-6.407719e+02)*S14+(-1.723080e+03)*S15+(-5.543790e+02)*S16+(-9.545898e-02)*S17+1.103715e+02*S18+(-2.397593e-01)*S19'
.param V15_part3='V15_part2+(-2.019064e-01)*S20+(-4.909970e-01)*S21+(-1.049428e+00)*S22+(-1.780332e-01)*S23+(-8.015023e+02)*S24+(-1.343628e+02)*S25+1.291563e+03*S26+(-3.969294e+02)*S27+(-1.182991e+03)*S28+(-6.182841e-01)*S29'
.param V15='V15_part3+(-8.938264e+03)*S30+(-2.240164e-01)*S31+(-3.325987e+03)*S32+(-8.080653e+03)*S33+(-2.111899e-01)*S34+(-6.529066e-01)*S35+(-6.112769e+03)*S36'
.param V16_part1='6.429504e-01*S0+5.872554e-01*S1+7.398157e+00*S2+5.721275e-01*S3+1.218061e+03*S4+1.163697e+00*S5+3.451777e-01*S6+6.226717e+01*S7+6.342735e-01*S8+2.376741e+01*S9'
.param V16_part2='V16_part1+9.960250e-01*S10+9.340832e+02*S11+8.321411e+02*S12+(-1.595284e+02)*S13+6.344869e+02*S14+7.128556e+03*S15+2.536966e+03*S16+3.621895e-01*S17+1.879370e+03*S18+4.079078e-01*S19'
.param V16_part3='V16_part2+1.469921e+00*S20+1.411126e+00*S21+1.494970e+00*S22+1.165148e+00*S23+9.285133e+02*S24+2.494749e+02*S25+(-5.129468e+02)*S26+3.446753e+02*S27+2.398120e+03*S28+1.826653e+00*S29'
.param V16='V16_part3+6.702819e+03*S30+1.630000e+00*S31+3.424471e+03*S32+5.002608e+03*S33+1.999076e+00*S34+1.999898e+00*S35+4.831425e+03*S36'
.param V17_part1='9.949088e-02*S0+1.599476e-01*S1+1.849945e+02*S2+2.332899e-01*S3+2.076539e+03*S4+6.198086e-02*S5+2.193364e-01*S6+6.996832e+00*S7+1.255278e-01*S8+2.167375e+01*S9'
.param V17_part2='V17_part1+1.603757e-01*S10+5.527475e+02*S11+4.252770e+02*S12+5.654680e+02*S13+5.965473e+02*S14+4.521117e+02*S15+4.871341e+02*S16+1.836928e-01*S17+1.226897e+03*S18+2.833952e-01*S19'
.param V17_part3='V17_part2+2.454752e-01*S20+3.837946e-01*S21+6.024695e-01*S22+1.932186e-01*S23+4.260144e+02*S24+1.581469e+02*S25+1.843708e+02*S26+4.133332e+02*S27+4.829115e+02*S28+5.093233e-01*S29'
.param V17='V17_part3+3.213836e+03*S30+2.698688e-01*S31+1.571832e+03*S32+3.518251e+03*S33+3.455652e-01*S34+5.426185e-01*S35+2.702626e+03*S36'
.param V18_part1='0.000000e+00*S0+5.643813e-03*S1+3.811886e+00*S2+(-3.915235e-02)*S3+(-1.978642e+01)*S4+2.260778e-01*S5+0.000000e+00*S6+5.260471e-01*S7+(-1.720121e-03)*S8+7.612613e-01*S9'
.param V18_part2='V18_part1+(-1.678175e-02)*S10+2.759373e+00*S11+(-8.445236e-01)*S12+7.617809e+00*S13+1.677629e+00*S14+(-1.352018e+00)*S15+2.468166e+00*S16+(-2.354906e-02)*S17+2.578876e+00*S18+0.000000e+00*S19'
.param V18_part3='V18_part2+(-2.285313e-02)*S20+(-6.658113e-02)*S21+(-6.939470e-02)*S22+1.729910e-02*S23+(-1.765335e-01)*S24+(-5.444092e-01)*S25+(-8.132826e+00)*S26+(-5.705764e-02)*S27+2.066502e+00*S28+4.774686e-02*S29'
.param V18='V18_part3+(-3.302003e+01)*S30+0.000000e+00*S31+1.365576e+01*S32+3.082385e+01*S33+2.378342e-02*S34+(-8.055366e-02)*S35+(-3.159364e+00)*S36'
.param V19_part1='0.000000e+00*S0+6.347549e-02*S1+1.355943e-02*S2+8.600531e-02*S3+1.068953e+02*S4+(-2.542954e-01)*S5+0.000000e+00*S6+1.709128e-02*S7+1.643468e-02*S8+9.952366e-02*S9'
.param V19_part2='V19_part1+8.685999e-02*S10+8.004273e+00*S11+1.684518e+01*S12+(-8.043260e+00)*S13+2.035195e+01*S14+3.810405e+01*S15+1.992200e+01*S16+7.229787e-02*S17+4.119826e+01*S18+0.000000e+00*S19'
.param V19_part3='V19_part2+8.128475e-02*S20+1.456801e-01*S21+1.117288e-01*S22+1.163311e-01*S23+1.152498e+01*S24+3.534840e+00*S25+(-4.425025e-01)*S26+9.391450e+00*S27+2.115750e+01*S28+9.855141e-02*S29'
.param V19='V19_part3+1.551120e+02*S30+0.000000e+00*S31+6.193623e+01*S32+1.060184e+02*S33+1.190662e-01*S34+2.302605e-01*S35+1.254062e+02*S36'
.param V20_part1='0.000000e+00*S0+1.206310e-02*S1+(-2.435234e+00)*S2+3.260493e-02*S3+(-1.772983e+01)*S4+1.872315e-02*S5+0.000000e+00*S6+2.737676e-02*S7+(-3.990655e-02)*S8+5.141264e-02*S9'
.param V20_part2='V20_part1+2.890281e-02*S10+(-7.084747e+00)*S11+(-1.719240e+00)*S12+5.511361e+01*S13+(-8.557262e+00)*S14+(-8.320645e+00)*S15+(-9.793337e+00)*S16+8.594554e-03*S17+(-1.125384e+01)*S18+0.000000e+00*S19'
.param V20_part3='V20_part2+7.133094e-02*S20+1.277135e-02*S21+(-1.302667e-02)*S22+1.725436e-02*S23+(-3.896270e+00)*S24+1.538425e-01*S25+3.331515e+01*S26+(-2.927829e+00)*S27+(-9.312914e+00)*S28+(-1.151696e-01)*S29'
.param V20='V20_part3+(-9.638155e+01)*S30+0.000000e+00*S31+(-5.209969e+01)*S32+(-1.450825e+02)*S33+6.159206e-02*S34+3.067303e-02*S35+(-1.027379e+02)*S36'
.param V21_part1='(-2.528566e-02)*S0+(-1.803017e-02)*S1+0.000000e+00*S2+(-3.300505e-02)*S3+9.431467e+01*S4+4.427523e+00*S5+1.773751e-02*S6+1.821479e+01*S7+8.955526e-03*S8+(-6.121078e-01)*S9'
.param V21_part2='V21_part1+6.671034e-02*S10+0.000000e+00*S11+2.335240e+02*S12+1.504711e+03*S13+7.239096e+01*S14+0.000000e+00*S15+0.000000e+00*S16+(-7.963439e-03)*S17+0.000000e+00*S18+9.992604e-03*S19'
.param V21_part3='V21_part2+7.024625e-02*S20+1.120080e-02*S21+9.844869e-02*S22+8.546427e-02*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+1.245674e-01*S29'
.param V21='V21_part3+0.000000e+00*S30+7.828706e-02*S31+0.000000e+00*S32+0.000000e+00*S33+1.727911e-01*S34+7.001192e-02*S35+0.000000e+00*S36'
.param V22_part1='6.318633e-03*S0+(-7.436802e-03)*S1+0.000000e+00*S2+7.027681e-03*S3+1.765893e+03*S4+(-1.026802e+01)*S5+1.642725e-02*S6+(-2.195255e+01)*S7+(-1.344817e-01)*S8+9.538593e+00*S9'
.param V22_part2='V22_part1+2.417519e-02*S10+0.000000e+00*S11+(-9.524690e+01)*S12+(-8.701084e+02)*S13+1.618533e+01*S14+0.000000e+00*S15+0.000000e+00*S16+4.227152e-02*S17+0.000000e+00*S18+2.207718e-02*S19'
.param V22_part3='V22_part2+6.945125e-02*S20+8.003568e-02*S21+2.346731e-03*S22+4.177157e-02*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+1.129765e-01*S29'
.param V22='V22_part3+0.000000e+00*S30+6.495593e-02*S31+0.000000e+00*S32+0.000000e+00*S33+1.408741e-01*S34+1.435279e-01*S35+0.000000e+00*S36'
.param V23_part1='6.524088e-02*S0+6.443809e-02*S1+0.000000e+00*S2+6.855382e-02*S3+(-1.487592e+02)*S4+3.148806e+00*S5+1.006187e-02*S6+6.332818e+00*S7+7.903697e-02*S8+6.863198e+00*S9'
.param V23_part2='V23_part1+8.767509e-02*S10+0.000000e+00*S11+(-7.249947e+01)*S12+(-2.090834e+02)*S13+(-2.239257e+01)*S14+0.000000e+00*S15+0.000000e+00*S16+5.576089e-02*S17+0.000000e+00*S18+4.769262e-02*S19'
.param V23_part3='V23_part2+8.558765e-02*S20+1.024552e-01*S21+8.504741e-02*S22+8.103332e-02*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+1.154325e-01*S29'
.param V23='V23_part3+0.000000e+00*S30+8.358917e-02*S31+0.000000e+00*S32+0.000000e+00*S33+1.018129e-01*S34+1.276402e-01*S35+0.000000e+00*S36'
.param V24_part1='6.045859e-01*S0+1.033665e+00*S1+9.403763e-01*S2+7.242001e-01*S3+8.321871e-01*S4+2.090504e+00*S5+6.052696e+00*S6+5.394935e-01*S7+(-4.557807e-01)*S8+6.650049e-01*S9'
.param V24_part2='V24_part1+1.118244e+00*S10+1.342262e+00*S11+1.118129e+00*S12+1.124725e+00*S13+1.345292e+00*S14+1.144009e+00*S15+1.288692e+00*S16+1.260310e+00*S17+1.201624e+00*S18+1.213487e+00*S19'
.param V24_part3='V24_part2+1.218062e+00*S20+1.369381e+00*S21+1.684343e+00*S22+1.526487e+00*S23+1.335913e+00*S24+1.152789e+00*S25+1.007341e+00*S26+1.799705e+00*S27+1.541443e+00*S28+2.605297e+00*S29'
.param V24='V24_part3+2.117792e+00*S30+1.529031e+00*S31+1.728554e+00*S32+1.798580e+00*S33+2.032023e+00*S34+1.602337e+00*S35+1.755214e+00*S36'
.param V25_part1='7.507891e-01*S0+3.900675e-01*S1+4.080287e-01*S2+5.473841e-01*S3+2.343611e-01*S4+4.618813e-01*S5+7.805730e-01*S6+1.983233e-01*S7+6.115539e+00*S8+3.281980e+00*S9'
.param V25_part2='V25_part1+1.464269e+00*S10+4.778314e-01*S11+6.957581e-01*S12+1.093250e+00*S13+3.952433e-01*S14+4.212896e-01*S15+2.993568e-01*S16+9.892575e-01*S17+5.627475e-01*S18+2.632487e-01*S19'
.param V25_part3='V25_part2+1.642699e+00*S20+1.960783e+00*S21+9.836510e-01*S22+1.487340e+00*S23+1.362358e+00*S24+1.682956e+00*S25+1.595705e+00*S26+6.870965e-01*S27+1.549974e+00*S28+2.095816e+00*S29'
.param V25='V25_part3+1.278887e+00*S30+1.413111e+00*S31+9.827587e-01*S32+8.934959e-01*S33+2.244586e+00*S34+2.937726e+00*S35+1.892038e+00*S36'
.param V26_part1='(-2.260075e-01)*S0+(-4.939030e-02)*S1+4.002041e-02*S2+3.595049e-02*S3+4.622656e-02*S4+(-6.566245e-01)*S5+(-4.023143e+00)*S6+3.324479e-02*S7+(-9.123353e-01)*S8+(-1.218443e+00)*S9'
.param V26_part2='V26_part1+(-1.863040e-01)*S10+(-2.912175e-01)*S11+(-1.682442e-01)*S12+(-1.069584e+00)*S13+(-7.268979e-02)*S14+(-1.674616e-01)*S15+(-2.553138e-01)*S16+(-1.396352e-01)*S17+(-3.407645e-01)*S18+(-1.469223e-01)*S19'
.param V26_part3='V26_part2+1.565416e-01*S20+(-1.422294e+00)*S21+(-1.216066e+00)*S22+(-1.616989e-01)*S23+1.335185e-01*S24+3.961576e-02*S25+(-1.159242e+00)*S26+4.186072e-02*S27+(-4.933535e-01)*S28+(-3.153335e+00)*S29'
.param V26='V26_part3+(-1.948673e+00)*S30+(-6.375363e-01)*S31+(-9.341795e-01)*S32+(-1.131420e+00)*S33+(-5.077758e-01)*S34+(-2.033687e+00)*S35+(-1.665446e+00)*S36'
.param V27_part1='2.650448e+00*S0+8.172523e+03*S1+3.768178e+00*S2+(-1.060278e+00)*S3+(-1.363696e+00)*S4+(-1.983924e+00)*S5+(-8.007341e+00)*S6+1.321883e-01*S7+9.283287e+00*S8+1.241313e+00*S9'
.param V27_part2='V27_part1+(-8.140756e+00)*S10+3.957590e+00*S11+(-2.363310e-01)*S12+(-3.099922e+00)*S13+(-5.640105e+00)*S14+2.113181e+01*S15+9.764300e+00*S16+2.159061e+00*S17+(-9.874548e+00)*S18+7.490406e+00*S19'
.param V27_part3='V27_part2+(-3.795402e+00)*S20+(-1.669387e+00)*S21+(-3.294367e-01)*S22+2.029860e+01*S23+(-2.017487e+00)*S24+1.742769e-02*S25+(-2.443223e-01)*S26+(-3.426776e+00)*S27+6.002092e+00*S28+9.572005e+01*S29'
.param V27='V27_part3+(-6.998631e+00)*S30+1.933793e+01*S31+4.265936e+01*S32+8.496396e+01*S33+4.044263e+02*S34+(-8.989411e+00)*S35+(-1.520898e+01)*S36'
.param V28_part1='6.073495e-01*S0+8.172523e+03*S1+(-4.794947e-01)*S2+3.883510e+00*S3+6.322480e+00*S4+(-1.139270e+01)*S5+(-3.509598e+00)*S6+1.084715e-01*S7+(-1.492765e+01)*S8+(-6.428997e-01)*S9'
.param V28_part2='V28_part1+2.646805e+01*S10+1.211362e+00*S11+1.133748e+01*S12+7.572401e+00*S13+1.366268e+01*S14+(-2.006217e+01)*S15+(-2.655708e+00)*S16+8.422581e+00*S17+1.600667e+01*S18+(-3.410966e-01)*S19'
.param V28_part3='V28_part2+2.592672e+01*S20+1.051863e+01*S21+9.726762e+00*S22+(-1.252724e-01)*S23+1.267514e+01*S24+6.527443e+00*S25+3.839975e+00*S26+1.243241e+01*S27+9.383103e+00*S28+(-2.050821e+01)*S29'
.param V28='V28_part3+2.035039e+01*S30+3.021476e+00*S31+(-1.295395e+01)*S32+(-5.320133e+00)*S33+(-2.933128e+02)*S34+2.149750e+01*S35+2.654276e+01*S36'
.param V29_part1='(-1.128722e+00)*S0+(-3.286583e+00)*S1+(-8.552584e-01)*S2+6.570560e+00*S3+3.139925e+00*S4+(-9.873774e+00)*S5+7.265015e-01*S6+(-2.691873e-01)*S7+(-1.516065e+01)*S8+(-2.600423e-01)*S9'
.param V29_part2='V29_part1+2.391645e+01*S10+(-1.353663e+00)*S11+1.841457e+00*S12+1.012057e+01*S13+1.114463e+01*S14+(-4.818681e+00)*S15+(-3.204116e+00)*S16+9.464785e-01*S17+2.381166e+01*S18+(-1.859417e+00)*S19'
.param V29_part3='V29_part2+1.404885e+01*S20+8.159405e+00*S21+5.892827e-01*S22+(-1.686858e+01)*S23+4.307946e+00*S24+8.396721e-01*S25+2.003928e+00*S26+4.150301e+00*S27+(-5.502560e+00)*S28+(-1.097026e+02)*S29'
.param V29='V29_part3+1.048109e+01*S30+(-1.760187e+01)*S31+(-2.542986e+01)*S32+(-1.066048e+02)*S33+(-4.378715e+02)*S34+2.087815e+01*S35+1.868136e+01*S36'
.param V30_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+1.200673e+01*S3+0.000000e+00*S4+1.246807e+00*S5+1.008778e+00*S6+1.611480e+01*S7+6.025347e+00*S8+1.844555e+01*S9'
.param V30_part2='V30_part1+0.000000e+00*S10+1.949108e+01*S11+0.000000e+00*S12+6.727427e+00*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V30_part3='V30_part2+1.266680e+01*S20+1.821371e+01*S21+8.399211e+01*S22+1.595383e+00*S23+1.057744e+01*S24+2.247208e+00*S25+3.930634e+01*S26+2.527897e+01*S27+4.307099e+01*S28+2.736069e+01*S29'
.param V30='V30_part3+1.246395e+02*S30+3.184204e+01*S31+3.572729e+01*S32+6.766789e+01*S33+2.153057e+01*S34+(-6.190068e+01)*S35+(-1.505004e+01)*S36'
.param V31_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+4.274170e+00*S3+0.000000e+00*S4+5.441936e+00*S5+4.651726e+00*S6+(-5.449248e+00)*S7+(-4.190858e+00)*S8+(-1.240537e+01)*S9'
.param V31_part2='V31_part1+0.000000e+00*S10+5.873723e+01*S11+0.000000e+00*S12+6.120391e+01*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V31_part3='V31_part2+9.444409e+01*S20+7.287708e+01*S21+(-8.209763e+00)*S22+6.922999e+01*S23+7.647074e+01*S24+8.720557e+01*S25+7.199240e+01*S26+5.601942e+01*S27+1.527145e+02*S28+(-1.437959e+01)*S29'
.param V31='V31_part3+(-4.463023e+01)*S30+7.254921e+01*S31+1.701945e+01*S32+1.091420e+01*S33+1.525648e+02*S34+2.038222e+02*S35+1.407221e+02*S36'
.param V32_part1='0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+(-2.410646e+01)*S3+0.000000e+00*S4+1.427679e+01*S5+1.275030e+01*S6+2.777793e+00*S7+1.076181e+01*S8+2.367315e+00*S9'
.param V32_part2='V32_part1+0.000000e+00*S10+(-7.091702e+01)*S11+0.000000e+00*S12+(-6.383004e+01)*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V32_part3='V32_part2+(-4.978978e+01)*S20+(-5.240794e+01)*S21+(-3.110418e+01)*S22+(-1.000857e+01)*S23+(-3.974371e+01)*S24+(-2.326756e+01)*S25+(-1.117460e+02)*S26+(-2.996530e+01)*S27+(-8.914045e+01)*S28+9.419122e+01*S29'
.param V32='V32_part3+(-1.934466e+00)*S30+(-8.013437e+01)*S31+(-2.104252e+01)*S32+(-3.456294e+01)*S33+(-2.933252e+01)*S34+1.300083e+01*S35+2.851181e+01*S36'
.param V33_part1='(-1.527990e+01)*S0+1.796925e+01*S1+(-1.374756e+01)*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V33_part2='V33_part1+(-1.820819e+01)*S10+0.000000e+00*S11+1.645961e+01*S12+(-4.378196e+01)*S13+(-2.292053e+00)*S14+0.000000e+00*S15+0.000000e+00*S16+(-2.100267e+01)*S17+3.171789e+01*S18+0.000000e+00*S19'
.param V33_part3='V33_part2+2.560703e+01*S20+0.000000e+00*S21+(-2.066718e+02)*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+(-4.630372e+01)*S27+0.000000e+00*S28+(-9.035285e+01)*S29'
.param V33='V33_part3+(-3.041790e+02)*S30+(-7.412489e+01)*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+8.416391e+01*S35+0.000000e+00*S36'
.param V34_part1='8.844836e+01*S0+8.706219e+01*S1+(-1.171161e+01)*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V34_part2='V34_part1+5.426962e+01*S10+0.000000e+00*S11+5.877932e+01*S12+1.631506e+01*S13+5.713665e+00*S14+0.000000e+00*S15+0.000000e+00*S16+(-1.183157e+01)*S17+2.251548e+01*S18+0.000000e+00*S19'
.param V34_part3='V34_part2+3.180417e+01*S20+0.000000e+00*S21+2.195924e+02*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+5.818496e+01*S27+0.000000e+00*S28+3.183529e+02*S29'
.param V34='V34_part3+3.788865e+02*S30+9.481493e+01*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+(-6.695848e+01)*S35+0.000000e+00*S36'
.param V35_part1='2.220023e+01*S0+(-8.679919e+01)*S1+4.398731e+01*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9'
.param V35_part2='V35_part1+6.762397e+01*S10+0.000000e+00*S11+5.057439e+01*S12+2.190512e+02*S13+2.595490e+01*S14+0.000000e+00*S15+0.000000e+00*S16+5.696627e+01*S17+(-7.010229e+01)*S18+0.000000e+00*S19'
.param V35_part3='V35_part2+(-1.165793e+01)*S20+0.000000e+00*S21+2.179696e+02*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+1.370568e+01*S27+0.000000e+00*S28+(-1.109975e+00)*S29'
.param V35='V35_part3+2.254542e+02*S30+2.442006e+02*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+1.242570e+02*S35+0.000000e+00*S36'
.param V36_part1='(-1.799772e+01)*S0+(-2.463387e+01)*S1+(-1.997622e+00)*S2+(-4.274404e+00)*S3+(-3.247762e+00)*S4+(-1.748693e+00)*S5+1.767212e+00*S6+1.439112e+00*S7+(-1.598541e-01)*S8+(-7.929616e-01)*S9'
.param V36_part2='V36_part1+(-1.192730e+00)*S10+(-7.508709e+00)*S11+(-1.310877e+01)*S12+(-5.134941e+01)*S13+(-9.792038e+00)*S14+(-3.369242e+00)*S15+(-4.298787e+00)*S16+(-2.465092e+00)*S17+(-8.806353e+00)*S18+(-2.319515e+00)*S19'
.param V36_part3='V36_part2+(-4.530019e+01)*S20+(-1.245697e+01)*S21+(-3.334785e+03)*S22+(-2.495348e+00)*S23+(-6.021957e+00)*S24+(-5.741722e+00)*S25+(-2.514715e+01)*S26+(-8.407477e+00)*S27+(-5.480895e+01)*S28+(-3.168691e+02)*S29'
.param V36='V36_part3+(-3.334531e+03)*S30+(-2.630161e+00)*S31+(-1.035395e+01)*S32+(-1.849590e+01)*S33+(-8.130966e+00)*S34+(-3.717714e+00)*S35+(-1.523531e+01)*S36'
.param V37_part1='(-3.342442e+00)*S0+1.138503e+00*S1+1.191799e+01*S2+7.206053e+00*S3+1.033965e+01*S4+4.460457e+00*S5+1.764043e-02*S6+2.144013e-01*S7+1.441989e+00*S8+1.911493e+00*S9'
.param V37_part2='V37_part1+2.391228e+01*S10+2.616166e+00*S11+2.652844e+01*S12+1.098291e+00*S13+2.149925e+01*S14+1.285448e+01*S15+1.711930e+01*S16+1.963622e+01*S17+9.856249e+00*S18+1.214799e+01*S19'
.param V37_part3='V37_part2+(-6.726515e-01)*S20+1.039640e+01*S21+3.131485e+00*S22+4.836425e+00*S23+1.156588e+00*S24+2.195907e+00*S25+4.497236e+00*S26+1.508708e+00*S27+(-4.872911e-01)*S28+1.768124e+00*S29'
.param V37='V37_part3+3.227762e+00*S30+7.098989e-01*S31+2.087061e+01*S32+2.205094e+01*S33+2.423880e+00*S34+(-3.084375e+00)*S35+6.006209e+00*S36'
.param V38_part1='6.102175e+01*S0+7.407144e+01*S1+1.204965e+00*S2+1.109615e+01*S3+5.061771e+00*S4+4.621244e+00*S5+(-1.111326e+00)*S6+(-2.490885e-01)*S7+9.123046e-01*S8+1.458289e+00*S9'
.param V38_part2='V38_part1+7.223794e+00*S10+2.713219e+01*S11+7.711038e+00*S12+1.534808e+02*S13+1.123104e+01*S14+9.408070e+00*S15+5.633342e+00*S16+9.117204e-01*S17+2.160867e+01*S18+5.096162e+00*S19'
.param V38_part3='V38_part2+1.382928e+02*S20+3.704166e+01*S21+1.000000e+04*S22+1.223277e+01*S23+2.213794e+01*S24+1.823234e+01*S25+7.086102e+01*S26+2.247525e+01*S27+1.668537e+02*S28+9.506440e+02*S29'
.param V38='V38_part3+1.000000e+04*S30+9.496059e+00*S31+1.857276e+01*S32+2.431680e+01*S33+2.810877e+01*S34+2.436349e+01*S35+5.240946e+01*S36'
.param V39_part1='(-1.586108e+00)*S0+6.110136e+00*S1+1.426634e+00*S2+3.276554e-01*S3+1.252248e+00*S4+1.315056e+01*S5+9.475041e+00*S6+2.445774e+01*S7+4.954741e+00*S8+5.081487e+00*S9'
.param V39_part2='V39_part1+1.710961e+01*S10+3.247398e-01*S11+9.869130e+00*S12+4.280451e+01*S13+(-2.207637e+00)*S14+2.529156e-01*S15+(-8.577171e-01)*S16+4.002374e+00*S17+3.680229e+00*S18+1.483556e+00*S19'
.param V39_part3='V39_part2+2.883532e+01*S20+(-7.695785e+00)*S21+4.670366e+01*S22+2.312776e+00*S23+2.696316e+00*S24+3.565664e+00*S25+1.409496e+01*S26+4.567322e+00*S27+3.108321e+01*S28+4.917684e+01*S29'
.param V39='V39_part3+3.558719e+01*S30+2.630017e+01*S31+1.690332e-01*S32+2.242075e-01*S33+2.631306e+00*S34+1.324482e+01*S35+(-2.003601e+01)*S36'
.param V40_part1='8.182183e+01*S0+4.659280e+01*S1+(-7.089086e-01)*S2+1.250171e+00*S3+1.060226e+00*S4+1.697736e+01*S5+(-9.234459e+00)*S6+(-1.944801e+01)*S7+(-4.866713e+00)*S8+(-4.096035e+00)*S9'
.param V40_part2='V40_part1+2.114857e+00*S10+2.203759e+00*S11+2.037388e+01*S12+2.199796e+01*S13+3.575559e+00*S14+(-6.644561e-01)*S15+8.820422e+00*S16+7.636991e-01*S17+2.125557e+00*S18+1.698294e+00*S19'
.param V40_part3='V40_part2+8.081174e+01*S20+7.211185e+00*S21+1.506305e+01*S22+1.378584e+01*S23+4.467489e+00*S24+3.321917e+00*S25+6.751297e+00*S26+2.912415e+00*S27+9.096316e+01*S28+3.185106e+01*S29'
.param V40='V40_part3+3.565122e+01*S30+8.907712e+01*S31+(-2.023966e-01)*S32+(-2.831187e-02)*S33+7.429200e+00*S34+5.806839e+01*S35+6.326420e+00*S36'
.param V41_part1='(-1.574659e+01)*S0+(-1.769559e+01)*S1+1.316482e+00*S2+1.000704e+00*S3+(-1.215485e+00)*S4+(-7.682409e+00)*S5+8.686377e+00*S6+(-4.964335e+00)*S7+1.962602e+00*S8+(-2.991424e-01)*S9'
.param V41_part2='V41_part1+9.576698e+00*S10+2.147376e-01*S11+(-9.173972e+00)*S12+(-1.494271e+01)*S13+8.856006e-01*S14+9.927803e+00*S15+(-8.389960e-01)*S16+1.814982e+00*S17+6.972257e-01*S18+(-1.659486e+00)*S19'
.param V41_part3='V41_part2+(-4.796400e+01)*S20+1.571590e+01*S21+8.328940e+00*S22+(-3.994215e+00)*S23+(-3.253222e+00)*S24+(-3.024452e+00)*S25+(-9.845219e+00)*S26+(-3.716718e+00)*S27+(-6.461327e+01)*S28+(-1.431405e+01)*S29'
.param V41='V41_part3+2.773705e+00*S30+(-4.802740e+01)*S31+4.842172e-01*S32+2.569350e-01*S33+(-5.324226e+00)*S34+(-1.992884e+01)*S35+5.185926e+01*S36'
.param V42_part1='0.000000e+00*S0+(-4.526250e+01)*S1+(-9.741270e+01)*S2+1.060598e+02*S3+(-1.077845e+02)*S4+0.000000e+00*S5+1.170229e+01*S6+(-4.514679e+00)*S7+1.356633e+00*S8+(-2.079245e+01)*S9'
.param V42_part2='V42_part1+(-9.560450e-01)*S10+(-1.608713e+02)*S11+(-7.008297e+01)*S12+0.000000e+00*S13+7.643979e+02*S14+(-3.016626e+01)*S15+8.014665e+01*S16+3.309318e+01*S17+(-5.471343e+01)*S18+7.248143e+01*S19'
.param V42_part3='V42_part2+(-7.598517e+01)*S20+3.574175e+02*S21+0.000000e+00*S22+3.610574e+01*S23+(-1.230292e+02)*S24+(-1.379470e+02)*S25+(-1.985885e+02)*S26+(-1.729835e+02)*S27+(-1.307697e+02)*S28+0.000000e+00*S29'
.param V42='V42_part3+0.000000e+00*S30+(-2.196347e+00)*S31+(-1.470718e+03)*S32+(-2.721295e+03)*S33+(-2.922454e+02)*S34+1.622903e+01*S35+3.652349e+02*S36'
.param V43_part1='0.000000e+00*S0+2.622268e+00*S1+4.613480e+02*S2+5.830200e+01*S3+2.233413e+02*S4+0.000000e+00*S5+7.063300e+00*S6+1.362136e+01*S7+3.082098e+01*S8+4.908557e+01*S9'
.param V43_part2='V43_part1+1.119097e+02*S10+(-2.165250e+01)*S11+1.768479e+02*S12+0.000000e+00*S13+3.142427e+00*S14+3.668141e+02*S15+8.507522e+01*S16+2.125377e+02*S17+8.909436e+01*S18+1.188219e+02*S19'
.param V43_part3='V43_part2+(-5.519498e+00)*S20+(-1.704413e+02)*S21+0.000000e+00*S22+(-3.558071e+01)*S23+(-2.762381e+01)*S24+(-6.909922e+00)*S25+2.873156e+01*S26+(-2.971468e+01)*S27+(-6.150028e+00)*S28+0.000000e+00*S29'
.param V43='V43_part3+0.000000e+00*S30+(-5.893495e+00)*S31+3.676688e+03*S32+3.285545e+03*S33+2.693570e+01*S34+(-3.736997e+01)*S35+(-1.056416e+02)*S36'
.param V44_part1='0.000000e+00*S0+1.348923e+02*S1+(-1.075991e+01)*S2+1.742949e+02*S3+3.839614e+02*S4+0.000000e+00*S5+(-2.192245e+01)*S6+(-1.271590e-01)*S7+(-1.086773e+01)*S8+1.347869e+01*S9'
.param V44_part2='V44_part1+2.436318e+01*S10+9.753300e+02*S11+3.322922e+01*S12+0.000000e+00*S13+2.641877e+01*S14+(-2.245344e+01)*S15+5.700962e+01*S16+(-6.205842e+01)*S17+2.395382e+02*S18+2.717733e+02*S19'
.param V44_part3='V44_part2+2.358831e+02*S20+1.229586e+02*S21+0.000000e+00*S22+1.393123e+02*S23+5.602296e+02*S24+4.859293e+02*S25+5.724981e+02*S26+5.485863e+02*S27+4.011604e+02*S28+0.000000e+00*S29'
.param V44='V44_part3+0.000000e+00*S30+1.557879e+01*S31+1.312722e+03*S32+2.557394e+03*S33+9.998615e+02*S34+3.658721e+01*S35+(-8.682581e+01)*S36'
.param V45_part1='(-8.051528e-01)*S0+3.421374e+00*S1+1.591845e+00*S2+(-1.108576e-01)*S3+(-3.137204e+00)*S4+(-3.521970e+00)*S5+(-6.136304e-02)*S6+(-1.441009e+00)*S7+(-1.627945e+00)*S8+(-6.225635e-01)*S9'
.param V45_part2='V45_part1+(-2.429134e+00)*S10+0.000000e+00*S11+(-2.575961e-01)*S12+(-7.233397e+00)*S13+0.000000e+00*S14+(-3.371559e-02)*S15+(-1.692960e+00)*S16+(-6.420431e+00)*S17+8.632935e-01*S18+(-8.857268e+00)*S19'
.param V45_part3='V45_part2+7.363075e+00*S20+0.000000e+00*S21+(-1.399344e+01)*S22+(-1.951760e+00)*S23+(-8.530934e-01)*S24+(-1.620456e+00)*S25+8.765652e+00*S26+(-5.210552e+00)*S27+1.308985e+01*S28+(-1.159015e+01)*S29'
.param V45='V45_part3+(-1.558772e+01)*S30+(-4.511984e+00)*S31+0.000000e+00*S32+2.048697e+01*S33+1.361668e+00*S34+(-1.269012e+01)*S35+(-1.111041e+01)*S36'
.param V46_part1='8.811881e+00*S0+9.427633e+00*S1+6.808398e-01*S2+3.951784e+00*S3+2.749025e+00*S4+7.364594e+00*S5+1.913900e+00*S6+6.887708e+00*S7+4.018669e+00*S8+4.006143e+00*S9'
.param V46_part2='V46_part1+2.772237e+00*S10+0.000000e+00*S11+5.219990e+00*S12+1.545702e+01*S13+0.000000e+00*S14+(-2.772809e+00)*S15+(-8.241680e-01)*S16+1.784088e+00*S17+6.345932e+00*S18+5.231444e+00*S19'
.param V46_part3='V46_part2+2.248865e+01*S20+0.000000e+00*S21+2.309615e+01*S22+1.509008e+01*S23+2.058015e+01*S24+2.377399e+01*S25+1.732111e+01*S26+2.427746e+01*S27+2.833500e+01*S28+2.759846e+01*S29'
.param V46='V46_part3+2.645054e+01*S30+2.484922e+01*S31+0.000000e+00*S32+(-1.516770e+01)*S33+2.987886e+01*S34+3.257901e+01*S35+2.347165e+01*S36'
.param V47_part1='7.757452e+00*S0+(-6.779936e+00)*S1+5.971398e+00*S2+(-5.923840e-01)*S3+5.704832e+00*S4+9.730005e+00*S5+8.221678e+00*S6+6.057337e+00*S7+8.340517e+00*S8+7.157744e+00*S9'
.param V47_part2='V47_part1+8.926256e+00*S10+0.000000e+00*S11+1.231544e+01*S12+2.811999e+01*S13+0.000000e+00*S14+5.202505e+00*S15+7.441707e+00*S16+1.530375e+01*S17+(-2.507320e+00)*S18+1.157660e+01*S19'
.param V47_part3='V47_part2+(-1.707974e+01)*S20+0.000000e+00*S21+3.852336e+01*S22+2.609134e+00*S23+(-6.397610e+00)*S24+(-4.388198e+00)*S25+(-2.888699e+01)*S26+6.514972e-01*S27+(-3.315479e+01)*S28+3.835773e+01*S29'
.param V47='V47_part3+4.883934e+01*S30+1.950646e+01*S31+0.000000e+00*S32+(-4.932878e+00)*S33+(-6.103719e+00)*S34+3.405179e+01*S35+1.488071e+01*S36'
.param V48_part1='0.000000e+00*S0+0.000000e+00*S1+7.912578e+00*S2+0.000000e+00*S3+1.392820e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+1.535572e-01*S8+1.086346e-02*S9'
.param V48_part2='V48_part1+1.057474e-01*S10+0.000000e+00*S11+1.301214e+01*S12+1.160431e+00*S13+0.000000e+00*S14+(-2.231557e-01)*S15+0.000000e+00*S16+4.103408e-01*S17+0.000000e+00*S18+2.254233e+00*S19'
.param V48_part3='V48_part2+(-5.699677e-01)*S20+0.000000e+00*S21+7.968591e-02*S22+7.767460e-01*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+1.443406e-01*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V48='V48_part3+0.000000e+00*S30+0.000000e+00*S31+(-8.762248e+00)*S32+0.000000e+00*S33+0.000000e+00*S34+2.910770e-02*S35+0.000000e+00*S36'
.param V49_part1='0.000000e+00*S0+0.000000e+00*S1+(-1.133716e-01)*S2+0.000000e+00*S3+(-3.693726e-01)*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+2.358834e-01*S8+1.844797e-01*S9'
.param V49_part2='V49_part1+4.510667e-02*S10+0.000000e+00*S11+3.979435e+01*S12+(-9.548987e-01)*S13+0.000000e+00*S14+8.120646e+00*S15+0.000000e+00*S16+1.174994e-01*S17+0.000000e+00*S18+(-7.040757e-01)*S19'
.param V49_part3='V49_part2+(-3.278831e-01)*S20+0.000000e+00*S21+(-4.853278e-03)*S22+(-1.694037e+00)*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+(-5.591588e-01)*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V49='V49_part3+0.000000e+00*S30+0.000000e+00*S31+1.630426e+03*S32+0.000000e+00*S33+0.000000e+00*S34+(-8.199943e-03)*S35+0.000000e+00*S36'
.param V50_part1='0.000000e+00*S0+0.000000e+00*S1+(-7.566958e+00)*S2+0.000000e+00*S3+(-4.564293e-01)*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+(-4.800556e-01)*S8+(-5.598650e-02)*S9'
.param V50_part2='V50_part1+8.548331e-02*S10+0.000000e+00*S11+2.146126e+01*S12+(-1.937522e-01)*S13+0.000000e+00*S14+(-2.740015e+00)*S15+0.000000e+00*S16+(-3.156208e-01)*S17+0.000000e+00*S18+(-1.075056e+00)*S19'
.param V50_part3='V50_part2+2.110584e+00*S20+0.000000e+00*S21+(-1.827978e-02)*S22+5.404073e-01*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+7.750703e-01*S27+0.000000e+00*S28+0.000000e+00*S29'
.param V50='V50_part3+0.000000e+00*S30+0.000000e+00*S31+3.501453e-01*S32+0.000000e+00*S33+0.000000e+00*S34+1.291064e-01*S35+0.000000e+00*S36'
.param V51_part1='1.000000e+04*S0+0.000000e+00*S1+(-1.018040e+02)*S2+0.000000e+00*S3+0.000000e+00*S4+2.330586e+03*S5+1.748013e+02*S6+0.000000e+00*S7+(-2.981781e+02)*S8+1.488108e+03*S9'
.param V51_part2='V51_part1+2.810451e+01*S10+0.000000e+00*S11+1.798021e+03*S12+(-1.581770e+03)*S13+3.084493e+03*S14+0.000000e+00*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V51_part3='V51_part2+0.000000e+00*S20+8.931375e+01*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+5.974402e-01*S29'
.param V51='V51_part3+6.579889e+02*S30+2.478158e+01*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36'
.param V52_part1='1.000000e+04*S0+0.000000e+00*S1+1.872819e+00*S2+0.000000e+00*S3+0.000000e+00*S4+1.000000e+04*S5+2.252289e+02*S6+0.000000e+00*S7+1.362577e+01*S8+(-1.118341e+03)*S9'
.param V52_part2='V52_part1+3.568573e+02*S10+0.000000e+00*S11+3.006383e+03*S12+4.142058e+03*S13+3.084493e+03*S14+0.000000e+00*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V52_part3='V52_part2+0.000000e+00*S20+6.233141e+02*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+(-4.395426e+02)*S29'
.param V52='V52_part3+8.403037e+03*S30+(-6.474152e+02)*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36'
.param V53_part1='1.000000e+04*S0+0.000000e+00*S1+3.015734e+02*S2+0.000000e+00*S3+0.000000e+00*S4+1.000000e+04*S5+1.276788e+02*S6+0.000000e+00*S7+1.080089e+03*S8+8.254745e-02*S9'
.param V53_part2='V53_part1+1.101202e+01*S10+0.000000e+00*S11+7.424737e+03*S12+8.519364e+00*S13+3.084493e+03*S14+0.000000e+00*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19'
.param V53_part3='V53_part2+0.000000e+00*S20+6.223888e+02*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+0.000000e+00*S26+0.000000e+00*S27+0.000000e+00*S28+9.374344e+02*S29'
.param V53='V53_part3+5.185897e+03*S30+1.083058e+03*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36'
.param _P0='V0+V1*radius_+V2*w_'
.param _P1='0.5*(_P0+sqrt(_P0*_P0+0.001))'
.param _P2='1e-09*_P1'
.param _P3='1e-09*_P1'
.param _P4='V3+V4*radius_+V5/w_'
.param _P5='0.5*(_P4+sqrt(_P4*_P4+0.001))'
.param _P6='V6+V7*radius_+V8*w_'
.param _P7='0.5*(_P6+sqrt(_P6*_P6+0.001))'
.param _P8='1e-09*_P7'
.param _P9='V9+V10*radius_+V11/w_'
.param _P10='0.5*(_P9+sqrt(_P9*_P9+0.001))'
.param _P11='V12+V13*radius_+V14*w_'
.param _P12='0.5*(_P11+sqrt(_P11*_P11+0.001))'
.param _P13='1e-09*_P12'
.param _P14='1e-09*_P12'
.param _P15='V15+V16*radius_+V17/w_'
.param _P16='0.5*(_P15+sqrt(_P15*_P15+0.001))'
.param _P17='V18+V19*radius_+V20*w_'
.param _P18='0.5*(_P17+sqrt(_P17*_P17+0.001))'
.param _P19='1e-09*_P18'
.param _P20='V21+V22*radius_+V23/w_'
.param _P21='0.5*(_P20+sqrt(_P20*_P20+0.001))'
.param _P22='V24+V25*radius_+V26*w_'
.param _P23='atan(_P22-0.5)/1.5708'
.param _P24='V27+V28*radius_+V29*w_'
.param _P25='atan(_P24-0.5)/1.5708'
.param _P26='0.5*_P23+0.5*_P25'
.param _P27='0.5*_P23-0.5*_P25'
.param _P28='V30+V31*radius_+V32*w_'
.param _P29='0.5*(_P28+sqrt(_P28*_P28+0.001))'
.param _P30='1e-15*_P29'
.param _P31='V33+V34*radius_+V35*w_'
.param _P32='0.5*(_P31+sqrt(_P31*_P31+0.001))'
.param _P33='1e-15*_P32'
.param _P34='1e-15*_P32'
.param _P35='V36+V37*radius_+V38*w_'
.param _P36='0.5*(_P35+sqrt(_P35*_P35+0.001))'
.param _P37='V39+V40*radius_+V41*w_'
.param _P38='0.5*(_P37+sqrt(_P37*_P37+0.001))'
.param _P39='V42+V43*radius_+V44*w_'
.param _P40='0.5*(_P39+sqrt(_P39*_P39+0.001))'
.param _P41='V45+V46*radius_+V47*w_'
.param _P42='0.5*(_P41+sqrt(_P41*_P41+0.001))'
.param _P43='V48+V49*radius_+V50*w_'
.param _P44='0.5*(_P43+sqrt(_P43*_P43+0.001))'
.param _P45='V51+V52*radius_+V53*w_'
.param _P46='0.5*(_P45+sqrt(_P45*_P45+0.001))'
.param _P47='1e-14*_P36'
.param _P48='100*_P38'
.param _P49='1e-15*_P40'
.param _P50='1e-14*_P36'
.param _P51='100*_P38'
.param _P52='1e-15*_P40'
.param _P53='1e-14*_P42'
.param _P54='100*_P44'
.param _P55='1e-15*_P46'
l1_sect1 PLUS _n1i_sect1 '_P2*(1+dls_diff_ind_3t_rf_pgs_psub_n)'
l2_sect1 _n2i_sect1 MINUS '_P3*(1+dls_diff_ind_3t_rf_pgs_psub_n)'
r1_sect1 _n1i_sect1 _n_sect1 '_P5*(1+drs_diff_ind_3t_rf_pgs_psub_n)' tc1=0.003
r2_sect1 _n_sect1 _n2i_sect1 '_P5*(1+drs_diff_ind_3t_rf_pgs_psub_n)' tc1=0.003
lc_sect1 _nc_sect1 CT '_P8*(1+dls_diff_ind_3t_rf_pgs_psub_n)'
rc_sect1 _n_sect1 _nc_sect1 '_P10*(1+drs_diff_ind_3t_rf_pgs_psub_n)' tc1=0.003
l1_sect2 PLUS _n1i_sect2 '_P13*(1+dls_diff_ind_3t_rf_pgs_psub_n)'
l2_sect2 _n2i_sect2 MINUS '_P14*(1+dls_diff_ind_3t_rf_pgs_psub_n)'
r1_sect2 _n1i_sect2 _n_sect2 '_P16*(1+drs_diff_ind_3t_rf_pgs_psub_n)' tc1=0.003
r2_sect2 _n_sect2 _n2i_sect2 '_P16*(1+drs_diff_ind_3t_rf_pgs_psub_n)' tc1=0.003
lc_sect2 _nc_sect2 CT '_P19*(1+dls_diff_ind_3t_rf_pgs_psub_n)'
rc_sect2 _n_sect2 _nc_sect2 '_P21*(1+drs_diff_ind_3t_rf_pgs_psub_n)' tc1=0.003
k12_sect1 l1_sect1 l2_sect1 K=_P26
k12_sect2 l1_sect2 l2_sect2 K=_P26
ks1s2_1 l1_sect1 l1_sect2 K=_P27
ks1s2_2 l2_sect1 l2_sect2 K=_P27
c12 PLUS MINUS '_P30'
c13 PLUS CT '_P33'
c23 MINUS CT '_P34'
c_1_sub PLUS _n1_1_sub '_P47'
rs_1_sub _n1_1_sub PSUB '_P48'
cs_1_sub _n1_1_sub PSUB '_P49'
c_2_sub MINUS _n1_2_sub '_P50'
rs_2_sub _n1_2_sub PSUB '_P51'
cs_2_sub _n1_2_sub PSUB '_P52'
c_3_sub CT _n1_3_sub '_P53'
rs_3_sub _n1_3_sub PSUB '_P54'
cs_3_sub _n1_3_sub PSUB '_P55'
kzero1 l1_sect1 l2_sect2 K=1e-6
kzero2 l1_sect2 l2_sect1 K=1e-6
.ends diff_ind_3t_rf_pgs_psub_n
