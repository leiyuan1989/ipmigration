
************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    DFFSR_X1
* View Name:    schematic
************************************************************************

.SUBCKT DFFSR_X1 CLK D Q RN SN VDD VSS
*.PININFO CLK:I D:I RN:I SN:I Q:O VDD:B VNW:B VPW:B VSS:B
mNM13 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM39 net5 rnb net4 VPW nch5 mr=1 l=600n w=220n nf=1
mM19 Q net2 VSS VPW nch5 mr=1 l=600n w=1.15u nf=1
mM38 net4 SN VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM17 net1 clkn net5 VPW nch5 mr=1 l=600n w=220n nf=1
mM25 net7 net10 net8 VPW nch5 mr=1 l=600n w=220n nf=1
mM31 net7 D net12 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM28 net12 clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM22 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM34 rnb RN VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM7 net9 SN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM32 net10 clkp net1 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM9 net2 net1 VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM10 net10 rnb net9 VPW nch5 mr=1 l=600n w=735n nf=1
mNM3 net10 net7 net9 VPW nch5 mr=1 l=600n w=735n nf=1
mM24 net8 clkp VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM42 net5 net2 net4 VPW nch5 mr=1 l=600n w=220n nf=1
mM29 net6 clkp VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM43 net5 net2 net3 VNW pch5 mr=1 l=500n w=220n nf=1
mM27 net13 clkn VDD VNW pch5 mr=1 l=500n w=220n nf=1
mPM13 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM16 net1 clkp net5 VNW pch5 mr=1 l=500n w=220n nf=1
mM35 rnb RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM26 net7 net10 net13 VNW pch5 mr=1 l=500n w=220n nf=1
mM23 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM40 net5 SN VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM33 net10 clkn net1 VNW pch5 mr=1 l=500n w=1.03u nf=1
mM18 Q net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM6 net10 SN VDD VNW pch5 mr=1 l=500n w=1.01u nf=1
mPM3 net10 net7 net11 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM11 net11 rnb VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM30 net7 D net6 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM41 net3 rnb VDD VNW pch5 mr=1 l=500n w=220n nf=1
mPM9 net2 net1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    EDFFR_X1
* View Name:    schematic
************************************************************************

.SUBCKT EDFFR_X1 CLK D E Q RN VDD VSS
*.PININFO CLK:I D:I E:I RN:I Q:O VDD:B VNW:B VPW:B VSS:B
mNM20 Q net2 VSS VPW nch5 mr=1 l=600n w=1.15u nf=1
mM22 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM16 net1 clkn VSS VPW nch5 mr=1 l=600n w=220n nf=1
mNM3 net11 D net12 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM17 net5 net6 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM13 net194 RN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM8 net10 E VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM5 net13 Q VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM4 net11 net10 net13 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM1 net2 net3 VSS VPW nch5 mr=1 l=600n w=780n nf=1
mNM2 net12 E VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM14 net7 net11 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM12 net5 clkp net3 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM9 net8 clkn net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM31 net9 clkp VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM30 net6 net5 net9 VPW nch5 mr=1 l=600n w=220n nf=1
mM12 net8 net7 net194 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM18 net3 net2 net1 VPW nch5 mr=1 l=600n w=220n nf=1
mNM15 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mPM20 Q net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM15 net7 net11 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM23 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM17 net14 clkp VDD VNW pch5 mr=1 l=500n w=300n nf=1
mPM5 net164 D VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM4 net164 E VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM2 net11 net10 net164 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM3 net11 Q net164 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM19 net3 net2 net14 VNW pch5 mr=1 l=500n w=300n nf=1
mPM15 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM17 net5 net6 VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mPM1 net2 net3 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM12 net5 clkn net3 VNW pch5 mr=1 l=500n w=1.68u nf=1
mPM9 net8 clkp net6 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM9 net10 E VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM10 net8 net7 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM11 net8 RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM28 net4 clkn VDD VNW pch5 mr=1 l=500n w=300n nf=1
mM29 net6 net5 net4 VNW pch5 mr=1 l=500n w=300n nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    CLKGTP_X1
* View Name:    schematic
************************************************************************

.SUBCKT CLKGTP_X1 CLK E GCLK VDD VSS
*.PININFO CLK:I E:I GCLK:O VDD:B VNW:B VPW:B VSS:B
mM22 net1 net10 net11 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM21 net10 net8 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM19 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM13 GCLK net1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM23 net11 clkp VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM7 net2 clkp net4 VNW pch5 mr=1 l=500n w=500n nf=1
mM6 net4 net8 VDD VNW pch5 mr=1 l=500n w=500n nf=1
mM1 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM3 net2 clkn net3 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM1 net8 net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM2 net3 E VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM20 net10 net8 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM11 net1 clkp VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM18 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM12 GCLK net1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM10 net1 net10 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM9 net2 clkn net7 VPW nch5 mr=1 l=600n w=220n nf=1
mM8 net7 net8 VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM5 net2 clkp net9 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM4 net9 E VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM0 net8 net2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    LATSR_X1
* View Name:    schematic
************************************************************************

.SUBCKT LATSR_X1 D G Q RN SN VDD VSS
*.PININFO D:I E:I RN:I SN:I Q:O VDD:B VNW:B VPW:B VSS:B
mM11 net8 net2 net4 VPW nch5 mr=1 l=600n w=220n nf=1
mM10 net4 en VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM18 net1 net2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM21 net2 rnb net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM7 net6 SN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM29 en G VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM25 net8 D net5 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM3 net2 net8 net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 Q net1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM34 rnb RN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM16 enb en VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM20 net5 enb VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM13 net3 enb VDD VNW pch5 mr=1 l=500n w=500n nf=1
mM12 net8 net2 net3 VNW pch5 mr=1 l=500n w=500n nf=1
mPM3 net2 net8 net10 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM22 net10 rnb VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM6 net2 SN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM29 en G VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM19 net1 net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM31 net8 D net7 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM17 enb en VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM35 rnb RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM1 Q net1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM33 net7 en VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    SDFFSR_X1
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSR_X1 CLK D Q RN SE SI SN VDD VSS
*.PININFO CLK:I D:I RN:I SE:I SI:I SN:I Q:O VDD:B VNW:B VPW:B VSS:B
mM9 net4 SEN net11 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM7 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.68u nf=1
mM48 SEN SE VDD VNW pch5 mr=1 l=500n w=1.68u nf=1
mM11 net4 SE net14 VNW pch5 mr=1 l=500n w=1.68u nf=1
mM51 net2 SN VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM10 net14 D VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM50 net2 net6 net16 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM61 net1 net8 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM64 Q net1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM59 net2 clkn net8 VNW pch5 mr=1 l=500n w=1.68u nf=1
mM56 net6 net2 net15 VNW pch5 mr=1 l=500n w=220n nf=1
mM8 net11 SI VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM69 net5 net1 net10 VNW pch5 mr=1 l=500n w=220n nf=1
mM42 net6 clkp net4 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM46 rnb RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM49 net16 rnb VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM68 net10 rnb VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM67 net5 SN VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM55 net15 clkn VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM66 net8 clkp net5 VNW pch5 mr=1 l=500n w=220n nf=1
mM5 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM62 net1 net8 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM47 SEN SE VSS VPW nch5 mr=1 l=600n w=1.15u nf=1
mM53 net2 rnb net3 VPW nch5 mr=1 l=600n w=1.15u nf=1
mM6 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM15 net13 D VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM52 net2 net6 net3 VPW nch5 mr=1 l=600n w=780n nf=1
mM41 net6 clkn net9 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM14 net7 SI VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM16 net9 SEN net13 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM60 net2 clkp net8 VPW nch5 mr=1 l=600n w=780n nf=1
mM63 Q net1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM54 net3 SN VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM4 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 net9 SE net7 VPW nch5 mr=1 l=600n w=1.15u nf=1
mM57 net6 net2 net17 VPW nch5 mr=1 l=600n w=220n nf=1
mM45 rnb RN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM58 net17 clkp VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM71 net5 rnb net12 VPW nch5 mr=1 l=600n w=220n nf=1
mM70 net5 net1 net12 VPW nch5 mr=1 l=600n w=220n nf=1
mM72 net12 SN VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM65 net8 clkn net5 VPW nch5 mr=1 l=600n w=220n nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    SEDFFSR_X1
* View Name:    schematic
************************************************************************

.SUBCKT SEDFFSR_X1 CLK D E Q RN SE SI SN VDD VSS
*.PININFO CLK:I D:I E:I RN:I SE:I SI:I SN:I Q:O VDD:B VNW:B VPW:B VSS:B
mNM9 net010 clkn net013 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM14 seb SE VSS VPW nch5 mr=1 l=600n w=1.15u nf=1
mNM12 net12 clkp net15 VPW nch5 mr=1 l=600n w=1.15u nf=1
mM61 net060 RN net017 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM48 net060 seb net010 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM37 net15 clkn net26 VPW nch5 mr=1 l=600n w=220n nf=1
mM24 Q net20 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM35 net013 clkp net28 VPW nch5 mr=1 l=600n w=220n nf=1
mM42 net12 net013 VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM36 net26 net20 VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM8 eb E VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM12 net010 SE net059 VPW nch5 mr=1 l=600n w=1.15u nf=1
mM44 net20 net15 VSS VPW nch5 mr=1 l=600n w=860n nf=1
mM49 net017 Q net047 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM3 net049 D VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM39 clkp clkn VSS VPW nch5 mr=1 l=600n w=780n nf=1
mNM1 clkn CLK VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM32 net28 net12 VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM1 snb SN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM4 net060 snb VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM50 net047 eb VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 net017 E net049 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM11 net059 SI VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM62 net058 SI VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mPM9 net010 clkp net013 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM40 net15 clkp net25 VNW pch5 mr=1 l=500n w=220n nf=1
mM33 net013 clkn net27 VNW pch5 mr=1 l=500n w=220n nf=1
mM15 seb SE VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM65 net048 eb net1 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM58 net010 seb net058 VNW pch5 mr=1 l=500n w=1.25u nf=1
mM43 net12 net013 VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM31 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM38 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM60 net046 E net1 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM64 net060 RN net1 VNW pch5 mr=1 l=500n w=1.31u nf=1
mPM1 net20 net15 VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM18 net1 snb VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM54 net060 D net048 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM9 eb E VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM63 net060 SE net010 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM66 net060 Q net046 VNW pch5 mr=1 l=500n w=1.68u nf=1
mPM12 net12 clkn net15 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM41 net25 net20 VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM34 net27 net12 VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM2 snb SN VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM45 Q net20 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
.ENDS