* SPICE INPUT		Tue Sep 18 13:23:08 2018	drfcrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfcrb0
.subckt drfcrb0 VDD VDDG GND Q QN RN D RETN CK
M1 GND N_9 N_5 GND mn15  l=0.13u w=0.2u m=1
M2 N_41 N_9 N_11 GND mn15  l=0.13u w=0.32u m=1
M3 N_41 D GND GND mn15  l=0.13u w=0.32u m=1
M4 GND CK N_9 GND mn15  l=0.13u w=0.22u m=1
M5 N_11 N_5 N_36 GND mn15  l=0.13u w=0.26u m=1
M6 GND N_16 N_36 GND mn15  l=0.13u w=0.26u m=1
M7 N_16 N_11 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_16 N_5 N_14 GND mn15  l=0.13u w=0.26u m=1
M9 N_14 N_19 GND GND mn15  l=0.13u w=0.26u m=1
M10 N_18 N_14 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_19 RN GND GND mn15  l=0.13u w=0.26u m=1
M12 N_50 N_24 GND GND mn15  l=0.13u w=0.26u m=1
M13 N_14 N_9 N_50 GND mn15  l=0.13u w=0.26u m=1
M14 N_24 RETN N_18 GND mn15  l=0.13u w=0.26u m=1
M15 Q N_18 GND GND mn15  l=0.13u w=0.26u m=1
M16 QN N_14 GND GND mn15  l=0.13u w=0.26u m=1
M17 N_30 RETN GND GND mn15  l=0.13u w=0.26u m=1
M18 N_29 N_24 GND GND mn15  l=0.13u w=0.26u m=1
M19 GND N_29 N_60 GND mn15  l=0.13u w=0.26u m=1
M20 N_24 N_30 N_60 GND mn15  l=0.13u w=0.26u m=1
M21 VDD N_9 N_5 VDD mp15  l=0.13u w=0.51u m=1
M22 N_73 D VDD VDD mp15  l=0.13u w=0.4u m=1
M23 N_11 N_9 N_72 VDD mp15  l=0.13u w=0.26u m=1
M24 N_9 CK VDD VDD mp15  l=0.13u w=0.56u m=1
M25 N_73 N_5 N_11 VDD mp15  l=0.13u w=0.4u m=1
M26 VDD N_16 N_72 VDD mp15  l=0.13u w=0.26u m=1
M27 N_18 N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_19 RN VDD VDD mp15  l=0.13u w=0.4u m=1
M29 N_16 N_11 N_70 VDD mp15  l=0.13u w=0.4u m=1
M30 N_74 N_24 N_70 VDD mp15  l=0.13u w=0.26u m=1
M31 N_16 N_9 N_14 VDD mp15  l=0.13u w=0.4u m=1
M32 N_70 N_19 VDD VDD mp15  l=0.13u w=0.4u m=1
M33 VDD N_19 N_70 VDD mp15  l=0.13u w=0.4u m=1
M34 N_74 N_5 N_14 VDD mp15  l=0.13u w=0.26u m=1
M35 Q N_18 VDD VDD mp15  l=0.13u w=0.4u m=1
M36 QN N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M37 VDDG N_29 N_75 VDDG mp15  l=0.13u w=0.26u m=1
M38 N_24 RETN N_75 VDDG mp15  l=0.13u w=0.26u m=1
M39 N_24 N_30 N_18 VDDG mp15  l=0.13u w=0.26u m=1
M40 N_30 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M41 N_29 N_24 VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends drfcrb0
* SPICE INPUT		Tue Sep 18 13:23:14 2018	drfcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfcrb1
.subckt drfcrb1 VDD VDDG GND Q QN RETN RN D CK
M1 GND N_9 N_5 GND mn15  l=0.13u w=0.2u m=1
M2 GND CK N_9 GND mn15  l=0.13u w=0.22u m=1
M3 N_41 D GND GND mn15  l=0.13u w=0.44u m=1
M4 N_41 N_9 N_11 GND mn15  l=0.13u w=0.44u m=1
M5 N_11 N_5 N_36 GND mn15  l=0.13u w=0.26u m=1
M6 GND N_15 N_36 GND mn15  l=0.13u w=0.26u m=1
M7 N_15 N_11 GND GND mn15  l=0.13u w=0.4u m=1
M8 GND N_19 N_13 GND mn15  l=0.13u w=0.4u m=1
M9 N_13 N_5 N_15 GND mn15  l=0.13u w=0.4u m=1
M10 N_19 RN GND GND mn15  l=0.13u w=0.3u m=1
M11 N_18 N_13 GND GND mn15  l=0.13u w=0.4u m=1
M12 N_13 N_9 N_50 GND mn15  l=0.13u w=0.26u m=1
M13 N_50 N_27 GND GND mn15  l=0.13u w=0.26u m=1
M14 Q N_18 GND GND mn15  l=0.13u w=0.46u m=1
M15 QN N_13 GND GND mn15  l=0.13u w=0.46u m=1
M16 N_27 RETN N_18 GND mn15  l=0.13u w=0.26u m=1
M17 N_30 RETN GND GND mn15  l=0.13u w=0.26u m=1
M18 N_29 N_27 GND GND mn15  l=0.13u w=0.26u m=1
M19 N_27 N_30 N_60 GND mn15  l=0.13u w=0.26u m=1
M20 GND N_29 N_60 GND mn15  l=0.13u w=0.26u m=1
M21 VDD N_9 N_5 VDD mp15  l=0.13u w=0.51u m=1
M22 VDD CK N_9 VDD mp15  l=0.13u w=0.56u m=1
M23 N_77 D VDD VDD mp15  l=0.13u w=0.6u m=1
M24 N_77 N_5 N_11 VDD mp15  l=0.13u w=0.6u m=1
M25 VDD N_15 N_76 VDD mp15  l=0.13u w=0.26u m=1
M26 N_11 N_9 N_76 VDD mp15  l=0.13u w=0.26u m=1
M27 N_19 RN VDD VDD mp15  l=0.13u w=0.5u m=1
M28 N_18 N_13 VDD VDD mp15  l=0.13u w=0.6u m=1
M29 N_15 N_9 N_13 VDD mp15  l=0.13u w=0.6u m=1
M30 N_66 N_11 N_15 VDD mp15  l=0.13u w=0.6u m=1
M31 N_66 N_19 VDD VDD mp15  l=0.13u w=0.6u m=1
M32 VDD N_19 N_66 VDD mp15  l=0.13u w=0.6u m=1
M33 N_78 N_5 N_13 VDD mp15  l=0.13u w=0.26u m=1
M34 N_78 N_27 N_66 VDD mp15  l=0.13u w=0.26u m=1
M35 Q N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 QN N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M37 N_30 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M38 N_29 N_27 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M39 N_27 N_30 N_18 VDDG mp15  l=0.13u w=0.26u m=1
M40 N_27 RETN N_79 VDDG mp15  l=0.13u w=0.26u m=1
M41 VDDG N_29 N_79 VDDG mp15  l=0.13u w=0.26u m=1
.ends drfcrb1
* SPICE INPUT		Tue Sep 18 13:23:21 2018	drfcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfcrb2
.subckt drfcrb2 VDD VDDG GND QN Q RETN RN D CK
M1 N_7 CK GND GND mn15  l=0.13u w=0.28u m=1
M2 GND N_7 N_5 GND mn15  l=0.13u w=0.22u m=1
M3 N_9 RN GND GND mn15  l=0.13u w=0.2u m=1
M4 GND RN N_9 GND mn15  l=0.13u w=0.2u m=1
M5 N_12 N_5 N_11 GND mn15  l=0.13u w=0.46u m=1
M6 N_48 N_5 N_14 GND mn15  l=0.13u w=0.26u m=1
M7 GND N_11 N_48 GND mn15  l=0.13u w=0.26u m=1
M8 GND N_14 N_11 GND mn15  l=0.13u w=0.46u m=1
M9 N_47 N_7 N_14 GND mn15  l=0.13u w=0.46u m=1
M10 N_47 D GND GND mn15  l=0.13u w=0.46u m=1
M11 QN N_12 GND GND mn15  l=0.13u w=0.46u m=1
M12 GND N_12 QN GND mn15  l=0.13u w=0.46u m=1
M13 GND N_9 N_12 GND mn15  l=0.13u w=0.46u m=1
M14 GND N_26 Q GND mn15  l=0.13u w=0.46u m=1
M15 GND N_26 Q GND mn15  l=0.13u w=0.46u m=1
M16 N_61 N_7 N_12 GND mn15  l=0.13u w=0.26u m=1
M17 GND N_27 N_61 GND mn15  l=0.13u w=0.26u m=1
M18 GND N_12 N_26 GND mn15  l=0.13u w=0.46u m=1
M19 N_27 RETN N_26 GND mn15  l=0.13u w=0.26u m=1
M20 N_33 RETN GND GND mn15  l=0.13u w=0.26u m=1
M21 N_32 N_27 GND GND mn15  l=0.13u w=0.26u m=1
M22 GND N_32 N_66 GND mn15  l=0.13u w=0.26u m=1
M23 N_27 N_33 N_66 GND mn15  l=0.13u w=0.26u m=1
M24 N_74 D VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_7 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD N_7 N_5 VDD mp15  l=0.13u w=0.56u m=1
M27 N_74 N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_11 N_77 VDD mp15  l=0.13u w=0.26u m=1
M29 N_14 N_7 N_77 VDD mp15  l=0.13u w=0.26u m=1
M30 N_9 RN VDD VDD mp15  l=0.13u w=0.3u m=1
M31 N_9 RN VDD VDD mp15  l=0.13u w=0.3u m=1
M32 N_11 N_14 N_70 VDD mp15  l=0.13u w=0.69u m=1
M33 N_11 N_7 N_12 VDD mp15  l=0.13u w=0.69u m=1
M34 VDD N_9 N_70 VDD mp15  l=0.13u w=0.69u m=1
M35 N_70 N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 N_12 N_5 N_78 VDD mp15  l=0.13u w=0.26u m=1
M37 N_70 N_27 N_78 VDD mp15  l=0.13u w=0.26u m=1
M38 QN N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 VDD N_12 QN VDD mp15  l=0.13u w=0.69u m=1
M40 Q N_26 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 Q N_26 VDD VDD mp15  l=0.13u w=0.69u m=1
M42 N_26 N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M43 N_33 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M44 N_32 N_27 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M45 N_27 RETN N_79 VDDG mp15  l=0.13u w=0.26u m=1
M46 VDDG N_32 N_79 VDDG mp15  l=0.13u w=0.26u m=1
M47 N_27 N_33 N_26 VDDG mp15  l=0.13u w=0.26u m=1
.ends drfcrb2
* SPICE INPUT		Tue Sep 18 13:23:27 2018	drfcrbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfcrbm
.subckt drfcrbm VDD VDDG GND Q QN RETN RN D CK
M1 GND N_9 N_5 GND mn15  l=0.13u w=0.2u m=1
M2 GND CK N_9 GND mn15  l=0.13u w=0.22u m=1
M3 N_41 D GND GND mn15  l=0.13u w=0.32u m=1
M4 N_41 N_9 N_11 GND mn15  l=0.13u w=0.32u m=1
M5 N_11 N_5 N_36 GND mn15  l=0.13u w=0.26u m=1
M6 GND N_16 N_36 GND mn15  l=0.13u w=0.26u m=1
M7 N_16 N_11 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_16 N_5 N_14 GND mn15  l=0.13u w=0.26u m=1
M9 N_14 N_19 GND GND mn15  l=0.13u w=0.26u m=1
M10 N_19 RN GND GND mn15  l=0.13u w=0.26u m=1
M11 N_18 N_14 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_14 N_9 N_50 GND mn15  l=0.13u w=0.26u m=1
M13 N_50 N_27 GND GND mn15  l=0.13u w=0.26u m=1
M14 Q N_18 GND GND mn15  l=0.13u w=0.36u m=1
M15 QN N_14 GND GND mn15  l=0.13u w=0.36u m=1
M16 N_27 RETN N_18 GND mn15  l=0.13u w=0.26u m=1
M17 N_30 RETN GND GND mn15  l=0.13u w=0.26u m=1
M18 N_29 N_27 GND GND mn15  l=0.13u w=0.26u m=1
M19 N_27 N_30 N_60 GND mn15  l=0.13u w=0.26u m=1
M20 GND N_29 N_60 GND mn15  l=0.13u w=0.26u m=1
M21 VDD N_9 N_5 VDD mp15  l=0.13u w=0.51u m=1
M22 N_9 CK VDD VDD mp15  l=0.13u w=0.56u m=1
M23 N_73 D VDD VDD mp15  l=0.13u w=0.4u m=1
M24 N_73 N_5 N_11 VDD mp15  l=0.13u w=0.4u m=1
M25 VDD N_16 N_72 VDD mp15  l=0.13u w=0.26u m=1
M26 N_11 N_9 N_72 VDD mp15  l=0.13u w=0.26u m=1
M27 N_19 RN VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_18 N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M29 N_16 N_9 N_14 VDD mp15  l=0.13u w=0.4u m=1
M30 N_16 N_11 N_66 VDD mp15  l=0.13u w=0.4u m=1
M31 N_74 N_5 N_14 VDD mp15  l=0.13u w=0.26u m=1
M32 N_74 N_27 N_66 VDD mp15  l=0.13u w=0.26u m=1
M33 N_66 N_19 VDD VDD mp15  l=0.13u w=0.4u m=1
M34 VDD N_19 N_66 VDD mp15  l=0.13u w=0.4u m=1
M35 Q N_18 VDD VDD mp15  l=0.13u w=0.55u m=1
M36 QN N_14 VDD VDD mp15  l=0.13u w=0.55u m=1
M37 N_30 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M38 N_29 N_27 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M39 N_27 N_30 N_18 VDDG mp15  l=0.13u w=0.26u m=1
M40 N_27 RETN N_75 VDDG mp15  l=0.13u w=0.26u m=1
M41 VDDG N_29 N_75 VDDG mp15  l=0.13u w=0.26u m=1
.ends drfcrbm
* SPICE INPUT		Tue Sep 18 13:23:33 2018	drfnrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfnrb0
.subckt drfnrb0 VDD VDDG GND QN Q RETN CK D
M1 N_34 N_18 N_7 GND mn15  l=0.13u w=0.26u m=1
M2 N_34 N_5 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_7 N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_38 N_9 N_7 GND mn15  l=0.13u w=0.28u m=1
M5 N_38 D GND GND mn15  l=0.13u w=0.28u m=1
M6 GND CK N_9 GND mn15  l=0.13u w=0.22u m=1
M7 QN N_14 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_14 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M9 GND N_9 N_18 GND mn15  l=0.13u w=0.2u m=1
M10 GND N_5 N_42 GND mn15  l=0.13u w=0.39u m=1
M11 N_17 N_18 N_42 GND mn15  l=0.13u w=0.39u m=1
M12 Q N_17 GND GND mn15  l=0.13u w=0.26u m=1
M13 N_51 N_9 N_17 GND mn15  l=0.13u w=0.26u m=1
M14 N_51 N_26 GND GND mn15  l=0.13u w=0.26u m=1
M15 N_23 RETN GND GND mn15  l=0.13u w=0.26u m=1
M16 GND N_26 N_28 GND mn15  l=0.13u w=0.26u m=1
M17 N_56 N_28 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_14 RETN N_26 GND mn15  l=0.13u w=0.26u m=1
M19 N_56 N_23 N_26 GND mn15  l=0.13u w=0.26u m=1
M20 N_126 N_18 N_7 VDD mp15  l=0.13u w=0.42u m=1
M21 N_127 N_9 N_7 VDD mp15  l=0.13u w=0.26u m=1
M22 N_126 D VDD VDD mp15  l=0.13u w=0.42u m=1
M23 N_127 N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
M24 N_9 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M25 N_5 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M26 QN N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M27 N_14 N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 VDD N_9 N_18 VDD mp15  l=0.13u w=0.49u m=1
M29 VDD N_5 N_128 VDD mp15  l=0.13u w=0.58u m=1
M30 N_128 N_9 N_17 VDD mp15  l=0.13u w=0.58u m=1
M31 Q N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M32 N_17 N_18 N_129 VDDG mp15  l=0.13u w=0.26u m=1
M33 VDD N_26 N_129 VDDG mp15  l=0.13u w=0.26u m=1
M34 VDDG N_26 N_28 VDDG mp15  l=0.13u w=0.26u m=1
M35 N_130 N_28 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M36 N_130 RETN N_26 VDDG mp15  l=0.13u w=0.26u m=1
M37 N_14 N_23 N_26 VDDG mp15  l=0.13u w=0.26u m=1
M38 N_23 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends drfnrb0
* SPICE INPUT		Tue Sep 18 13:23:39 2018	drfnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfnrb1
.subckt drfnrb1 VDDG VDD GND QN Q RETN CK D
M1 N_34 N_5 N_7 GND mn15  l=0.13u w=0.4u m=1
M2 N_34 D GND GND mn15  l=0.13u w=0.4u m=1
M3 GND CK N_5 GND mn15  l=0.13u w=0.22u m=1
M4 N_38 N_18 N_7 GND mn15  l=0.13u w=0.26u m=1
M5 N_38 N_9 GND GND mn15  l=0.13u w=0.26u m=1
M6 GND N_7 N_9 GND mn15  l=0.13u w=0.4u m=1
M7 QN N_14 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_14 N_17 GND GND mn15  l=0.13u w=0.4u m=1
M9 GND N_5 N_18 GND mn15  l=0.13u w=0.2u m=1
M10 GND N_9 N_42 GND mn15  l=0.13u w=0.46u m=1
M11 N_17 N_18 N_42 GND mn15  l=0.13u w=0.46u m=1
M12 Q N_17 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_51 N_5 N_17 GND mn15  l=0.13u w=0.26u m=1
M14 N_51 N_26 GND GND mn15  l=0.13u w=0.26u m=1
M15 N_23 RETN GND GND mn15  l=0.13u w=0.26u m=1
M16 N_56 N_23 N_26 GND mn15  l=0.13u w=0.26u m=1
M17 GND N_26 N_28 GND mn15  l=0.13u w=0.26u m=1
M18 N_56 N_28 GND GND mn15  l=0.13u w=0.26u m=1
M19 N_14 RETN N_26 GND mn15  l=0.13u w=0.26u m=1
M20 N_64 N_18 N_7 VDD mp15  l=0.13u w=0.6u m=1
M21 N_65 N_5 N_7 VDD mp15  l=0.13u w=0.26u m=1
M22 N_64 D VDD VDD mp15  l=0.13u w=0.6u m=1
M23 N_65 N_9 VDD VDD mp15  l=0.13u w=0.26u m=1
M24 N_5 CK VDD VDD mp15  l=0.13u w=0.56u m=1
M25 VDD N_7 N_9 VDD mp15  l=0.13u w=0.6u m=1
M26 N_18 N_5 VDD VDD mp15  l=0.13u w=0.51u m=1
M27 VDD N_14 QN VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_9 N_66 VDD mp15  l=0.13u w=0.69u m=1
M29 N_66 N_5 N_17 VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_17 N_14 VDD mp15  l=0.13u w=0.6u m=1
M31 VDD N_17 Q VDD mp15  l=0.13u w=0.69u m=1
M32 N_17 N_18 N_67 VDDG mp15  l=0.13u w=0.26u m=1
M33 VDD N_26 N_67 VDDG mp15  l=0.13u w=0.26u m=1
M34 N_14 N_23 N_26 VDDG mp15  l=0.13u w=0.26u m=1
M35 VDDG N_26 N_28 VDDG mp15  l=0.13u w=0.26u m=1
M36 N_68 N_28 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M37 N_68 RETN N_26 VDDG mp15  l=0.13u w=0.26u m=1
M38 N_23 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends drfnrb1
* SPICE INPUT		Tue Sep 18 13:23:46 2018	drfnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfnrb2
.subckt drfnrb2 VDDG VDD GND QN Q RETN CK D
M1 N_36 N_24 N_7 GND mn15  l=0.13u w=0.26u m=1
M2 N_36 N_5 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_7 N_5 GND mn15  l=0.13u w=0.4u m=1
M4 N_40 N_10 N_7 GND mn15  l=0.13u w=0.46u m=1
M5 N_40 D GND GND mn15  l=0.13u w=0.46u m=1
M6 N_10 CK GND GND mn15  l=0.13u w=0.28u m=1
M7 QN N_14 GND GND mn15  l=0.13u w=0.46u m=1
M8 QN N_14 GND GND mn15  l=0.13u w=0.46u m=1
M9 N_14 N_23 GND GND mn15  l=0.13u w=0.46u m=1
M10 GND N_17 N_19 GND mn15  l=0.13u w=0.26u m=1
M11 N_49 N_19 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_14 RETN N_17 GND mn15  l=0.13u w=0.26u m=1
M13 N_49 N_30 N_17 GND mn15  l=0.13u w=0.26u m=1
M14 GND N_10 N_24 GND mn15  l=0.13u w=0.22u m=1
M15 GND N_5 N_50 GND mn15  l=0.13u w=0.46u m=1
M16 N_23 N_24 N_50 GND mn15  l=0.13u w=0.46u m=1
M17 GND N_23 Q GND mn15  l=0.13u w=0.46u m=1
M18 GND N_23 Q GND mn15  l=0.13u w=0.46u m=1
M19 N_60 N_10 N_23 GND mn15  l=0.13u w=0.26u m=1
M20 N_60 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M21 N_30 RETN GND GND mn15  l=0.13u w=0.26u m=1
M22 N_136 N_24 N_7 VDD mp15  l=0.13u w=0.69u m=1
M23 N_137 N_10 N_7 VDD mp15  l=0.13u w=0.26u m=1
M24 N_136 D VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_137 N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
M26 VDD CK N_10 VDD mp15  l=0.13u w=0.69u m=1
M27 N_5 N_7 VDD VDD mp15  l=0.13u w=0.6u m=1
M28 QN N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 QN N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_23 N_14 VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_10 N_24 VDD mp15  l=0.13u w=0.56u m=1
M32 VDD N_5 N_138 VDD mp15  l=0.13u w=0.69u m=1
M33 N_23 N_10 N_138 VDD mp15  l=0.13u w=0.69u m=1
M34 Q N_23 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_23 Q VDD mp15  l=0.13u w=0.69u m=1
M36 N_23 N_24 N_139 VDDG mp15  l=0.13u w=0.26u m=1
M37 VDD N_17 N_139 VDDG mp15  l=0.13u w=0.26u m=1
M38 VDDG N_17 N_19 VDDG mp15  l=0.13u w=0.26u m=1
M39 N_140 N_19 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M40 N_140 RETN N_17 VDDG mp15  l=0.13u w=0.26u m=1
M41 N_14 N_30 N_17 VDDG mp15  l=0.13u w=0.26u m=1
M42 N_30 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends drfnrb2
* SPICE INPUT		Tue Sep 18 13:23:53 2018	drfnrbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfnrbm
.subckt drfnrbm VDD VDDG GND QN Q RETN CK D
M1 N_34 N_18 N_7 GND mn15  l=0.13u w=0.26u m=1
M2 N_34 N_5 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_7 N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_38 N_9 N_7 GND mn15  l=0.13u w=0.28u m=1
M5 N_38 D GND GND mn15  l=0.13u w=0.28u m=1
M6 GND CK N_9 GND mn15  l=0.13u w=0.22u m=1
M7 QN N_14 GND GND mn15  l=0.13u w=0.36u m=1
M8 N_14 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M9 GND N_9 N_18 GND mn15  l=0.13u w=0.2u m=1
M10 GND N_5 N_42 GND mn15  l=0.13u w=0.4u m=1
M11 N_17 N_18 N_42 GND mn15  l=0.13u w=0.4u m=1
M12 Q N_17 GND GND mn15  l=0.13u w=0.36u m=1
M13 N_51 N_9 N_17 GND mn15  l=0.13u w=0.26u m=1
M14 N_51 N_26 GND GND mn15  l=0.13u w=0.26u m=1
M15 N_23 RETN GND GND mn15  l=0.13u w=0.26u m=1
M16 GND N_26 N_28 GND mn15  l=0.13u w=0.26u m=1
M17 N_56 N_28 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_14 RETN N_26 GND mn15  l=0.13u w=0.26u m=1
M19 N_56 N_23 N_26 GND mn15  l=0.13u w=0.26u m=1
M20 N_126 N_18 N_7 VDD mp15  l=0.13u w=0.42u m=1
M21 N_127 N_9 N_7 VDD mp15  l=0.13u w=0.26u m=1
M22 N_126 D VDD VDD mp15  l=0.13u w=0.42u m=1
M23 N_127 N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
M24 N_9 CK VDD VDD mp15  l=0.13u w=0.56u m=1
M25 N_5 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M26 QN N_14 VDD VDD mp15  l=0.13u w=0.55u m=1
M27 N_14 N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 VDD N_9 N_18 VDD mp15  l=0.13u w=0.51u m=1
M29 VDD N_5 N_128 VDD mp15  l=0.13u w=0.6u m=1
M30 N_128 N_9 N_17 VDD mp15  l=0.13u w=0.6u m=1
M31 Q N_17 VDD VDD mp15  l=0.13u w=0.55u m=1
M32 N_17 N_18 N_129 VDDG mp15  l=0.13u w=0.26u m=1
M33 VDD N_26 N_129 VDDG mp15  l=0.13u w=0.26u m=1
M34 VDDG N_26 N_28 VDDG mp15  l=0.13u w=0.26u m=1
M35 N_130 N_28 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M36 N_130 RETN N_26 VDDG mp15  l=0.13u w=0.26u m=1
M37 N_14 N_23 N_26 VDDG mp15  l=0.13u w=0.26u m=1
M38 N_23 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends drfnrbm
* SPICE INPUT		Tue Sep 18 13:23:59 2018	drfprb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfprb0
.subckt drfprb0 VDDG VDD GND Q QN RETN SN CK D
M1 N_7 CK GND GND mn15  l=0.13u w=0.21u m=1
M2 GND N_7 N_5 GND mn15  l=0.13u w=0.19u m=1
M3 N_40 D GND GND mn15  l=0.13u w=0.28u m=1
M4 N_12 N_7 N_40 GND mn15  l=0.13u w=0.28u m=1
M5 N_38 N_18 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_12 N_5 N_38 GND mn15  l=0.13u w=0.26u m=1
M7 N_14 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_16 N_12 N_18 GND mn15  l=0.13u w=0.3u m=1
M9 N_16 SN GND GND mn15  l=0.13u w=0.3u m=1
M10 N_16 SN GND GND mn15  l=0.13u w=0.3u m=1
M11 N_18 N_5 N_17 GND mn15  l=0.13u w=0.26u m=1
M12 Q N_14 GND GND mn15  l=0.13u w=0.26u m=1
M13 QN N_17 GND GND mn15  l=0.13u w=0.26u m=1
M14 N_17 N_7 N_52 GND mn15  l=0.13u w=0.26u m=1
M15 N_16 N_27 N_52 GND mn15  l=0.13u w=0.26u m=1
M16 N_27 RETN N_14 GND mn15  l=0.13u w=0.26u m=1
M17 N_30 RETN GND GND mn15  l=0.13u w=0.26u m=1
M18 N_29 N_27 GND GND mn15  l=0.13u w=0.26u m=1
M19 N_27 N_30 N_60 GND mn15  l=0.13u w=0.26u m=1
M20 GND N_29 N_60 GND mn15  l=0.13u w=0.26u m=1
M21 N_7 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M22 VDD N_7 N_5 VDD mp15  l=0.13u w=0.49u m=1
M23 N_73 D VDD VDD mp15  l=0.13u w=0.42u m=1
M24 N_74 N_18 VDD VDD mp15  l=0.13u w=0.26u m=1
M25 N_73 N_5 N_12 VDD mp15  l=0.13u w=0.42u m=1
M26 N_74 N_7 N_12 VDD mp15  l=0.13u w=0.26u m=1
M27 N_14 N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_17 N_7 N_18 VDD mp15  l=0.13u w=0.4u m=1
M29 VDD N_12 N_18 VDD mp15  l=0.13u w=0.4u m=1
M30 N_17 SN VDD VDD mp15  l=0.13u w=0.4u m=1
M31 N_75 N_5 N_17 VDD mp15  l=0.13u w=0.26u m=1
M32 N_75 N_27 VDD VDD mp15  l=0.13u w=0.26u m=1
M33 Q N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M34 QN N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M35 N_27 N_30 N_14 VDDG mp15  l=0.13u w=0.26u m=1
M36 N_27 RETN N_76 VDDG mp15  l=0.13u w=0.26u m=1
M37 VDDG N_29 N_76 VDDG mp15  l=0.13u w=0.26u m=1
M38 N_30 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M39 N_29 N_27 VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends drfprb0
* SPICE INPUT		Tue Sep 18 13:24:05 2018	drfprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfprb1
.subckt drfprb1 VDDG VDD GND Q QN RETN SN CK D
M1 N_7 CK GND GND mn15  l=0.13u w=0.22u m=1
M2 GND N_7 N_5 GND mn15  l=0.13u w=0.19u m=1
M3 N_41 D GND GND mn15  l=0.13u w=0.39u m=1
M4 N_41 N_7 N_11 GND mn15  l=0.13u w=0.39u m=1
M5 N_38 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_11 N_5 N_38 GND mn15  l=0.13u w=0.26u m=1
M7 N_14 N_16 GND GND mn15  l=0.13u w=0.39u m=1
M8 N_15 N_11 N_17 GND mn15  l=0.13u w=0.4u m=1
M9 GND SN N_15 GND mn15  l=0.13u w=0.4u m=1
M10 N_15 SN GND GND mn15  l=0.13u w=0.4u m=1
M11 N_17 N_5 N_16 GND mn15  l=0.13u w=0.39u m=1
M12 QN N_16 GND GND mn15  l=0.13u w=0.46u m=1
M13 Q N_14 GND GND mn15  l=0.13u w=0.46u m=1
M14 N_16 N_7 N_52 GND mn15  l=0.13u w=0.26u m=1
M15 N_15 N_28 N_52 GND mn15  l=0.13u w=0.26u m=1
M16 N_28 N_33 N_55 GND mn15  l=0.13u w=0.26u m=1
M17 GND N_32 N_55 GND mn15  l=0.13u w=0.26u m=1
M18 N_28 RETN N_14 GND mn15  l=0.13u w=0.26u m=1
M19 N_33 RETN GND GND mn15  l=0.13u w=0.26u m=1
M20 N_32 N_28 GND GND mn15  l=0.13u w=0.26u m=1
M21 N_7 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M22 VDD N_7 N_5 VDD mp15  l=0.13u w=0.49u m=1
M23 N_73 D VDD VDD mp15  l=0.13u w=0.58u m=1
M24 N_74 N_17 VDD VDD mp15  l=0.13u w=0.26u m=1
M25 N_73 N_5 N_11 VDD mp15  l=0.13u w=0.58u m=1
M26 N_74 N_7 N_11 VDD mp15  l=0.13u w=0.26u m=1
M27 N_17 N_7 N_16 VDD mp15  l=0.13u w=0.58u m=1
M28 N_17 N_11 VDD VDD mp15  l=0.13u w=0.58u m=1
M29 N_16 SN VDD VDD mp15  l=0.13u w=0.58u m=1
M30 N_14 N_16 VDD VDD mp15  l=0.13u w=0.58u m=1
M31 N_16 N_5 N_75 VDD mp15  l=0.13u w=0.26u m=1
M32 N_75 N_28 VDD VDD mp15  l=0.13u w=0.26u m=1
M33 QN N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M34 Q N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 N_33 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M36 N_32 N_28 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M37 N_28 N_33 N_14 VDDG mp15  l=0.13u w=0.26u m=1
M38 N_28 RETN N_76 VDDG mp15  l=0.13u w=0.26u m=1
M39 VDDG N_32 N_76 VDDG mp15  l=0.13u w=0.26u m=1
.ends drfprb1
* SPICE INPUT		Tue Sep 18 13:24:11 2018	drfprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfprb2
.subckt drfprb2 VDDG VDD GND Q QN RETN SN CK D
M1 N_7 CK GND GND mn15  l=0.13u w=0.28u m=1
M2 GND N_7 N_5 GND mn15  l=0.13u w=0.22u m=1
M3 N_42 D GND GND mn15  l=0.13u w=0.46u m=1
M4 N_42 N_7 N_11 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_16 N_38 GND mn15  l=0.13u w=0.26u m=1
M6 N_11 N_5 N_38 GND mn15  l=0.13u w=0.26u m=1
M7 N_14 N_11 N_16 GND mn15  l=0.13u w=0.46u m=1
M8 N_14 SN GND GND mn15  l=0.13u w=0.46u m=1
M9 N_14 SN GND GND mn15  l=0.13u w=0.46u m=1
M10 N_16 N_5 N_15 GND mn15  l=0.13u w=0.46u m=1
M11 GND N_15 QN GND mn15  l=0.13u w=0.46u m=1
M12 QN N_15 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_15 N_20 GND mn15  l=0.13u w=0.46u m=1
M14 GND N_20 Q GND mn15  l=0.13u w=0.46u m=1
M15 GND N_20 Q GND mn15  l=0.13u w=0.46u m=1
M16 N_26 N_29 N_54 GND mn15  l=0.13u w=0.26u m=1
M17 GND N_28 N_54 GND mn15  l=0.13u w=0.26u m=1
M18 N_29 RETN GND GND mn15  l=0.13u w=0.26u m=1
M19 N_28 N_26 GND GND mn15  l=0.13u w=0.26u m=1
M20 N_26 RETN N_20 GND mn15  l=0.13u w=0.26u m=1
M21 N_15 N_7 N_62 GND mn15  l=0.13u w=0.26u m=1
M22 N_14 N_26 N_62 GND mn15  l=0.13u w=0.26u m=1
M23 N_7 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_7 N_5 VDD mp15  l=0.13u w=0.54u m=1
M25 N_71 D VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_72 N_16 VDD VDD mp15  l=0.13u w=0.26u m=1
M27 N_71 N_5 N_11 VDD mp15  l=0.13u w=0.69u m=1
M28 N_72 N_7 N_11 VDD mp15  l=0.13u w=0.26u m=1
M29 N_15 N_7 N_16 VDD mp15  l=0.13u w=0.69u m=1
M30 N_16 N_11 VDD VDD mp15  l=0.13u w=0.35u m=1
M31 N_16 N_11 VDD VDD mp15  l=0.13u w=0.34u m=1
M32 VDD N_15 QN VDD mp15  l=0.13u w=0.69u m=1
M33 QN N_15 VDD VDD mp15  l=0.13u w=0.69u m=1
M34 VDD N_15 N_20 VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_20 Q VDD mp15  l=0.13u w=0.69u m=1
M36 VDD N_20 Q VDD mp15  l=0.13u w=0.69u m=1
M37 N_15 SN VDD VDD mp15  l=0.13u w=0.34u m=1
M38 N_15 SN VDD VDD mp15  l=0.13u w=0.35u m=1
M39 N_15 N_5 N_73 VDD mp15  l=0.13u w=0.26u m=1
M40 N_73 N_26 VDD VDD mp15  l=0.13u w=0.26u m=1
M41 N_26 N_29 N_20 VDDG mp15  l=0.13u w=0.26u m=1
M42 N_26 RETN N_74 VDDG mp15  l=0.13u w=0.26u m=1
M43 VDDG N_28 N_74 VDDG mp15  l=0.13u w=0.26u m=1
M44 N_29 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M45 N_28 N_26 VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends drfprb2
* SPICE INPUT		Tue Sep 18 13:24:17 2018	drfprbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=drfprbm
.subckt drfprbm VDDG VDD GND Q QN RETN SN CK D
M1 N_7 CK GND GND mn15  l=0.13u w=0.21u m=1
M2 GND N_7 N_5 GND mn15  l=0.13u w=0.2u m=1
M3 N_40 D GND GND mn15  l=0.13u w=0.28u m=1
M4 N_12 N_7 N_40 GND mn15  l=0.13u w=0.28u m=1
M5 N_38 N_18 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_12 N_5 N_38 GND mn15  l=0.13u w=0.26u m=1
M7 N_14 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_16 N_12 N_18 GND mn15  l=0.13u w=0.3u m=1
M9 N_16 SN GND GND mn15  l=0.13u w=0.3u m=1
M10 N_16 SN GND GND mn15  l=0.13u w=0.3u m=1
M11 N_18 N_5 N_17 GND mn15  l=0.13u w=0.26u m=1
M12 Q N_14 GND GND mn15  l=0.13u w=0.35u m=1
M13 QN N_17 GND GND mn15  l=0.13u w=0.35u m=1
M14 N_17 N_7 N_52 GND mn15  l=0.13u w=0.26u m=1
M15 N_16 N_27 N_52 GND mn15  l=0.13u w=0.26u m=1
M16 N_27 RETN N_14 GND mn15  l=0.13u w=0.26u m=1
M17 N_30 RETN GND GND mn15  l=0.13u w=0.26u m=1
M18 N_29 N_27 GND GND mn15  l=0.13u w=0.26u m=1
M19 N_27 N_30 N_60 GND mn15  l=0.13u w=0.26u m=1
M20 GND N_29 N_60 GND mn15  l=0.13u w=0.26u m=1
M21 N_7 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M22 VDD N_7 N_5 VDD mp15  l=0.13u w=0.49u m=1
M23 N_73 D VDD VDD mp15  l=0.13u w=0.42u m=1
M24 N_74 N_18 VDD VDD mp15  l=0.13u w=0.26u m=1
M25 N_73 N_5 N_12 VDD mp15  l=0.13u w=0.42u m=1
M26 N_74 N_7 N_12 VDD mp15  l=0.13u w=0.26u m=1
M27 N_14 N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_17 N_7 N_18 VDD mp15  l=0.13u w=0.4u m=1
M29 VDD N_12 N_18 VDD mp15  l=0.13u w=0.4u m=1
M30 N_17 SN VDD VDD mp15  l=0.13u w=0.4u m=1
M31 N_75 N_5 N_17 VDD mp15  l=0.13u w=0.26u m=1
M32 N_75 N_27 VDD VDD mp15  l=0.13u w=0.26u m=1
M33 Q N_14 VDD VDD mp15  l=0.13u w=0.53u m=1
M34 QN N_17 VDD VDD mp15  l=0.13u w=0.53u m=1
M35 N_27 N_30 N_14 VDDG mp15  l=0.13u w=0.26u m=1
M36 N_27 RETN N_76 VDDG mp15  l=0.13u w=0.26u m=1
M37 VDDG N_29 N_76 VDDG mp15  l=0.13u w=0.26u m=1
M38 N_30 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M39 N_29 N_27 VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends drfprbm
* SPICE INPUT		Tue Sep 18 13:24:23 2018	gpgbuffd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpgbuffd16
.subckt gpgbuffd16 Y VDDG GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.72u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.72u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.72u m=1
M4 N_4 A GND GND mn15  l=0.13u w=0.72u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.84u m=1
M6 Y N_4 GND GND mn15  l=0.13u w=0.84u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.84u m=1
M8 Y N_4 GND GND mn15  l=0.13u w=0.84u m=1
M9 GND N_4 Y GND mn15  l=0.13u w=0.84u m=1
M10 Y N_4 GND GND mn15  l=0.13u w=0.84u m=1
M11 GND N_4 Y GND mn15  l=0.13u w=0.84u m=1
M12 Y N_4 GND GND mn15  l=0.13u w=0.72u m=1
M13 Y N_4 GND GND mn15  l=0.13u w=0.76u m=1
M14 VDDG A N_4 VDDG mp15  l=0.13u w=1.51u m=1
M15 VDDG A N_4 VDDG mp15  l=0.13u w=1.51u m=1
M16 VDDG A N_4 VDDG mp15  l=0.13u w=1.47u m=1
M17 VDDG N_4 Y VDDG mp15  l=0.13u w=1.47u m=1
M18 VDDG N_4 Y VDDG mp15  l=0.13u w=1.47u m=1
M19 VDDG N_4 Y VDDG mp15  l=0.13u w=1.47u m=1
M20 VDDG N_4 Y VDDG mp15  l=0.13u w=1.47u m=1
M21 Y N_4 VDDG VDDG mp15  l=0.13u w=1.33u m=1
M22 VDDG N_4 Y VDDG mp15  l=0.13u w=1.33u m=1
M23 Y N_4 VDDG VDDG mp15  l=0.13u w=1.33u m=1
M24 VDDG N_4 Y VDDG mp15  l=0.13u w=1.33u m=1
.ends gpgbuffd16
* SPICE INPUT		Tue Sep 18 13:24:29 2018	gpgbuffd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpgbuffd2
.subckt gpgbuffd2 VDDG Y GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 N_4 A VDDG VDDG mp15  l=0.13u w=0.56u m=1
M5 Y N_4 VDDG VDDG mp15  l=0.13u w=1.4u m=1
.ends gpgbuffd2
* SPICE INPUT		Tue Sep 18 13:24:36 2018	gpgbuffd32
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpgbuffd32
.subckt gpgbuffd32 Y VDDG GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.72u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.72u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.72u m=1
M4 N_4 A GND GND mn15  l=0.13u w=0.72u m=1
M5 GND A N_4 GND mn15  l=0.13u w=0.72u m=1
M6 N_4 A GND GND mn15  l=0.13u w=0.72u m=1
M7 GND A N_4 GND mn15  l=0.13u w=0.72u m=1
M8 N_4 A GND GND mn15  l=0.13u w=0.72u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.895u m=1
M10 Y N_4 GND GND mn15  l=0.13u w=0.895u m=1
M11 GND N_4 Y GND mn15  l=0.13u w=0.89u m=1
M12 Y N_4 GND GND mn15  l=0.13u w=0.89u m=1
M13 GND N_4 Y GND mn15  l=0.13u w=0.89u m=1
M14 Y N_4 GND GND mn15  l=0.13u w=0.89u m=1
M15 GND N_4 Y GND mn15  l=0.13u w=0.89u m=1
M16 Y N_4 GND GND mn15  l=0.13u w=0.89u m=1
M17 GND N_4 Y GND mn15  l=0.13u w=0.89u m=1
M18 Y N_4 GND GND mn15  l=0.13u w=0.89u m=1
M19 GND N_4 Y GND mn15  l=0.13u w=0.89u m=1
M20 Y N_4 GND GND mn15  l=0.13u w=0.89u m=1
M21 GND N_4 Y GND mn15  l=0.13u w=0.89u m=1
M22 Y N_4 GND GND mn15  l=0.13u w=0.89u m=1
M23 GND N_4 Y GND mn15  l=0.13u w=0.89u m=1
M24 Y N_4 GND GND mn15  l=0.13u w=0.89u m=1
M25 Y N_4 GND GND mn15  l=0.13u w=0.47u m=1
M26 VDDG A N_4 VDDG mp15  l=0.13u w=1.76u m=1
M27 VDDG A N_4 VDDG mp15  l=0.13u w=1.44u m=1
M28 N_4 A VDDG VDDG mp15  l=0.13u w=1.44u m=1
M29 VDDG A N_4 VDDG mp15  l=0.13u w=1.44u m=1
M30 N_4 A VDDG VDDG mp15  l=0.13u w=1.44u m=1
M31 VDDG A N_4 VDDG mp15  l=0.13u w=1.44u m=1
M32 Y N_4 VDDG VDDG mp15  l=0.13u w=1.68u m=1
M33 Y N_4 VDDG VDDG mp15  l=0.13u w=1.68u m=1
M34 VDDG N_4 Y VDDG mp15  l=0.13u w=1.68u m=1
M35 Y N_4 VDDG VDDG mp15  l=0.13u w=1.68u m=1
M36 VDDG N_4 Y VDDG mp15  l=0.13u w=1.74u m=1
M37 VDDG N_4 Y VDDG mp15  l=0.13u w=1.74u m=1
M38 VDDG N_4 Y VDDG mp15  l=0.13u w=1.74u m=1
M39 Y N_4 VDDG VDDG mp15  l=0.13u w=1.74u m=1
M40 VDDG N_4 Y VDDG mp15  l=0.13u w=1.74u m=1
M41 Y N_4 VDDG VDDG mp15  l=0.13u w=1.74u m=1
M42 VDDG N_4 Y VDDG mp15  l=0.13u w=1.32u m=1
M43 Y N_4 VDDG VDDG mp15  l=0.13u w=1.32u m=1
M44 VDDG N_4 Y VDDG mp15  l=0.13u w=1.32u m=1
M45 Y N_4 VDDG VDDG mp15  l=0.13u w=1.32u m=1
.ends gpgbuffd32
* SPICE INPUT		Tue Sep 18 13:24:42 2018	gpgbuffd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpgbuffd4
.subckt gpgbuffd4 Y VDDG GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.36u m=1
M3 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 VDDG A N_4 VDDG mp15  l=0.13u w=1.12u m=1
M8 VDDG N_4 Y VDDG mp15  l=0.13u w=1.4u m=1
M9 VDDG N_4 Y VDDG mp15  l=0.13u w=1.4u m=1
.ends gpgbuffd4
* SPICE INPUT		Tue Sep 18 13:24:48 2018	gpgbuffd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpgbuffd8
.subckt gpgbuffd8 Y VDDG GND VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.72u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.72u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 VDDG A N_5 VDDG mp15  l=0.13u w=1.12u m=1
M12 N_5 A VDDG VDDG mp15  l=0.13u w=1.12u m=1
M13 VDDG N_5 Y VDDG mp15  l=0.13u w=1.4u m=1
M14 VDDG N_5 Y VDDG mp15  l=0.13u w=1.4u m=1
M15 VDDG N_5 Y VDDG mp15  l=0.13u w=1.4u m=1
M16 Y N_5 VDDG VDDG mp15  l=0.13u w=1.4u m=1
.ends gpgbuffd8
* SPICE INPUT		Tue Sep 18 13:24:54 2018	gpginvd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpginvd16
.subckt gpginvd16 VDDG Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.735u m=1
M2 GND A Y GND mn15  l=0.13u w=0.735u m=1
M3 GND A Y GND mn15  l=0.13u w=0.735u m=1
M4 Y A GND GND mn15  l=0.13u w=0.735u m=1
M5 GND A Y GND mn15  l=0.13u w=0.735u m=1
M6 Y A GND GND mn15  l=0.13u w=0.735u m=1
M7 GND A Y GND mn15  l=0.13u w=0.735u m=1
M8 Y A GND GND mn15  l=0.13u w=0.735u m=1
M9 GND A Y GND mn15  l=0.13u w=0.735u m=1
M10 Y A GND GND mn15  l=0.13u w=0.735u m=1
M11 Y A VDDG VDDG mp15  l=0.13u w=1.87u m=1
M12 Y A VDDG VDDG mp15  l=0.13u w=1.87u m=1
M13 VDDG A Y VDDG mp15  l=0.13u w=1.87u m=1
M14 Y A VDDG VDDG mp15  l=0.13u w=1.87u m=1
M15 VDDG A Y VDDG mp15  l=0.13u w=1.87u m=1
M16 Y A VDDG VDDG mp15  l=0.13u w=1.85u m=1
.ends gpginvd16
* SPICE INPUT		Tue Sep 18 13:25:00 2018	gpginvd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpginvd2
.subckt gpginvd2 Y GND VDDG VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 Y A VDDG VDDG mp15  l=0.13u w=1.4u m=1
.ends gpginvd2
* SPICE INPUT		Tue Sep 18 13:25:06 2018	gpginvd32
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpginvd32
.subckt gpginvd32 Y GND VDD A VDDG
M1 Y A GND GND mn15  l=0.13u w=1.68u m=1
M2 Y A GND GND mn15  l=0.13u w=1.68u m=1
M3 Y A GND GND mn15  l=0.13u w=0.71u m=1
M4 Y A GND GND mn15  l=0.13u w=0.71u m=1
M5 GND A Y GND mn15  l=0.13u w=0.71u m=1
M6 Y A GND GND mn15  l=0.13u w=0.71u m=1
M7 GND A Y GND mn15  l=0.13u w=0.71u m=1
M8 Y A GND GND mn15  l=0.13u w=0.71u m=1
M9 GND A Y GND mn15  l=0.13u w=0.71u m=1
M10 Y A GND GND mn15  l=0.13u w=0.71u m=1
M11 GND A Y GND mn15  l=0.13u w=0.71u m=1
M12 Y A GND GND mn15  l=0.13u w=0.71u m=1
M13 GND A Y GND mn15  l=0.13u w=0.71u m=1
M14 Y A GND GND mn15  l=0.13u w=0.71u m=1
M15 GND A Y GND mn15  l=0.13u w=0.71u m=1
M16 Y A GND GND mn15  l=0.13u w=0.71u m=1
M17 GND A Y GND mn15  l=0.13u w=0.71u m=1
M18 Y A GND GND mn15  l=0.13u w=0.71u m=1
M19 Y A VDDG VDDG mp15  l=0.13u w=1.87u m=1
M20 Y A VDDG VDDG mp15  l=0.13u w=1.87u m=1
M21 VDDG A Y VDDG mp15  l=0.13u w=1.87u m=1
M22 Y A VDDG VDDG mp15  l=0.13u w=1.87u m=1
M23 VDDG A Y VDDG mp15  l=0.13u w=1.87u m=1
M24 Y A VDDG VDDG mp15  l=0.13u w=1.87u m=1
M25 VDDG A Y VDDG mp15  l=0.13u w=1.87u m=1
M26 Y A VDDG VDDG mp15  l=0.13u w=1.87u m=1
M27 VDDG A Y VDDG mp15  l=0.13u w=1.87u m=1
M28 Y A VDDG VDDG mp15  l=0.13u w=1.87u m=1
M29 VDDG A Y VDDG mp15  l=0.13u w=1.87u m=1
M30 Y A VDDG VDDG mp15  l=0.13u w=1.83u m=1
.ends gpginvd32
* SPICE INPUT		Tue Sep 18 13:25:12 2018	gpginvd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpginvd4
.subckt gpginvd4 Y VDDG GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 VDDG A Y VDDG mp15  l=0.13u w=1.4u m=1
M6 VDDG A Y VDDG mp15  l=0.13u w=1.4u m=1
.ends gpginvd4
* SPICE INPUT		Tue Sep 18 13:25:19 2018	gpginvd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=gpginvd8
.subckt gpginvd8 Y VDDG GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A Y GND mn15  l=0.13u w=0.46u m=1
M8 Y A GND GND mn15  l=0.13u w=0.46u m=1
M9 VDDG A Y VDDG mp15  l=0.13u w=1.87u m=1
M10 VDDG A Y VDDG mp15  l=0.13u w=1.87u m=1
M11 VDDG A Y VDDG mp15  l=0.13u w=1.86u m=1
.ends gpginvd8
* SPICE INPUT		Tue Sep 18 13:25:25 2018	head1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=head1
.subckt head1 GND SLEEPOUT VDDG VDD SLEEP
M1 N_4 SLEEP GND GND mn15  l=0.13u w=0.26u m=1
M2 SLEEPOUT N_4 GND GND mn15  l=0.13u w=0.52u m=1
M3 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2u m=1
M4 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2u m=1
M5 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2u m=1
M6 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2u m=1
M7 N_4 SLEEP VDDG VDDG mp15  l=0.13u w=0.4u m=1
M8 SLEEPOUT N_4 VDDG VDDG mp15  l=0.13u w=0.8u m=1
.ends head1
* SPICE INPUT		Tue Sep 18 13:25:31 2018	head2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=head2
.subckt head2 SLEEPOUT GND VDDG VDD SLEEP
M1 GND SLEEP N_4 GND mn15  l=0.13u w=0.4u m=1
M2 GND N_4 SLEEPOUT GND mn15  l=0.13u w=0.55u m=1
M3 GND N_4 SLEEPOUT GND mn15  l=0.13u w=0.55u m=1
M4 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2.4u m=1
M5 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2.4u m=1
M6 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2.4u m=1
M7 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2.4u m=1
M8 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2.4u m=1
M9 N_4 SLEEP VDDG VDDG mp15  l=0.13u w=0.6u m=1
M10 SLEEPOUT N_4 VDDG VDDG mp15  l=0.13u w=0.825u m=1
M11 VDDG N_4 SLEEPOUT VDDG mp15  l=0.13u w=0.825u m=1
.ends head2
* SPICE INPUT		Tue Sep 18 13:25:37 2018	head4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=head4
.subckt head4 GND SLEEPOUT VDDG VDD SLEEP
M1 N_5 SLEEP GND GND mn15  l=0.13u w=0.8u m=1
M2 SLEEPOUT N_5 GND GND mn15  l=0.13u w=0.8u m=1
M3 SLEEPOUT N_5 GND GND mn15  l=0.13u w=0.7u m=1
M4 SLEEPOUT N_5 GND GND mn15  l=0.13u w=0.7u m=1
M5 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2.4u m=1
M6 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2.4u m=1
M7 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2.4u m=1
M8 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2.4u m=1
M9 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2.4u m=1
M10 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2.4u m=1
M11 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2.4u m=1
M12 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2.4u m=1
M13 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2.4u m=1
M14 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2.4u m=1
M15 N_5 SLEEP VDDG VDDG mp15  l=0.13u w=1.2u m=1
M16 SLEEPOUT N_5 VDDG VDDG mp15  l=0.13u w=1.1u m=1
M17 SLEEPOUT N_5 VDDG VDDG mp15  l=0.13u w=1.1u m=1
M18 SLEEPOUT N_5 VDDG VDDG mp15  l=0.13u w=1.1u m=1
.ends head4
* SPICE INPUT		Tue Sep 18 13:25:43 2018	headm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=headm
.subckt headm GND SLEEPOUT VDDG VDD SLEEP
M1 N_4 SLEEP GND GND mn15  l=0.13u w=0.26u m=1
M2 SLEEPOUT N_4 GND GND mn15  l=0.13u w=0.52u m=1
M3 VDD SLEEP VDDG VDDG mp15  l=0.13u w=2u m=1
M4 VDDG SLEEP VDD VDDG mp15  l=0.13u w=2u m=1
M5 N_4 SLEEP VDDG VDDG mp15  l=0.13u w=0.4u m=1
M6 SLEEPOUT N_4 VDDG VDDG mp15  l=0.13u w=0.8u m=1
.ends headm
* SPICE INPUT		Tue Sep 18 13:25:49 2018	isohd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=isohd1
.subckt isohd1 GND Y EN A VDD
M1 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 EN GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_9 A N_5 VDD mp15  l=0.13u w=0.6u m=1
M5 N_9 EN VDD VDD mp15  l=0.13u w=0.6u m=1
M6 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends isohd1
* SPICE INPUT		Tue Sep 18 13:25:55 2018	isohd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=isohd2
.subckt isohd2 Y VDD GND EN A
M1 N_4 A GND GND mn15  l=0.13u w=0.36u m=1
M2 GND EN N_4 GND mn15  l=0.13u w=0.36u m=1
M3 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 N_6 A N_4 VDD mp15  l=0.13u w=0.69u m=1
M6 VDD EN N_6 VDD mp15  l=0.13u w=0.69u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends isohd2
* SPICE INPUT		Tue Sep 18 13:26:01 2018	isohd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=isohd4
.subckt isohd4 Y GND VDD EN A
M1 N_6 EN GND GND mn15  l=0.13u w=0.36u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.36u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.36u m=1
M4 N_6 EN GND GND mn15  l=0.13u w=0.36u m=1
M5 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M9 N_16 EN VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_17 A N_6 VDD mp15  l=0.13u w=0.69u m=1
M11 N_6 A N_16 VDD mp15  l=0.13u w=0.69u m=1
M12 N_17 EN VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends isohd4
* SPICE INPUT		Tue Sep 18 13:26:08 2018	isohdm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=isohdm
.subckt isohdm GND Y EN A VDD
M1 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 EN GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.33u m=1
M4 N_10 A N_5 VDD mp15  l=0.13u w=0.52u m=1
M5 N_10 EN VDD VDD mp15  l=0.13u w=0.52u m=1
M6 VDD N_5 Y VDD mp15  l=0.13u w=0.5u m=1
.ends isohdm
* SPICE INPUT		Tue Sep 18 13:26:14 2018	isold1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=isold1
.subckt isold1 GND Y VDD E A
M1 N_5 A N_4 GND mn15  l=0.13u w=0.33u m=1
M2 N_5 E GND GND mn15  l=0.13u w=0.33u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M5 N_4 E VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends isold1
* SPICE INPUT		Tue Sep 18 13:26:21 2018	isold2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=isold2
.subckt isold2 Y GND VDD E A
M1 N_6 A N_4 GND mn15  l=0.13u w=0.46u m=1
M2 GND E N_6 GND mn15  l=0.13u w=0.46u m=1
M3 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.6u m=1
M6 N_4 E VDD VDD mp15  l=0.13u w=0.6u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends isold2
* SPICE INPUT		Tue Sep 18 13:26:27 2018	isold4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=isold4
.subckt isold4 Y GND VDD E A
M1 N_9 E GND GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND E N_10 GND mn15  l=0.13u w=0.46u m=1
M7 N_10 A N_5 GND mn15  l=0.13u w=0.46u m=1
M8 N_5 A N_9 GND mn15  l=0.13u w=0.46u m=1
M9 N_5 E VDD VDD mp15  l=0.13u w=0.6u m=1
M10 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M13 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD E N_5 VDD mp15  l=0.13u w=0.6u m=1
M15 N_5 A VDD VDD mp15  l=0.13u w=0.6u m=1
M16 VDD A N_5 VDD mp15  l=0.13u w=0.6u m=1
.ends isold4
* SPICE INPUT		Tue Sep 18 13:26:33 2018	isoldm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=isoldm
.subckt isoldm GND Y VDD E A
M1 N_5 A N_4 GND mn15  l=0.13u w=0.26u m=1
M2 N_5 E GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.33u m=1
M4 N_4 A VDD VDD mp15  l=0.13u w=0.26u m=1
M5 N_4 E VDD VDD mp15  l=0.13u w=0.26u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
.ends isoldm
* SPICE INPUT		Tue Sep 18 13:28:46 2018	sdrcrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrcrb0
.subckt sdrcrb0 VDD VDDG GND Q QN RETN RN SI CK D SE
M1 GND SE N_5 GND mn15  l=0.13u w=0.26u m=1
M2 N_46 N_5 GND GND mn15  l=0.13u w=0.4u m=1
M3 N_46 D N_10 GND mn15  l=0.13u w=0.4u m=1
M4 N_10 SE N_43 GND mn15  l=0.13u w=0.26u m=1
M5 N_43 SI GND GND mn15  l=0.13u w=0.26u m=1
M6 N_14 CK GND GND mn15  l=0.13u w=0.21u m=1
M7 GND N_14 N_12 GND mn15  l=0.13u w=0.19u m=1
M8 N_10 N_14 N_17 GND mn15  l=0.13u w=0.4u m=1
M9 N_17 N_12 N_50 GND mn15  l=0.13u w=0.26u m=1
M10 GND N_21 N_50 GND mn15  l=0.13u w=0.26u m=1
M11 N_21 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M12 GND N_25 N_19 GND mn15  l=0.13u w=0.26u m=1
M13 N_19 N_12 N_21 GND mn15  l=0.13u w=0.26u m=1
M14 GND N_19 N_23 GND mn15  l=0.13u w=0.26u m=1
M15 N_25 RN GND GND mn15  l=0.13u w=0.26u m=1
M16 N_19 N_14 N_62 GND mn15  l=0.13u w=0.26u m=1
M17 N_62 N_33 GND GND mn15  l=0.13u w=0.26u m=1
M18 QN N_19 GND GND mn15  l=0.13u w=0.26u m=1
M19 Q N_23 GND GND mn15  l=0.13u w=0.26u m=1
M20 N_33 RETN N_23 GND mn15  l=0.13u w=0.26u m=1
M21 N_36 RETN GND GND mn15  l=0.13u w=0.26u m=1
M22 N_35 N_33 GND GND mn15  l=0.13u w=0.26u m=1
M23 N_33 N_36 N_72 GND mn15  l=0.13u w=0.26u m=1
M24 GND N_35 N_72 GND mn15  l=0.13u w=0.26u m=1
M25 VDD SE N_5 VDD mp15  l=0.13u w=0.39u m=1
M26 N_75 N_5 N_82 VDD mp15  l=0.13u w=0.26u m=1
M27 N_87 D N_75 VDD mp15  l=0.13u w=0.58u m=1
M28 N_87 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M29 N_82 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M30 N_14 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M31 VDD N_14 N_12 VDD mp15  l=0.13u w=0.49u m=1
M32 N_17 N_12 N_75 VDD mp15  l=0.13u w=0.58u m=1
M33 VDD N_21 N_88 VDD mp15  l=0.13u w=0.26u m=1
M34 N_17 N_14 N_88 VDD mp15  l=0.13u w=0.26u m=1
M35 N_23 N_19 VDD VDD mp15  l=0.13u w=0.4u m=1
M36 N_25 RN VDD VDD mp15  l=0.13u w=0.4u m=1
M37 N_21 N_14 N_19 VDD mp15  l=0.13u w=0.4u m=1
M38 N_21 N_17 N_79 VDD mp15  l=0.13u w=0.4u m=1
M39 N_79 N_25 VDD VDD mp15  l=0.13u w=0.4u m=1
M40 VDD N_25 N_79 VDD mp15  l=0.13u w=0.4u m=1
M41 N_89 N_12 N_19 VDD mp15  l=0.13u w=0.26u m=1
M42 N_89 N_33 N_79 VDD mp15  l=0.13u w=0.26u m=1
M43 QN N_19 VDD VDD mp15  l=0.13u w=0.4u m=1
M44 Q N_23 VDD VDD mp15  l=0.13u w=0.4u m=1
M45 N_36 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M46 N_35 N_33 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M47 N_33 RETN N_90 VDDG mp15  l=0.13u w=0.26u m=1
M48 N_33 N_36 N_23 VDDG mp15  l=0.13u w=0.26u m=1
M49 VDDG N_35 N_90 VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrcrb0
* SPICE INPUT		Tue Sep 18 13:28:52 2018	sdrcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrcrb1
.subckt sdrcrb1 VDD VDDG GND Q QN SI CK D SE RN RETN
M1 N_7 N_10 N_40 GND mn15  l=0.13u w=0.26u m=1
M2 GND N_9 N_40 GND mn15  l=0.13u w=0.26u m=1
M3 N_9 N_7 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_10 RETN GND GND mn15  l=0.13u w=0.26u m=1
M5 N_7 RETN N_11 GND mn15  l=0.13u w=0.26u m=1
M6 Q N_11 GND GND mn15  l=0.13u w=0.46u m=1
M7 QN N_18 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_52 N_7 GND GND mn15  l=0.13u w=0.26u m=1
M9 N_18 N_28 N_52 GND mn15  l=0.13u w=0.26u m=1
M10 GND N_18 N_11 GND mn15  l=0.13u w=0.39u m=1
M11 N_21 RN GND GND mn15  l=0.13u w=0.3u m=1
M12 GND N_38 N_57 GND mn15  l=0.13u w=0.26u m=1
M13 N_24 N_26 N_57 GND mn15  l=0.13u w=0.26u m=1
M14 N_25 N_28 N_24 GND mn15  l=0.13u w=0.44u m=1
M15 GND N_28 N_26 GND mn15  l=0.13u w=0.19u m=1
M16 N_28 CK GND GND mn15  l=0.13u w=0.21u m=1
M17 N_65 SI GND GND mn15  l=0.13u w=0.26u m=1
M18 N_25 SE N_65 GND mn15  l=0.13u w=0.26u m=1
M19 N_68 D N_25 GND mn15  l=0.13u w=0.44u m=1
M20 N_68 N_34 GND GND mn15  l=0.13u w=0.44u m=1
M21 GND SE N_34 GND mn15  l=0.13u w=0.26u m=1
M22 N_18 N_26 N_38 GND mn15  l=0.13u w=0.39u m=1
M23 GND N_21 N_18 GND mn15  l=0.13u w=0.4u m=1
M24 N_38 N_24 GND GND mn15  l=0.13u w=0.4u m=1
M25 Q N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 QN N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_87 N_7 N_83 VDD mp15  l=0.13u w=0.26u m=1
M28 N_87 N_26 N_18 VDD mp15  l=0.13u w=0.26u m=1
M29 N_83 N_21 VDD VDD mp15  l=0.13u w=0.58u m=1
M30 VDD N_21 N_83 VDD mp15  l=0.13u w=0.58u m=1
M31 N_83 N_24 N_38 VDD mp15  l=0.13u w=0.58u m=1
M32 N_38 N_28 N_18 VDD mp15  l=0.13u w=0.58u m=1
M33 N_11 N_18 VDD VDD mp15  l=0.13u w=0.58u m=1
M34 N_21 RN VDD VDD mp15  l=0.13u w=0.5u m=1
M35 N_24 N_28 N_88 VDD mp15  l=0.13u w=0.26u m=1
M36 VDD N_38 N_88 VDD mp15  l=0.13u w=0.26u m=1
M37 N_24 N_26 N_78 VDD mp15  l=0.13u w=0.58u m=1
M38 VDD N_28 N_26 VDD mp15  l=0.13u w=0.49u m=1
M39 N_28 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M40 N_75 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M41 N_89 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M42 N_89 D N_78 VDD mp15  l=0.13u w=0.58u m=1
M43 N_78 N_34 N_75 VDD mp15  l=0.13u w=0.26u m=1
M44 VDD SE N_34 VDD mp15  l=0.13u w=0.39u m=1
M45 N_7 RETN N_90 VDDG mp15  l=0.13u w=0.26u m=1
M46 N_7 N_10 N_11 VDDG mp15  l=0.13u w=0.26u m=1
M47 VDDG N_9 N_90 VDDG mp15  l=0.13u w=0.26u m=1
M48 N_9 N_7 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M49 N_10 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrcrb1
* SPICE INPUT		Tue Sep 18 13:28:59 2018	sdrcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrcrb2
.subckt sdrcrb2 VDD VDDG GND QN Q RN RETN CK SI SE D
M1 GND SE N_5 GND mn15  l=0.13u w=0.26u m=1
M2 N_48 N_5 GND GND mn15  l=0.13u w=0.44u m=1
M3 N_48 D N_10 GND mn15  l=0.13u w=0.44u m=1
M4 N_10 SE N_45 GND mn15  l=0.13u w=0.26u m=1
M5 N_45 SI GND GND mn15  l=0.13u w=0.26u m=1
M6 N_14 CK GND GND mn15  l=0.13u w=0.27u m=1
M7 GND N_14 N_12 GND mn15  l=0.13u w=0.21u m=1
M8 N_56 N_12 N_17 GND mn15  l=0.13u w=0.26u m=1
M9 GND N_15 N_56 GND mn15  l=0.13u w=0.26u m=1
M10 GND N_17 N_15 GND mn15  l=0.13u w=0.46u m=1
M11 N_10 N_14 N_17 GND mn15  l=0.13u w=0.44u m=1
M12 N_16 N_12 N_15 GND mn15  l=0.13u w=0.46u m=1
M13 GND RN N_24 GND mn15  l=0.13u w=0.2u m=1
M14 N_24 RN GND GND mn15  l=0.13u w=0.19u m=1
M15 GND N_16 QN GND mn15  l=0.13u w=0.586u m=1
M16 GND N_16 QN GND mn15  l=0.13u w=0.334u m=1
M17 GND N_24 N_16 GND mn15  l=0.13u w=0.46u m=1
M18 N_68 N_14 N_16 GND mn15  l=0.13u w=0.26u m=1
M19 GND N_29 N_68 GND mn15  l=0.13u w=0.26u m=1
M20 GND N_16 N_28 GND mn15  l=0.13u w=0.46u m=1
M21 N_29 RETN N_28 GND mn15  l=0.13u w=0.26u m=1
M22 GND N_28 Q GND mn15  l=0.13u w=0.46u m=1
M23 GND N_28 Q GND mn15  l=0.13u w=0.46u m=1
M24 N_38 RETN GND GND mn15  l=0.13u w=0.26u m=1
M25 N_37 N_29 GND GND mn15  l=0.13u w=0.26u m=1
M26 N_29 N_38 N_76 GND mn15  l=0.13u w=0.26u m=1
M27 GND N_37 N_76 GND mn15  l=0.13u w=0.26u m=1
M28 VDD SE N_5 VDD mp15  l=0.13u w=0.39u m=1
M29 N_80 N_5 N_86 VDD mp15  l=0.13u w=0.26u m=1
M30 N_90 D N_80 VDD mp15  l=0.13u w=0.69u m=1
M31 N_90 SE VDD VDD mp15  l=0.13u w=0.69u m=1
M32 VDD SI N_86 VDD mp15  l=0.13u w=0.26u m=1
M33 N_14 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M34 VDD N_14 N_12 VDD mp15  l=0.13u w=0.54u m=1
M35 N_17 N_12 N_80 VDD mp15  l=0.13u w=0.69u m=1
M36 VDD N_15 N_91 VDD mp15  l=0.13u w=0.26u m=1
M37 N_17 N_14 N_91 VDD mp15  l=0.13u w=0.26u m=1
M38 N_24 RN VDD VDD mp15  l=0.13u w=0.29u m=1
M39 N_24 RN VDD VDD mp15  l=0.13u w=0.29u m=1
M40 N_82 N_17 N_15 VDD mp15  l=0.13u w=0.69u m=1
M41 N_15 N_14 N_16 VDD mp15  l=0.13u w=0.69u m=1
M42 VDD N_24 N_82 VDD mp15  l=0.13u w=0.69u m=1
M43 N_82 N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M44 N_16 N_12 N_92 VDD mp15  l=0.13u w=0.26u m=1
M45 N_82 N_29 N_92 VDD mp15  l=0.13u w=0.26u m=1
M46 QN N_16 VDD VDD mp15  l=0.13u w=1.12u m=1
M47 QN N_16 VDD VDD mp15  l=0.13u w=0.26u m=1
M48 VDD N_28 Q VDD mp15  l=0.13u w=0.69u m=1
M49 VDD N_28 Q VDD mp15  l=0.13u w=0.69u m=1
M50 N_28 N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M51 N_38 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M52 N_37 N_29 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M53 N_29 N_38 N_28 VDDG mp15  l=0.13u w=0.26u m=1
M54 VDDG N_37 N_93 VDDG mp15  l=0.13u w=0.26u m=1
M55 N_29 RETN N_93 VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrcrb2
* SPICE INPUT		Tue Sep 18 13:29:05 2018	sdrcrbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrcrbm
.subckt sdrcrbm VDD VDDG GND Q QN RETN RN SI CK D SE
M1 GND SE N_5 GND mn15  l=0.13u w=0.26u m=1
M2 N_46 N_5 GND GND mn15  l=0.13u w=0.4u m=1
M3 N_46 D N_10 GND mn15  l=0.13u w=0.4u m=1
M4 N_10 SE N_43 GND mn15  l=0.13u w=0.26u m=1
M5 N_43 SI GND GND mn15  l=0.13u w=0.26u m=1
M6 N_14 CK GND GND mn15  l=0.13u w=0.21u m=1
M7 GND N_14 N_12 GND mn15  l=0.13u w=0.19u m=1
M8 N_10 N_14 N_17 GND mn15  l=0.13u w=0.4u m=1
M9 N_17 N_12 N_50 GND mn15  l=0.13u w=0.26u m=1
M10 GND N_21 N_50 GND mn15  l=0.13u w=0.26u m=1
M11 N_21 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M12 GND N_25 N_19 GND mn15  l=0.13u w=0.26u m=1
M13 N_19 N_12 N_21 GND mn15  l=0.13u w=0.26u m=1
M14 GND N_19 N_23 GND mn15  l=0.13u w=0.26u m=1
M15 N_25 RN GND GND mn15  l=0.13u w=0.26u m=1
M16 N_19 N_14 N_62 GND mn15  l=0.13u w=0.26u m=1
M17 N_62 N_33 GND GND mn15  l=0.13u w=0.26u m=1
M18 QN N_19 GND GND mn15  l=0.13u w=0.36u m=1
M19 Q N_23 GND GND mn15  l=0.13u w=0.36u m=1
M20 N_33 RETN N_23 GND mn15  l=0.13u w=0.26u m=1
M21 N_36 RETN GND GND mn15  l=0.13u w=0.26u m=1
M22 N_35 N_33 GND GND mn15  l=0.13u w=0.26u m=1
M23 N_33 N_36 N_72 GND mn15  l=0.13u w=0.26u m=1
M24 GND N_35 N_72 GND mn15  l=0.13u w=0.26u m=1
M25 VDD SE N_5 VDD mp15  l=0.13u w=0.39u m=1
M26 N_75 N_5 N_82 VDD mp15  l=0.13u w=0.26u m=1
M27 N_87 D N_75 VDD mp15  l=0.13u w=0.58u m=1
M28 N_87 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M29 N_82 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M30 N_14 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M31 VDD N_14 N_12 VDD mp15  l=0.13u w=0.49u m=1
M32 N_17 N_12 N_75 VDD mp15  l=0.13u w=0.58u m=1
M33 VDD N_21 N_88 VDD mp15  l=0.13u w=0.26u m=1
M34 N_17 N_14 N_88 VDD mp15  l=0.13u w=0.26u m=1
M35 N_23 N_19 VDD VDD mp15  l=0.13u w=0.4u m=1
M36 N_25 RN VDD VDD mp15  l=0.13u w=0.4u m=1
M37 N_21 N_14 N_19 VDD mp15  l=0.13u w=0.4u m=1
M38 N_21 N_17 N_79 VDD mp15  l=0.13u w=0.4u m=1
M39 N_79 N_25 VDD VDD mp15  l=0.13u w=0.4u m=1
M40 VDD N_25 N_79 VDD mp15  l=0.13u w=0.4u m=1
M41 N_89 N_12 N_19 VDD mp15  l=0.13u w=0.26u m=1
M42 N_89 N_33 N_79 VDD mp15  l=0.13u w=0.26u m=1
M43 QN N_19 VDD VDD mp15  l=0.13u w=0.55u m=1
M44 Q N_23 VDD VDD mp15  l=0.13u w=0.55u m=1
M45 N_36 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M46 N_35 N_33 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M47 N_33 RETN N_90 VDDG mp15  l=0.13u w=0.26u m=1
M48 N_33 N_36 N_23 VDDG mp15  l=0.13u w=0.26u m=1
M49 VDDG N_35 N_90 VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrcrbm
* SPICE INPUT		Tue Sep 18 13:29:12 2018	sdrnrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrnrb0
.subckt sdrnrb0 VDD VDDG GND Q QN RETN SI SE CK D
M1 N_6 SE GND GND mn15  l=0.13u w=0.26u m=1
M2 N_9 CK GND GND mn15  l=0.13u w=0.21u m=1
M3 GND N_9 N_7 GND mn15  l=0.13u w=0.19u m=1
M4 N_46 D N_12 GND mn15  l=0.13u w=0.36u m=1
M5 N_46 N_6 GND GND mn15  l=0.13u w=0.36u m=1
M6 N_48 SI GND GND mn15  l=0.13u w=0.26u m=1
M7 N_48 SE N_12 GND mn15  l=0.13u w=0.26u m=1
M8 N_17 N_9 N_12 GND mn15  l=0.13u w=0.36u m=1
M9 N_50 N_11 GND GND mn15  l=0.13u w=0.26u m=1
M10 N_11 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_50 N_7 N_17 GND mn15  l=0.13u w=0.26u m=1
M12 N_20 N_23 GND GND mn15  l=0.13u w=0.26u m=1
M13 Q N_23 GND GND mn15  l=0.13u w=0.26u m=1
M14 GND N_11 N_54 GND mn15  l=0.13u w=0.39u m=1
M15 N_23 N_7 N_54 GND mn15  l=0.13u w=0.39u m=1
M16 GND N_20 QN GND mn15  l=0.13u w=0.26u m=1
M17 N_23 N_9 N_59 GND mn15  l=0.13u w=0.26u m=1
M18 GND N_32 N_59 GND mn15  l=0.13u w=0.26u m=1
M19 N_31 RETN GND GND mn15  l=0.13u w=0.26u m=1
M20 GND N_32 N_34 GND mn15  l=0.13u w=0.26u m=1
M21 N_68 N_34 GND GND mn15  l=0.13u w=0.26u m=1
M22 N_20 RETN N_32 GND mn15  l=0.13u w=0.26u m=1
M23 N_68 N_31 N_32 GND mn15  l=0.13u w=0.26u m=1
M24 VDD SE N_6 VDD mp15  l=0.13u w=0.4u m=1
M25 N_84 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M26 N_72 D N_84 VDD mp15  l=0.13u w=0.58u m=1
M27 N_72 N_6 N_83 VDD mp15  l=0.13u w=0.26u m=1
M28 N_83 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M29 N_9 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M30 N_7 N_9 VDD VDD mp15  l=0.13u w=0.49u m=1
M31 N_85 N_9 N_17 VDD mp15  l=0.13u w=0.26u m=1
M32 N_85 N_11 VDD VDD mp15  l=0.13u w=0.26u m=1
M33 N_11 N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M34 N_72 N_7 N_17 VDD mp15  l=0.13u w=0.58u m=1
M35 Q N_23 VDD VDD mp15  l=0.13u w=0.4u m=1
M36 N_20 N_23 VDD VDD mp15  l=0.13u w=0.4u m=1
M37 QN N_20 VDD VDD mp15  l=0.13u w=0.4u m=1
M38 N_23 N_9 N_86 VDD mp15  l=0.13u w=0.58u m=1
M39 VDD N_11 N_86 VDD mp15  l=0.13u w=0.58u m=1
M40 N_23 N_7 N_87 VDDG mp15  l=0.13u w=0.26u m=1
M41 VDD N_32 N_87 VDDG mp15  l=0.13u w=0.26u m=1
M42 VDDG N_32 N_34 VDDG mp15  l=0.13u w=0.26u m=1
M43 N_88 N_34 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M44 N_88 RETN N_32 VDDG mp15  l=0.13u w=0.26u m=1
M45 N_20 N_31 N_32 VDDG mp15  l=0.13u w=0.26u m=1
M46 N_31 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrnrb0
* SPICE INPUT		Tue Sep 18 13:29:19 2018	sdrnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrnrb1
.subckt sdrnrb1 VDD VDDG GND Q QN RETN SI SE CK D
M1 N_6 SE GND GND mn15  l=0.13u w=0.26u m=1
M2 N_9 CK GND GND mn15  l=0.13u w=0.21u m=1
M3 GND N_9 N_7 GND mn15  l=0.13u w=0.19u m=1
M4 N_47 D N_12 GND mn15  l=0.13u w=0.4u m=1
M5 GND N_6 N_47 GND mn15  l=0.13u w=0.4u m=1
M6 N_50 SI GND GND mn15  l=0.13u w=0.26u m=1
M7 N_50 SE N_12 GND mn15  l=0.13u w=0.26u m=1
M8 N_17 N_9 N_12 GND mn15  l=0.13u w=0.4u m=1
M9 N_52 N_11 GND GND mn15  l=0.13u w=0.26u m=1
M10 N_11 N_17 GND GND mn15  l=0.13u w=0.39u m=1
M11 N_52 N_7 N_17 GND mn15  l=0.13u w=0.26u m=1
M12 Q N_25 GND GND mn15  l=0.13u w=0.235u m=1
M13 GND N_25 Q GND mn15  l=0.13u w=0.225u m=1
M14 N_20 N_25 GND GND mn15  l=0.13u w=0.2u m=1
M15 GND N_25 N_20 GND mn15  l=0.13u w=0.2u m=1
M16 GND N_11 N_58 GND mn15  l=0.13u w=0.46u m=1
M17 N_25 N_7 N_58 GND mn15  l=0.13u w=0.46u m=1
M18 GND N_20 QN GND mn15  l=0.13u w=0.46u m=1
M19 N_25 N_9 N_63 GND mn15  l=0.13u w=0.26u m=1
M20 GND N_34 N_63 GND mn15  l=0.13u w=0.26u m=1
M21 N_33 RETN GND GND mn15  l=0.13u w=0.26u m=1
M22 GND N_34 N_36 GND mn15  l=0.13u w=0.26u m=1
M23 N_72 N_36 GND GND mn15  l=0.13u w=0.26u m=1
M24 N_20 RETN N_34 GND mn15  l=0.13u w=0.26u m=1
M25 N_72 N_33 N_34 GND mn15  l=0.13u w=0.26u m=1
M26 VDD SE N_6 VDD mp15  l=0.13u w=0.4u m=1
M27 N_88 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M28 N_76 D N_88 VDD mp15  l=0.13u w=0.58u m=1
M29 N_76 N_6 N_87 VDD mp15  l=0.13u w=0.26u m=1
M30 N_87 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M31 N_9 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M32 N_7 N_9 VDD VDD mp15  l=0.13u w=0.49u m=1
M33 N_89 N_9 N_17 VDD mp15  l=0.13u w=0.26u m=1
M34 N_89 N_11 VDD VDD mp15  l=0.13u w=0.26u m=1
M35 N_11 N_17 VDD VDD mp15  l=0.13u w=0.58u m=1
M36 N_76 N_7 N_17 VDD mp15  l=0.13u w=0.58u m=1
M37 Q N_25 VDD VDD mp15  l=0.13u w=0.69u m=1
M38 N_20 N_25 VDD VDD mp15  l=0.13u w=0.6u m=1
M39 VDD N_20 QN VDD mp15  l=0.13u w=0.345u m=1
M40 VDD N_20 QN VDD mp15  l=0.13u w=0.345u m=1
M41 N_25 N_9 N_90 VDD mp15  l=0.13u w=0.69u m=1
M42 VDD N_11 N_90 VDD mp15  l=0.13u w=0.69u m=1
M43 N_25 N_7 N_91 VDDG mp15  l=0.13u w=0.26u m=1
M44 VDD N_34 N_91 VDDG mp15  l=0.13u w=0.26u m=1
M45 VDDG N_34 N_36 VDDG mp15  l=0.13u w=0.26u m=1
M46 N_92 N_36 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M47 N_92 RETN N_34 VDDG mp15  l=0.13u w=0.26u m=1
M48 N_20 N_33 N_34 VDDG mp15  l=0.13u w=0.26u m=1
M49 N_33 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrnrb1
* SPICE INPUT		Tue Sep 18 13:29:25 2018	sdrnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrnrb2
.subckt sdrnrb2 VDD VDDG GND Q QN SE SI D CK RETN
M1 N_7 N_10 N_40 GND mn15  l=0.13u w=0.26u m=1
M2 GND N_9 N_40 GND mn15  l=0.13u w=0.26u m=1
M3 N_9 N_7 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_10 RETN GND GND mn15  l=0.13u w=0.26u m=1
M5 Q N_18 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_18 Q GND mn15  l=0.13u w=0.46u m=1
M7 N_7 RETN N_14 GND mn15  l=0.13u w=0.26u m=1
M8 GND N_7 N_51 GND mn15  l=0.13u w=0.26u m=1
M9 N_18 N_26 N_51 GND mn15  l=0.13u w=0.26u m=1
M10 GND N_18 N_14 GND mn15  l=0.13u w=0.46u m=1
M11 N_57 N_29 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_57 N_27 N_18 GND mn15  l=0.13u w=0.46u m=1
M13 GND SE N_23 GND mn15  l=0.13u w=0.26u m=1
M14 N_27 N_26 GND GND mn15  l=0.13u w=0.21u m=1
M15 N_26 CK GND GND mn15  l=0.13u w=0.28u m=1
M16 N_71 N_27 N_35 GND mn15  l=0.13u w=0.26u m=1
M17 N_29 N_35 GND GND mn15  l=0.13u w=0.39u m=1
M18 N_71 N_29 GND GND mn15  l=0.13u w=0.26u m=1
M19 N_35 N_26 N_30 GND mn15  l=0.13u w=0.44u m=1
M20 N_30 SE N_68 GND mn15  l=0.13u w=0.26u m=1
M21 N_68 SI GND GND mn15  l=0.13u w=0.26u m=1
M22 N_67 N_23 GND GND mn15  l=0.13u w=0.44u m=1
M23 N_67 D N_30 GND mn15  l=0.13u w=0.44u m=1
M24 GND N_14 QN GND mn15  l=0.13u w=0.46u m=1
M25 GND N_14 QN GND mn15  l=0.13u w=0.46u m=1
M26 N_14 N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_84 N_29 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 N_84 N_26 N_18 VDD mp15  l=0.13u w=0.69u m=1
M29 Q N_18 VDD VDD mp15  l=0.13u w=0.47u m=1
M30 Q N_18 VDD VDD mp15  l=0.13u w=0.47u m=1
M31 VDD N_18 Q VDD mp15  l=0.13u w=0.44u m=1
M32 VDD N_14 QN VDD mp15  l=0.13u w=0.78u m=1
M33 QN N_14 VDD VDD mp15  l=0.13u w=0.6u m=1
M34 N_77 N_27 N_35 VDD mp15  l=0.13u w=0.58u m=1
M35 N_29 N_35 VDD VDD mp15  l=0.13u w=0.58u m=1
M36 N_85 N_29 VDD VDD mp15  l=0.13u w=0.26u m=1
M37 N_85 N_26 N_35 VDD mp15  l=0.13u w=0.26u m=1
M38 N_27 N_26 VDD VDD mp15  l=0.13u w=0.54u m=1
M39 N_87 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M40 N_26 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M41 N_86 SE VDD VDD mp15  l=0.13u w=0.69u m=1
M42 VDD SE N_23 VDD mp15  l=0.13u w=0.4u m=1
M43 N_87 N_23 N_77 VDD mp15  l=0.13u w=0.26u m=1
M44 N_86 D N_77 VDD mp15  l=0.13u w=0.69u m=1
M45 N_7 RETN N_88 VDDG mp15  l=0.13u w=0.26u m=1
M46 N_88 N_9 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M47 N_9 N_7 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M48 N_10 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M49 VDD N_7 N_89 VDDG mp15  l=0.13u w=0.26u m=1
M50 N_18 N_27 N_89 VDDG mp15  l=0.13u w=0.26u m=1
M51 N_14 N_10 N_7 VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrnrb2
* SPICE INPUT		Tue Sep 18 13:29:31 2018	sdrnrbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrnrbm
.subckt sdrnrbm VDD VDDG GND Q QN RETN SI SE CK D
M1 N_6 SE GND GND mn15  l=0.13u w=0.26u m=1
M2 N_9 CK GND GND mn15  l=0.13u w=0.21u m=1
M3 GND N_9 N_7 GND mn15  l=0.13u w=0.19u m=1
M4 N_47 D N_12 GND mn15  l=0.13u w=0.36u m=1
M5 N_47 N_6 GND GND mn15  l=0.13u w=0.36u m=1
M6 N_49 SI GND GND mn15  l=0.13u w=0.26u m=1
M7 N_49 SE N_12 GND mn15  l=0.13u w=0.26u m=1
M8 N_17 N_9 N_12 GND mn15  l=0.13u w=0.36u m=1
M9 N_51 N_11 GND GND mn15  l=0.13u w=0.26u m=1
M10 N_11 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_51 N_7 N_17 GND mn15  l=0.13u w=0.26u m=1
M12 N_20 N_24 GND GND mn15  l=0.13u w=0.26u m=1
M13 Q N_24 GND GND mn15  l=0.13u w=0.18u m=1
M14 Q N_24 GND GND mn15  l=0.13u w=0.18u m=1
M15 GND N_11 N_56 GND mn15  l=0.13u w=0.39u m=1
M16 N_24 N_7 N_56 GND mn15  l=0.13u w=0.39u m=1
M17 GND N_20 QN GND mn15  l=0.13u w=0.36u m=1
M18 N_24 N_9 N_61 GND mn15  l=0.13u w=0.26u m=1
M19 GND N_33 N_61 GND mn15  l=0.13u w=0.26u m=1
M20 N_32 RETN GND GND mn15  l=0.13u w=0.26u m=1
M21 GND N_33 N_35 GND mn15  l=0.13u w=0.26u m=1
M22 N_70 N_35 GND GND mn15  l=0.13u w=0.26u m=1
M23 N_20 RETN N_33 GND mn15  l=0.13u w=0.26u m=1
M24 N_70 N_32 N_33 GND mn15  l=0.13u w=0.26u m=1
M25 VDD SE N_6 VDD mp15  l=0.13u w=0.4u m=1
M26 N_86 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M27 N_74 D N_86 VDD mp15  l=0.13u w=0.58u m=1
M28 N_74 N_6 N_85 VDD mp15  l=0.13u w=0.26u m=1
M29 N_85 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M30 N_9 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M31 N_7 N_9 VDD VDD mp15  l=0.13u w=0.49u m=1
M32 N_87 N_9 N_17 VDD mp15  l=0.13u w=0.26u m=1
M33 N_87 N_11 VDD VDD mp15  l=0.13u w=0.26u m=1
M34 N_11 N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M35 N_74 N_7 N_17 VDD mp15  l=0.13u w=0.58u m=1
M36 Q N_24 VDD VDD mp15  l=0.13u w=0.55u m=1
M37 N_20 N_24 VDD VDD mp15  l=0.13u w=0.4u m=1
M38 QN N_20 VDD VDD mp15  l=0.13u w=0.55u m=1
M39 N_24 N_9 N_88 VDD mp15  l=0.13u w=0.58u m=1
M40 VDD N_11 N_88 VDD mp15  l=0.13u w=0.58u m=1
M41 N_24 N_7 N_89 VDDG mp15  l=0.13u w=0.26u m=1
M42 VDD N_33 N_89 VDDG mp15  l=0.13u w=0.26u m=1
M43 VDDG N_33 N_35 VDDG mp15  l=0.13u w=0.26u m=1
M44 N_90 N_35 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M45 N_90 RETN N_33 VDDG mp15  l=0.13u w=0.26u m=1
M46 N_20 N_32 N_33 VDDG mp15  l=0.13u w=0.26u m=1
M47 N_32 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrnrbm
* SPICE INPUT		Tue Sep 18 13:29:37 2018	sdrprb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrprb0
.subckt sdrprb0 VDD VDDG GND QN Q RETN SN SI SE CK D
M1 N_6 SE GND GND mn15  l=0.13u w=0.26u m=1
M2 N_9 CK GND GND mn15  l=0.13u w=0.21u m=1
M3 GND N_9 N_7 GND mn15  l=0.13u w=0.19u m=1
M4 N_45 D N_12 GND mn15  l=0.13u w=0.36u m=1
M5 GND N_6 N_45 GND mn15  l=0.13u w=0.36u m=1
M6 N_48 SI GND GND mn15  l=0.13u w=0.26u m=1
M7 N_48 SE N_12 GND mn15  l=0.13u w=0.26u m=1
M8 N_17 N_9 N_12 GND mn15  l=0.13u w=0.36u m=1
M9 N_43 N_21 GND GND mn15  l=0.13u w=0.26u m=1
M10 N_17 N_7 N_43 GND mn15  l=0.13u w=0.26u m=1
M11 N_19 N_32 GND GND mn15  l=0.13u w=0.26u m=1
M12 QN N_32 GND GND mn15  l=0.13u w=0.26u m=1
M13 N_22 N_17 N_21 GND mn15  l=0.13u w=0.3u m=1
M14 GND N_23 N_25 GND mn15  l=0.13u w=0.26u m=1
M15 N_59 N_25 GND GND mn15  l=0.13u w=0.26u m=1
M16 N_59 N_36 N_23 GND mn15  l=0.13u w=0.26u m=1
M17 N_19 RETN N_23 GND mn15  l=0.13u w=0.26u m=1
M18 GND N_19 Q GND mn15  l=0.13u w=0.26u m=1
M19 N_21 N_7 N_32 GND mn15  l=0.13u w=0.26u m=1
M20 N_66 N_9 N_32 GND mn15  l=0.13u w=0.26u m=1
M21 GND SN N_22 GND mn15  l=0.13u w=0.6u m=1
M22 N_66 N_23 N_22 GND mn15  l=0.13u w=0.26u m=1
M23 N_36 RETN GND GND mn15  l=0.13u w=0.26u m=1
M24 VDD SE N_6 VDD mp15  l=0.13u w=0.39u m=1
M25 N_84 SE VDD VDD mp15  l=0.13u w=0.55u m=1
M26 N_84 D N_73 VDD mp15  l=0.13u w=0.55u m=1
M27 N_73 N_6 N_83 VDD mp15  l=0.13u w=0.26u m=1
M28 N_83 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M29 N_9 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M30 N_7 N_9 VDD VDD mp15  l=0.13u w=0.49u m=1
M31 QN N_32 VDD VDD mp15  l=0.13u w=0.4u m=1
M32 N_19 N_32 VDD VDD mp15  l=0.13u w=0.4u m=1
M33 N_85 N_9 N_17 VDD mp15  l=0.13u w=0.26u m=1
M34 VDD N_21 N_85 VDD mp15  l=0.13u w=0.26u m=1
M35 VDD N_17 N_21 VDD mp15  l=0.13u w=0.4u m=1
M36 N_32 N_9 N_21 VDD mp15  l=0.13u w=0.4u m=1
M37 N_73 N_7 N_17 VDD mp15  l=0.13u w=0.55u m=1
M38 VDD N_19 Q VDD mp15  l=0.13u w=0.4u m=1
M39 N_86 N_7 N_32 VDD mp15  l=0.13u w=0.26u m=1
M40 N_32 SN VDD VDD mp15  l=0.13u w=0.4u m=1
M41 N_86 N_23 VDD VDD mp15  l=0.13u w=0.26u m=1
M42 N_36 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M43 VDDG N_23 N_25 VDDG mp15  l=0.13u w=0.26u m=1
M44 N_87 N_25 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M45 N_19 N_36 N_23 VDDG mp15  l=0.13u w=0.26u m=1
M46 N_87 RETN N_23 VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrprb0
* SPICE INPUT		Tue Sep 18 13:29:44 2018	sdrprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrprb1
.subckt sdrprb1 VDDG VDD GND QN Q RETN SN SI SE CK D
M1 N_6 SE GND GND mn15  l=0.13u w=0.26u m=1
M2 N_9 CK GND GND mn15  l=0.13u w=0.21u m=1
M3 GND N_9 N_7 GND mn15  l=0.13u w=0.19u m=1
M4 N_11 N_39 N_10 GND mn15  l=0.13u w=0.4u m=1
M5 GND N_22 QN GND mn15  l=0.13u w=0.23u m=1
M6 QN N_22 GND GND mn15  l=0.13u w=0.23u m=1
M7 GND N_22 N_13 GND mn15  l=0.13u w=0.2u m=1
M8 N_13 N_22 GND GND mn15  l=0.13u w=0.19u m=1
M9 GND N_13 Q GND mn15  l=0.13u w=0.46u m=1
M10 N_22 N_7 N_10 GND mn15  l=0.13u w=0.39u m=1
M11 N_58 N_9 N_22 GND mn15  l=0.13u w=0.26u m=1
M12 N_11 SN GND GND mn15  l=0.13u w=0.4u m=1
M13 N_11 SN GND GND mn15  l=0.13u w=0.4u m=1
M14 N_11 N_27 N_58 GND mn15  l=0.13u w=0.26u m=1
M15 N_26 RETN GND GND mn15  l=0.13u w=0.26u m=1
M16 GND N_27 N_29 GND mn15  l=0.13u w=0.26u m=1
M17 N_66 N_29 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_13 RETN N_27 GND mn15  l=0.13u w=0.26u m=1
M19 N_66 N_26 N_27 GND mn15  l=0.13u w=0.26u m=1
M20 N_70 D N_34 GND mn15  l=0.13u w=0.4u m=1
M21 GND N_6 N_70 GND mn15  l=0.13u w=0.4u m=1
M22 N_73 SI GND GND mn15  l=0.13u w=0.26u m=1
M23 N_73 SE N_34 GND mn15  l=0.13u w=0.26u m=1
M24 N_39 N_9 N_34 GND mn15  l=0.13u w=0.4u m=1
M25 N_68 N_10 GND GND mn15  l=0.13u w=0.26u m=1
M26 N_39 N_7 N_68 GND mn15  l=0.13u w=0.26u m=1
M27 VDD SE N_6 VDD mp15  l=0.13u w=0.4u m=1
M28 N_90 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M29 N_90 D N_79 VDD mp15  l=0.13u w=0.58u m=1
M30 N_79 N_6 N_89 VDD mp15  l=0.13u w=0.26u m=1
M31 N_89 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M32 N_9 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M33 N_7 N_9 VDD VDD mp15  l=0.13u w=0.49u m=1
M34 N_91 N_9 N_39 VDD mp15  l=0.13u w=0.26u m=1
M35 VDD N_10 N_91 VDD mp15  l=0.13u w=0.26u m=1
M36 VDD N_39 N_10 VDD mp15  l=0.13u w=0.58u m=1
M37 N_22 N_9 N_10 VDD mp15  l=0.13u w=0.58u m=1
M38 N_79 N_7 N_39 VDD mp15  l=0.13u w=0.58u m=1
M39 VDD N_13 Q VDD mp15  l=0.13u w=0.43u m=1
M40 VDD N_13 Q VDD mp15  l=0.13u w=0.26u m=1
M41 N_92 N_7 N_22 VDD mp15  l=0.13u w=0.26u m=1
M42 N_22 SN VDD VDD mp15  l=0.13u w=0.26u m=1
M43 N_92 N_27 VDD VDD mp15  l=0.13u w=0.26u m=1
M44 QN N_22 VDD VDD mp15  l=0.13u w=0.69u m=1
M45 N_13 N_22 VDD VDD mp15  l=0.13u w=0.58u m=1
M46 N_26 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M47 VDDG N_27 N_29 VDDG mp15  l=0.13u w=0.26u m=1
M48 N_93 N_29 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M49 N_93 RETN N_27 VDDG mp15  l=0.13u w=0.26u m=1
M50 N_13 N_26 N_27 VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrprb1
* SPICE INPUT		Tue Sep 18 13:29:50 2018	sdrprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrprb2
.subckt sdrprb2 VDD VDDG GND Q QN RETN SN SI SE D CK
M1 GND SE N_5 GND mn15  l=0.13u w=0.26u m=1
M2 N_9 N_8 GND GND mn15  l=0.13u w=0.21u m=1
M3 N_8 CK GND GND mn15  l=0.13u w=0.27u m=1
M4 GND N_31 Q GND mn15  l=0.13u w=0.46u m=1
M5 GND N_31 Q GND mn15  l=0.13u w=0.46u m=1
M6 N_17 D N_15 GND mn15  l=0.13u w=0.44u m=1
M7 N_17 N_5 GND GND mn15  l=0.13u w=0.44u m=1
M8 N_18 SI GND GND mn15  l=0.13u w=0.26u m=1
M9 N_15 SE N_18 GND mn15  l=0.13u w=0.26u m=1
M10 N_15 N_8 N_19 GND mn15  l=0.13u w=0.44u m=1
M11 GND N_25 N_13 GND mn15  l=0.13u w=0.26u m=1
M12 N_19 N_9 N_13 GND mn15  l=0.13u w=0.26u m=1
M13 N_25 N_19 N_22 GND mn15  l=0.13u w=0.46u m=1
M14 N_25 N_9 N_24 GND mn15  l=0.13u w=0.46u m=1
M15 N_26 N_8 N_24 GND mn15  l=0.13u w=0.26u m=1
M16 N_22 SN GND GND mn15  l=0.13u w=0.46u m=1
M17 N_22 SN GND GND mn15  l=0.13u w=0.46u m=1
M18 N_22 N_39 N_26 GND mn15  l=0.13u w=0.26u m=1
M19 QN N_24 GND GND mn15  l=0.13u w=0.46u m=1
M20 GND N_24 QN GND mn15  l=0.13u w=0.46u m=1
M21 GND N_24 N_31 GND mn15  l=0.13u w=0.46u m=1
M22 N_35 RETN GND GND mn15  l=0.13u w=0.26u m=1
M23 N_34 N_39 GND GND mn15  l=0.13u w=0.26u m=1
M24 N_39 RETN N_31 GND mn15  l=0.13u w=0.26u m=1
M25 N_39 N_35 N_36 GND mn15  l=0.13u w=0.26u m=1
M26 GND N_34 N_36 GND mn15  l=0.13u w=0.26u m=1
M27 N_9 N_8 VDD VDD mp15  l=0.13u w=0.54u m=1
M28 N_90 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M29 VDD SE N_5 VDD mp15  l=0.13u w=0.4u m=1
M30 N_8 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M31 N_90 D N_79 VDD mp15  l=0.13u w=0.58u m=1
M32 N_79 N_5 N_89 VDD mp15  l=0.13u w=0.26u m=1
M33 N_89 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M34 N_79 N_9 N_19 VDD mp15  l=0.13u w=0.58u m=1
M35 N_19 N_8 N_91 VDD mp15  l=0.13u w=0.26u m=1
M36 VDD N_25 N_91 VDD mp15  l=0.13u w=0.26u m=1
M37 VDD N_19 N_25 VDD mp15  l=0.13u w=0.69u m=1
M38 Q N_31 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 Q N_31 VDD VDD mp15  l=0.13u w=0.69u m=1
M40 QN N_24 VDD VDD mp15  l=0.13u w=0.48u m=1
M41 VDD N_24 QN VDD mp15  l=0.13u w=0.47u m=1
M42 QN N_24 VDD VDD mp15  l=0.13u w=0.43u m=1
M43 N_25 N_8 N_24 VDD mp15  l=0.13u w=0.69u m=1
M44 N_92 N_9 N_24 VDD mp15  l=0.13u w=0.26u m=1
M45 N_24 SN VDD VDD mp15  l=0.13u w=0.345u m=1
M46 VDD SN N_24 VDD mp15  l=0.13u w=0.345u m=1
M47 VDD N_24 N_31 VDD mp15  l=0.13u w=0.345u m=1
M48 VDD N_24 N_31 VDD mp15  l=0.13u w=0.345u m=1
M49 VDD N_39 N_92 VDD mp15  l=0.13u w=0.26u m=1
M50 N_39 N_35 N_31 VDDG mp15  l=0.13u w=0.26u m=1
M51 N_35 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M52 N_34 N_39 VDDG VDDG mp15  l=0.13u w=0.26u m=1
M53 N_39 RETN N_93 VDDG mp15  l=0.13u w=0.26u m=1
M54 N_93 N_34 VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrprb2
* SPICE INPUT		Tue Sep 18 13:29:57 2018	sdrprbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdrprbm
.subckt sdrprbm VDDG VDD GND QN Q SN RETN SI SE CK D
M1 N_6 SE GND GND mn15  l=0.13u w=0.26u m=1
M2 N_9 CK GND GND mn15  l=0.13u w=0.21u m=1
M3 GND N_9 N_7 GND mn15  l=0.13u w=0.19u m=1
M4 N_13 D N_12 GND mn15  l=0.13u w=0.36u m=1
M5 GND N_6 N_13 GND mn15  l=0.13u w=0.36u m=1
M6 N_16 SI GND GND mn15  l=0.13u w=0.26u m=1
M7 N_16 SE N_12 GND mn15  l=0.13u w=0.26u m=1
M8 N_17 N_9 N_12 GND mn15  l=0.13u w=0.36u m=1
M9 N_11 N_21 GND GND mn15  l=0.13u w=0.26u m=1
M10 N_17 N_7 N_11 GND mn15  l=0.13u w=0.26u m=1
M11 QN N_27 GND GND mn15  l=0.13u w=0.36u m=1
M12 N_19 N_27 GND GND mn15  l=0.13u w=0.26u m=1
M13 N_22 N_17 N_21 GND mn15  l=0.13u w=0.3u m=1
M14 GND N_19 Q GND mn15  l=0.13u w=0.36u m=1
M15 N_21 N_7 N_27 GND mn15  l=0.13u w=0.26u m=1
M16 N_29 N_9 N_27 GND mn15  l=0.13u w=0.26u m=1
M17 GND SN N_22 GND mn15  l=0.13u w=0.6u m=1
M18 N_29 N_32 N_22 GND mn15  l=0.13u w=0.26u m=1
M19 N_31 RETN GND GND mn15  l=0.13u w=0.26u m=1
M20 N_19 RETN N_32 GND mn15  l=0.13u w=0.26u m=1
M21 N_36 N_31 N_32 GND mn15  l=0.13u w=0.26u m=1
M22 GND N_32 N_34 GND mn15  l=0.13u w=0.26u m=1
M23 N_36 N_34 GND GND mn15  l=0.13u w=0.26u m=1
M24 VDD SE N_6 VDD mp15  l=0.13u w=0.4u m=1
M25 N_84 SE VDD VDD mp15  l=0.13u w=0.55u m=1
M26 N_84 D N_72 VDD mp15  l=0.13u w=0.55u m=1
M27 N_72 N_6 N_83 VDD mp15  l=0.13u w=0.26u m=1
M28 N_83 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M29 N_9 CK VDD VDD mp15  l=0.13u w=0.54u m=1
M30 N_7 N_9 VDD VDD mp15  l=0.13u w=0.49u m=1
M31 QN N_27 VDD VDD mp15  l=0.13u w=0.55u m=1
M32 N_19 N_27 VDD VDD mp15  l=0.13u w=0.4u m=1
M33 N_85 N_9 N_17 VDD mp15  l=0.13u w=0.26u m=1
M34 VDD N_21 N_85 VDD mp15  l=0.13u w=0.26u m=1
M35 VDD N_17 N_21 VDD mp15  l=0.13u w=0.4u m=1
M36 N_27 N_9 N_21 VDD mp15  l=0.13u w=0.4u m=1
M37 N_72 N_7 N_17 VDD mp15  l=0.13u w=0.55u m=1
M38 VDD N_19 Q VDD mp15  l=0.13u w=0.55u m=1
M39 N_86 N_7 N_27 VDD mp15  l=0.13u w=0.26u m=1
M40 N_27 SN VDD VDD mp15  l=0.13u w=0.4u m=1
M41 N_86 N_32 VDD VDD mp15  l=0.13u w=0.26u m=1
M42 N_31 RETN VDDG VDDG mp15  l=0.13u w=0.26u m=1
M43 N_87 RETN N_32 VDDG mp15  l=0.13u w=0.26u m=1
M44 N_19 N_31 N_32 VDDG mp15  l=0.13u w=0.26u m=1
M45 VDDG N_32 N_34 VDDG mp15  l=0.13u w=0.26u m=1
M46 N_87 N_34 VDDG VDDG mp15  l=0.13u w=0.26u m=1
.ends sdrprbm
