* 
* No part of this file can be released without the consent of SMIC.
*
* Note: SMIC recommends that users set VNTOL=1E-9 at .option for more smooth convergence.
*************************************************************************************************************
* 0.11um Mixed Signal 1P8M with MIM Salicide 1.2V/3.3V RF SPICE Model (for HSPICE only)  *
*************************************************************************************************************
** * release version    : 1.14
** * 
** * release date       : 03/30/2016
** * 
** * simulation tool    : Synopsys Star-HSPICE version C-2009.09 
** * 
*  Inductor   :
*
*        *-------------------------------------------------------------------------------------------------* 
*        | Inductor subckt |   diff_ind_rf   | diff_ind_rf_pgs | diff_ind_rf_psub   | diff_ind_rf_pgs_psub |
*        *-------------------------------------------------------------------------------------------------*
**********************************
* 0.11um differential Inductor *
**********************************
* 1=port1(M8), 2=port2(M8)
* R means inner redius; N means turns
* Spacing is fixed at 1.5um and width is fixed at 8um
.subckt diff_ind_rf 1 2 R=radius N=turns 
* inductor scalable model parameters
.param
+L00  = 'max((88.81e-12*pwr((R*1e+4),1.29)+12.90e-12)*pwr(N,2)+(128.0e-12*(R*1e+4)-59.23e-12),1e-12)'
+R00 = 'max((0.3257*pwr((R*1e+4),0.9274)+0.1961)*N+(0.09286*(R*1e+4)-0.3465),1e-3)'
+L01  = 'max((61.08e-12*pwr((R*1e+4),2.257)+58.39e-12)*N+(-12.82e-12*pwr((R*1e+4),-0.4249)-83.58e-12),1e-12)'
+COXM = 'max((31.31e-15*pwr((R*1e+4),0.707)+1.520e-15)*pwr(N,1.2)+(27.95e-15*(R*1e+4)-12.55e-15),1e-18)'
+RSM = 'max((58.77e+3*pwr((R*1e+6),-1)+13.65)*pwr(N,-1)+(1.091e+3*pwr((R*1e+6),-0.5028)+39.07),1e-3)'
+CSM    = 1e-15
+CPASS = 'max((15.97e-15*pwr((R*1e+4),1.171)+7.596e-15)*pwr(N,1.2)+(-13.35e-15*pwr((R*1e+4),2.0)-18.82e-15),1e-18)'
+COXI  = 'max((0.2715e-15*pwr((R*1e+4),1.341)+0.5962e-15)*pwr(N,2)+(23.74e-15*pwr((R*1e+4),1.5)+4.7e-15),1e-18)'
+RSI = 300  
+CSI    = 'max(2.0e-15*pwr(N,1.2)+(77.23e-15*pwr((R*1e+4),0.7531)),1e-18)'
+COXO  = 'COXI'
+RSO    = 'RSI-5.0'
+CSO    = 'CSI'
+kk = 'max((-0.1962*pwr((R*1e+6),0.1493)+0.4354),1e-3)'
* equivalent circuit
L00_rf  1 N1    'L00*(1+DL00_RF)' 
R00_rf  N1 NM   'R00*(1+DR00_RF)' tc1=3.69e-03
L01_rf  N1 N11  L01 
R01_rf  N11 NM  '2.0*R00*(1+DR00_RF)' tc1=3.69e-03
L10_rf  NM N2   'L00*(1+DL00_RF)'  
R10_rf  N2 2    'R00*(1+DR00_RF)' tc1=3.69e-03
L11_rf  N2 N21  L01
R11_rf  N21 2   '2.0*R00*(1+DR00_RF)' tc1=3.69e-03
COXM_rf  NM NSM COXM
RSM_rf  NSM 0   RSM  
CSM_rf  NSM 0   CSM
CPASS_rf  1 2   CPASS 
CCI_rf  1 NM    0.1e-15 
CCO_rf  NM 2    0.1e-15  
RCI_rf  NSI NSM 1e+6  
RCO_rf  NSM NSO 1e+6  
COXI_rf 1 NSI   COXI
RSI_rf  NSI 0   RSI  
CSI_rf  NSI 0   CSI 
COXO_rf 2 NSO   COXO
RSO_rf  NSO 0   RSO  
CSO_rf  NSO 0   CSO
K01 L10_rf L01_rf kk
K11 L00_rf L11_rf kk
K12 L00_rf L10_rf 0.85
.ends diff_ind_rf
*****************************************
* 0.11um differential Inductor with PGS *
*****************************************
* 1=port1(M8), 2=port2(M8)
* R means inner redius; N means turns
* Spacing is fixed at 1.5um and width is fixed at 8um
.subckt diff_ind_rf_pgs 1 2 R=radius N=turns 
* inductor scalable model parameters
.param
+L00  = 'max((88.81e-12*pwr((R*1e+4),1.29)+12.90e-12)*pwr(N,2)+(128.0e-12*(R*1e+4)-59.23e-12),1e-12)'
+R00 = 'max((0.3257*pwr((R*1e+4),0.9274)+0.1961)*N+(0.09286*(R*1e+4)-0.3465),1e-3)'
+L01  = 'max((61.08e-12*pwr((R*1e+4),2.257)+58.39e-12)*N+(-12.82e-12*pwr((R*1e+4),-0.4249)-83.58e-12),1e-12)'
+COXM = 'max(((31.31e-15*pwr((R*1e+4),0.707)+1.520e-15)*pwr(N,1.2)+(27.95e-15*(R*1e+4)-12.55e-15))*1.16,1e-18)'
+RSM = 10
+CSM    = 1e-15
+CPASS = 'max((15.97e-15*pwr((R*1e+4),1.171)+7.596e-15)*pwr(N,1.2)+(-13.35e-15*pwr((R*1e+4),2.0)-18.82e-15),1e-18)'
+COXI  = 'max(((0.2715e-15*pwr((R*1e+4),1.341)+0.5962e-15)*pwr(N,2)+(23.74e-15*pwr((R*1e+4),1.5)+4.7e-15))*0.95,1e-18)'
+RSI = 150  
+CSI    = 'max(2.0e-15*pwr(N,1.2)+(77.23e-15*pwr((R*1e+4),0.7531)),1e-18)'
+COXO  = 'COXI'
+RSO    = 'RSI-1.0'
+CSO    = 'CSI'
+kk = 'max((-0.1962*pwr((R*1e+6),0.1493)+0.4354),1e-3)'
* equivalent circuit
L00_rf  1 N1    'L00*(1+DL00_RF)' 
R00_rf  N1 NM   'R00*(1+DR00_RF)' tc1=3.69e-03
L01_rf  N1 N11  L01 
R01_rf  N11 NM  '2.0*R00*(1+DR00_RF)' tc1=3.69e-03
L10_rf  NM N2   'L00*(1+DL00_RF)'  
R10_rf  N2 2    'R00*(1+DR00_RF)' tc1=3.69e-03
L11_rf  N2 N21  L01
R11_rf  N21 2   '2.0*R00*(1+DR00_RF)' tc1=3.69e-03
COXM_rf  NM NSM COXM
RSM_rf  NSM 0   RSM  
CSM_rf  NSM 0   CSM
CPASS_rf  1 2   CPASS 
CCI_rf  1 NM    0.1e-15 
CCO_rf  NM 2    0.1e-15  
RCI_rf  NSI NSM 1e+6  
RCO_rf  NSM NSO 1e+6  
COXI_rf 1 NSI   COXI
RSI_rf  NSI 0   RSI  
CSI_rf  NSI 0   CSI 
COXO_rf 2 NSO   COXO
RSO_rf  NSO 0   RSO  
CSO_rf  NSO 0   CSO
K01 L10_rf L01_rf kk
K11 L00_rf L11_rf kk
K12 L00_rf L10_rf 0.85
.ends diff_ind_rf_pgs
****************************************************
* 0.11um differential Inductor with psub terminals *
****************************************************
* 1=port1(M8), 2=port2(M8)
* R means inner redius; N means turns
* Spacing is fixed at 1.5um and width is fixed at 8um
.subckt diff_ind_rf_psub 1 2 psub R=radius N=turns 
* inductor scalable model parameters
.param
+L00  = 'max((88.81e-12*pwr((R*1e+4),1.29)+12.90e-12)*pwr(N,2)+(128.0e-12*(R*1e+4)-59.23e-12),1e-12)'
+R00 = 'max((0.3257*pwr((R*1e+4),0.9274)+0.1961)*N+(0.09286*(R*1e+4)-0.3465),1e-3)'
+L01  = 'max((61.08e-12*pwr((R*1e+4),2.257)+58.39e-12)*N+(-12.82e-12*pwr((R*1e+4),-0.4249)-83.58e-12),1e-12)'
+COXM = 'max((31.31e-15*pwr((R*1e+4),0.707)+1.520e-15)*pwr(N,1.2)+(27.95e-15*(R*1e+4)-12.55e-15),1e-18)'
+RSM = 'max((58.77e+3*pwr((R*1e+6),-1)+13.65)*pwr(N,-1)+(1.091e+3*pwr((R*1e+6),-0.5028)+39.07),1e-3)'
+CSM    = 1e-15
+CPASS = 'max((15.97e-15*pwr((R*1e+4),1.171)+7.596e-15)*pwr(N,1.2)+(-13.35e-15*pwr((R*1e+4),2.0)-18.82e-15),1e-18)'
+COXI  = 'max((0.2715e-15*pwr((R*1e+4),1.341)+0.5962e-15)*pwr(N,2)+(23.74e-15*pwr((R*1e+4),1.5)+4.7e-15),1e-18)'
+RSI = 300  
+CSI    = 'max(2.0e-15*pwr(N,1.2)+(77.23e-15*pwr((R*1e+4),0.7531)),1e-18)'
+COXO  = 'COXI'
+RSO    = 'RSI-5.0'
+CSO    = 'CSI'
+kk = 'max((-0.1962*pwr((R*1e+6),0.1493)+0.4354),1e-3)'
* equivalent circuit
L00_rf  1 N1    'L00*(1+DL00_RF)' 
R00_rf  N1 NM   'R00*(1+DR00_RF)' tc1=3.69e-03
L01_rf  N1 N11  L01 
R01_rf  N11 NM  '2.0*R00*(1+DR00_RF)' tc1=3.69e-03
L10_rf  NM N2   'L00*(1+DL00_RF)'  
R10_rf  N2 2    'R00*(1+DR00_RF)' tc1=3.69e-03
L11_rf  N2 N21  L01
R11_rf  N21 2   '2.0*R00*(1+DR00_RF)' tc1=3.69e-03
COXM_rf  NM NSM COXM
RSM_rf  NSM psub   RSM  
CSM_rf  NSM psub   CSM
CPASS_rf  1 2   CPASS 
CCI_rf  1 NM    0.1e-15 
CCO_rf  NM 2    0.1e-15  
RCI_rf  NSI NSM 1e+6  
RCO_rf  NSM NSO 1e+6  
COXI_rf 1 NSI   COXI
RSI_rf  NSI psub   RSI  
CSI_rf  NSI psub   CSI 
COXO_rf 2 NSO   COXO
RSO_rf  NSO psub   RSO  
CSO_rf  NSO psub   CSO
K01 L10_rf L01_rf kk
K11 L00_rf L11_rf kk
K12 L00_rf L10_rf 0.85
.ends diff_ind_rf_psub
************************************************************
* 0.11um differential Inductor with PGS and psub terminals *
************************************************************
* 1=port1(M8), 2=port2(M8)
* R means inner redius; N means turns
* Spacing is fixed at 1.5um and width is fixed at 8um
.subckt diff_ind_rf_pgs_psub 1 2 psub R=radius N=turns 
* inductor scalable model parameters
.param
+L00  = 'max((88.81e-12*pwr((R*1e+4),1.29)+12.90e-12)*pwr(N,2)+(128.0e-12*(R*1e+4)-59.23e-12),1e-12)'
+R00 = 'max((0.3257*pwr((R*1e+4),0.9274)+0.1961)*N+(0.09286*(R*1e+4)-0.3465),1e-3)'
+L01  = 'max((61.08e-12*pwr((R*1e+4),2.257)+58.39e-12)*N+(-12.82e-12*pwr((R*1e+4),-0.4249)-83.58e-12),1e-12)'
+COXM = 'max(((31.31e-15*pwr((R*1e+4),0.707)+1.520e-15)*pwr(N,1.2)+(27.95e-15*(R*1e+4)-12.55e-15))*1.16,1e-18)'
+RSM = 10
+CSM    = 1e-15
+CPASS = 'max((15.97e-15*pwr((R*1e+4),1.171)+7.596e-15)*pwr(N,1.2)+(-13.35e-15*pwr((R*1e+4),2.0)-18.82e-15),1e-18)'
+COXI  = 'max(((0.2715e-15*pwr((R*1e+4),1.341)+0.5962e-15)*pwr(N,2)+(23.74e-15*pwr((R*1e+4),1.5)+4.7e-15))*0.95,1e-18)'
+RSI = 150  
+CSI    = 'max(2.0e-15*pwr(N,1.2)+(77.23e-15*pwr((R*1e+4),0.7531)),1e-18)'
+COXO  = 'COXI'
+RSO    = 'RSI-1.0'
+CSO    = 'CSI'
+kk = 'max((-0.1962*pwr((R*1e+6),0.1493)+0.4354),1e-3)'
* equivalent circuit
L00_rf  1 N1    'L00*(1+DL00_RF)' 
R00_rf  N1 NM   'R00*(1+DR00_RF)' tc1=3.69e-03
L01_rf  N1 N11  L01 
R01_rf  N11 NM  '2.0*R00*(1+DR00_RF)' tc1=3.69e-03
L10_rf  NM N2   'L00*(1+DL00_RF)'  
R10_rf  N2 2    'R00*(1+DR00_RF)' tc1=3.69e-03
L11_rf  N2 N21  L01
R11_rf  N21 2   '2.0*R00*(1+DR00_RF)' tc1=3.69e-03
COXM_rf  NM NSM COXM
RSM_rf  NSM psub   RSM  
CSM_rf  NSM psub   CSM
CPASS_rf  1 2   CPASS 
CCI_rf  1 NM    0.1e-15 
CCO_rf  NM 2    0.1e-15  
RCI_rf  NSI NSM 1e+6  
RCO_rf  NSM NSO 1e+6  
COXI_rf 1 NSI   COXI
RSI_rf  NSI psub   RSI  
CSI_rf  NSI psub   CSI 
COXO_rf 2 NSO   COXO
RSO_rf  NSO psub   RSO  
CSO_rf  NSO psub   CSO
K01 L10_rf L01_rf kk
K11 L00_rf L11_rf kk
K12 L00_rf L10_rf 0.85
.ends diff_ind_rf_pgs_psub


