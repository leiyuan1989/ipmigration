************************************************************************
* auCdl Netlist:
* 
* Library Name:  prima_sc180bcd_5v_9t_sch
* Top Cell Name: NAND2_X2
* View Name:     schematic
* Netlisted on:  Apr 22 13:37:41 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    NAND2_X2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2_X2 A1 A2 VDD VNW VPW VSS ZN
*.PININFO A1:I A2:I ZN:O VDD:B VNW:B VPW:B VSS:B
mM3 net3 A2 VSS VPW nch5 mr=1 l=600n w=2.42u nf=2
mM1 ZN A1 net3 VPW nch5 mr=1 l=600n w=2.42u nf=2
mM4 ZN A2 VDD VNW pch5 mr=1 l=500n w=3.48u nf=2
mM0 ZN A1 VDD VNW pch5 mr=1 l=500n w=3.48u nf=2
.ENDS

