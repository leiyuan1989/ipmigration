************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    DFFR_X1
* View Name:    schematic
************************************************************************

.SUBCKT DFFR_X1 CLK D Q RN VDD VSS
*.PININFO CLK:I D:I RN:I Q:O VDD:B VNW:B VPW:B VSS:B
mNM13 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 net2 clkp net16 VPW nch5 mr=1 l=600n w=220n nf=1
mM12 net4 net10 VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM9 net2 D net5 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM2 net17 RN VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM3 net16 net6 net17 VPW nch5 mr=1 l=600n w=220n nf=1
mM8 net5 clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM22 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM17 net7 clkn net4 VPW nch5 mr=1 l=600n w=220n nf=1
mM19 Q net10 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM10 net6 net2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM15 net10 net7 net3 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM14 net3 RN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM6 net6 clkp net7 VPW nch5 mr=1 l=600n w=1.21u nf=1
mPM13 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM1 net2 clkn net16 VNW pch5 mr=1 l=500n w=300n nf=1
mM13 net4 net10 VDD VNW pch5 mr=1 l=500n w=300n nf=1
mM4 net16 net6 VDD VNW pch5 mr=1 l=500n w=300n nf=1
mM18 Q net10 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM21 net8 clkp VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM16 net7 clkp net4 VNW pch5 mr=1 l=500n w=300n nf=1
mM11 net6 net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM5 net16 RN VDD VNW pch5 mr=1 l=500n w=300n nf=1
mM25 net10 net7 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM24 net10 RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM20 net2 D net8 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM7 net6 clkn net7 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM23 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
.ENDS
