//* 
//* No part of this file can be released without the consent of SMIC.
//*
//******************************************************************************************
//* 0.11um Mixed Signal 1P8M with MIM Salicide 1.2V/3.3V RF SPICE Model (for SPECTRE only) *
//******************************************************************************************
//*
//* Release version    : 1.14
//*
//* Release date       : 31/03/2013
//*
//* Simulation tool    : Cadence spectre V10.0
//*
//*
//*  MIM Capacitor   :
//*
//*        *------------------------------------------------------------------------------------------------------* 
//*        | 1fF/um^2 subckt   |  mim1_rf       |  mim1_shield_rf         | mim1_shield_rf_3t                     | 
//*        *------------------------------------------------------------------------------------------------------* 
//*        | 1.5fF/um^2 subckt |  mim15_rf      |  mim15_shield_rf        | mim15_rf_3t    | mim15_shield_rf_3t   | 
//*        *------------------------------------------------------------------------------------------------------* 
//*        | 2fF/um^2 subckt   |  mim2_rf_2mask |  mim2_shield_rf_2mask   | mim2_shield_rf_2mask_3t               |
//*        *------------------------------------------------------------------------------------------------------*
//*        | 3fF/um^2 subckt   |  mim3_rf                                                                         | 
//*        *------------------------------------------------------------------------------------------------------* 
simulator lang=spectre  insensitive=yes
//*******************************                  
//* 0.11um 1fF/um^2 MIM Capacitor
//*******************************
//* 1=port1, 2=port2
subckt mim1_rf (1 2)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
//*** mismatch paramters
parameters ac0 = 0.0384    
parameters cc0 = 1.2717 
parameters ar_c0 = ((lr*0.9)*(wr*0.9)*mr*1e12)  
parameters geo_fac=(1/sqrt(ar_c0))
parameters dmim1_mis_rf  = (ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//*** 
parameters c0_a = 0.971
parameters cvc1 = 8.03e-6            
parameters cvc2 = 3.74e-6  
parameters ctc1 = 4.088E-05 
//*parameters ar_c0 = ((lr*0.9)*(wr*0.9)*mr*1e12)  
parameters c0    = (c0_a*ar_c0)
parameters tcoef = (1.0+ctc1*(temp-25.0)) 
parameters cf_rf = c0*(1+dmim1_RF)*(1+dmim1_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
//* equivalent circuit
ls    (1 11)  inductor   l=max((0.1709-5.88E-06*(lr*0.9)*(wr*0.9)*1E12)*1E-9*(0.0095*pwr(lr*wr*0.81,-0.1852)), 1E-13)   m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))
rs    (11 22) resistor   r=max(189.3258/((lr*0.9)*(wr*0.9)*1E12)*(0.9985*exp(547415735.7484*lr*wr*0.81)), 1E-6)  m=mr
rsub1 (10 0)  resistor   r=max(3.0E+04-2.0*(lr*0.9)*(wr*0.9)*1E12, 1E-3) m=mr
csub1 (10 0)  capacitor  c=max((0.08*(lr*0.9)*1E6)*1E-15, 1E-18)   m=mr
cox1  (1 10)  capacitor  c=max((2.5E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)   m=mr
rsub2 (20 0)  resistor   r=max(4.88E+03-6.495E-3*(lr*0.9)*(wr*0.9)*1E12, 1E-3)  m=mr
csub2 (20 0)  capacitor  c=max((0.1*(lr*0.9)*1E6)*1E-15, 1E-18)           m=mr
cox2  (2 20)  capacitor  c=max((6.38E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)  m=mr
ends mim1_rf
//*********************


//****************************************************
//* 0.11um 1fF/um^2 MIM Capacitor with shielding layer
//****************************************************
//* 1=port1, 2=port2
subckt mim1_shield_rf (1 2)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
//*** mismatch paramters
parameters ac0 = 0.0384    
parameters cc0 = 1.2717
parameters ar_c0 = ((lr*0.9)*(wr*0.9)*mr*1e12)  
parameters geo_fac=(1/sqrt(ar_c0))
parameters dmim1_mis_rf  = (ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//***
parameters c0_a = 0.971
parameters cvc1 = 8.03e-6            
parameters cvc2 = 3.74e-6  
parameters ctc1 = 4.088E-05 
parameters c0    = (c0_a*ar_c0)
parameters tcoef = (1.0+ctc1*(temp-25.0)) 
parameters cf_rf = c0*(1+dmim1_shield_RF)*(1+dmim1_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
//* equivalent circuit
ls    (1 11)  inductor   l=max((0.1709-5.88E-06*(lr*0.9)*(wr*0.9)*1E12)*1E-9*(0.0095*pwr(lr*wr*0.81,-0.1852)), 1E-13)   m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))
rs    (11 22) resistor   r=max(189.3258/((lr*0.9)*(wr*0.9)*1E12)*(0.9985*exp(547415735.7484*lr*wr*0.81))*(1.9845*pwr((lr*0.9)*(wr*0.9),0.02675)), 1E-6) m=mr
rsub1 (10 0)  resistor   r=max(3.0E+04-2.0*(lr*0.9)*(wr*0.9)*1E12, 1E-3) m=mr
csub1 (10 0)  capacitor  c=max((0.08*(lr*0.9)*1E6)*1E-15, 1E-18)  m=mr
cox1  (1 10)  capacitor  c=max((2.5E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)   m=mr
rsub2 (20 0)  resistor   r=max((4.88E+03-6.495E-3*(lr*0.9)*(wr*0.9)*1E12)/(875777*pwr((lr*0.9)*(wr*0.9),0.38965)), 1E-3)   m=mr
csub2 (20 0)  capacitor  c=max((0.1*(lr*0.9)*1E6)*1E-15, 1E-18)  m=mr
cox2  (2 20)  capacitor  c=max((6.38E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15+(0.105*(lr*0.9)*(wr*0.9)*1E12+0.9)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)  m=mr
ends mim1_shield_rf


//****************************************************
//* 0.11um 1fF/um^2 MIM Capacitor with shielding layer (3-terminal)
//****************************************************
//* 1=port1, 2=port2
subckt mim1_shield_rf_3t (1 2 p)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
//*** mismatch paramters
parameters ac0 = 0.0384    
parameters cc0 = 1.2717
parameters ar_c0 = ((lr*0.9)*(wr*0.9)*mr*1e12)  
parameters geo_fac=(1/sqrt(ar_c0))
parameters dmim1_mis_rf  = (ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//***
parameters c0_a = 0.971
parameters cvc1 = 8.03e-6            
parameters cvc2 = 3.74e-6  
parameters ctc1 = 4.088E-05 
parameters c0    = (c0_a*ar_c0)
parameters tcoef = (1.0+ctc1*(temp-25.0)) 
parameters cf_rf = c0*(1+dmim1_shield_RF)*(1+dmim1_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
//* equivalent circuit
ls    (1 11)  inductor   l=max((0.1709-5.88E-06*(lr*0.9)*(wr*0.9)*1E12)*1E-9*(0.0095*pwr(lr*wr*0.81,-0.1852)), 1E-13)   m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))
rs    (11 22) resistor   r=max(189.3258/((lr*0.9)*(wr*0.9)*1E12)*(0.9985*exp(547415735.7484*lr*wr*0.81))*(1.9845*pwr((lr*0.9)*(wr*0.9),0.02675)), 1E-6) m=mr
rsub1 (10 p)  resistor   r=max(3.0E+04-2.0*(lr*0.9)*(wr*0.9)*1E12, 1E-3) m=mr
csub1 (10 p)  capacitor  c=max((0.08*(lr*0.9)*1E6)*1E-15, 1E-18)  m=mr
cox1  (1 10)  capacitor  c=max((2.5E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)   m=mr
rsub2 (20 p)  resistor   r=max((4.88E+03-6.495E-3*(lr*0.9)*(wr*0.9)*1E12)/(875777*pwr((lr*0.9)*(wr*0.9),0.38965)), 1E-3)   m=mr
csub2 (20 p)  capacitor  c=max((0.1*(lr*0.9)*1E6)*1E-15, 1E-18)  m=mr
cox2  (2 20)  capacitor  c=max((6.38E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15+(0.105*(lr*0.9)*(wr*0.9)*1E12+0.9)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)  m=mr
ends mim1_shield_rf_3t

//*********************************
//* 0.11um 1.5fF/um^2 MIM Capacitor
//*********************************
//* 1=port1, 2=port2
subckt mim15_rf (1 2)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
//*** mismatch paramters
parameters ac0 = 2.2793E-02    
parameters cc0 = 1.1757
parameters ar_c0 = ((lr*0.9)*(wr*0.9)*mr*1e12)  
parameters geo_fac=(1/sqrt(ar_c0))
parameters dmim15_mis_rf      = (ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//***
parameters c0_a = 1.449
parameters cvc1  = 9.68e-6            
parameters cvc2 = 6.72e-6   
parameters ctc1 = 3.758E-05
parameters c0    = (c0_a*ar_c0)
parameters tcoef = (1.0+ctc1*(temp-25.0))  
parameters cf_rf = c0*(1+dmim15_RF)*(1+dmim15_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
//* equivalent circuit
ls    (1 11)  inductor   l=max((0.1709-5.88E-06*(lr*0.9)*(wr*0.9)*1E12)*1E-9, 1E-13)  m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))
rs    (11 22) resistor   r=max(189.3258/((lr*0.9)*(wr*0.9)*1E12), 1E-6) m=mr
rsub1 (10 0)  resistor   r=max(3.0E+04-2.0*(lr*0.9)*(wr*0.9)*1E12, 1E-3) m=mr
csub1 (10 0)  capacitor  c=max((0.08*(lr*0.9)*1E6)*1E-15, 1E-18)   m=mr
cox1  (1 10)  capacitor  c=max((0.08*pwr(wr*lr*0.81*1e12,0.5)+0.02)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)  m=mr
rsub2 (20 0)  resistor   r=max(4.88E+03-6.495E-3*(lr*0.9)*(wr*0.9)*1E12, 1E-3)  m=mr
csub2 (20 0)  capacitor  c=max((0.1*(lr*0.9)*1E6)*1E-15, 1E-18)          m=mr
cox2  (2 20)  capacitor  c=max((0.2*pwr(wr*lr*0.81*1e12,0.5)+0.46)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)  m=mr
ends mim15_rf

//************************************************
//* 0.11um 1.5fF/um^2 MIM Capacitor (3-terminal)
//************************************************
//* 1=port1, 2=port2
subckt mim15_rf_3t (1 2 p)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
//*** mismatch paramters
parameters ac0 = 2.2793E-02    
parameters cc0 = 1.1757
parameters ar_c0 = ((lr*0.9)*(wr*0.9)*mr*1e12)  
parameters geo_fac=(1/sqrt(ar_c0))
parameters dmim15_mis_rf      = (ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//***
parameters c0_a = 1.449
parameters cvc1  = 9.68e-6            
parameters cvc2 = 6.72e-6   
parameters ctc1 = 3.758E-05
parameters c0    = (c0_a*ar_c0)
parameters tcoef = (1.0+ctc1*(temp-25.0))  
parameters cf_rf = c0*(1+dmim15_RF)*(1+dmim15_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
//* equivalent circuit
ls    (1 11)  inductor   l=max((0.1709-5.88E-06*(lr*0.9)*(wr*0.9)*1E12)*1E-9, 1E-13)  m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))
rs    (11 22) resistor   r=max(189.3258/((lr*0.9)*(wr*0.9)*1E12), 1E-6) m=mr
rsub1 (10 p)  resistor   r=max(3.0E+04-2.0*(lr*0.9)*(wr*0.9)*1E12, 1E-3) m=mr
csub1 (10 p)  capacitor  c=max((0.08*(lr*0.9)*1E6)*1E-15, 1E-18)   m=mr
cox1  (1 10)  capacitor  c=max((0.08*pwr(wr*lr*0.81*1e12,0.5)+0.02)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)  m=mr
rsub2 (20 p)  resistor   r=max(4.88E+03-6.495E-3*(lr*0.9)*(wr*0.9)*1E12, 1E-3)  m=mr
csub2 (20 p)  capacitor  c=max((0.1*(lr*0.9)*1E6)*1E-15, 1E-18)          m=mr
cox2  (2 20)  capacitor  c=max((0.2*pwr(wr*lr*0.81*1e12,0.5)+0.46)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)  m=mr
ends mim15_rf_3t

//******************************************************
//* 0.11um 1.5fF/um^2 MIM Capacitor with shielding layer
//******************************************************
//* 1=port1, 2=port2
subckt mim15_shield_rf (1 2)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
//*** mismatch paramters
parameters ac0 = 2.2793E-02    
parameters cc0 = 1.1757 
parameters ar_c0 = ((lr*0.9)*(wr*0.9)*mr*1e12)  
parameters geo_fac=(1/sqrt(ar_c0))
parameters dmim15_mis_rf      = (ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//***  
parameters c0_a = 1.449
parameters cvc1  = 9.68e-6            
parameters cvc2 = 6.72e-6   
parameters ctc1 = 3.758E-05
parameters c0    = (c0_a*ar_c0)
parameters tcoef = (1.0+ctc1*(temp-25.0))  
parameters cf_rf = c0*(1+dmim15_shield_RF)*(1+dmim15_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
//* equivalent circuit
ls    (1 11)  inductor   l=max((0.1709-5.88E-06*(lr*0.9)*(wr*0.9)*1E12)*1E-9, 1E-13)    m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))    
rs    (11 22) resistor   r=max(189.3258/((lr*0.9)*(wr*0.9)*1E12)*(1.9845*pwr((lr*0.9)*(wr*0.9),0.02675)), 1E-6) m=mr
rsub1 (10 0)  resistor   r=max(3.0E+04-2.0*(lr*0.9)*(wr*0.9)*1E12, 1E-3) m=mr
csub1 (10 0)  capacitor  c=max((0.08*(lr*0.9)*1E6)*1E-15, 1E-18)   m=mr
cox1  (1 10)  capacitor  c=max((0.08*pwr(wr*lr*0.81*1e12,0.5)+0.02)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)   m=mr
rsub2 (20 0)  resistor   r=max((4.88E+03-6.495E-3*(lr*0.9)*(wr*0.9)*1E12)/(613044*pwr((lr*0.9)*(wr*0.9),0.38965)), 1E-3)    m=mr
csub2 (20 0)  capacitor  c=max((0.1*(lr*0.9)*1E6)*1E-15, 1E-18) m=mr
cox2  (2 20)  capacitor  c=max((6.38E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15+(0.105*(lr*0.9)*(wr*0.9)*1E12+0.9)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)  m=mr
ends mim15_shield_rf

//*********************************************************************
//* 0.11um 1.5fF/um^2 MIM Capacitor with shielding layer (3-terminal)
//*********************************************************************
//* 1=port1, 2=port2
subckt mim15_shield_rf_3t (1 2 p)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
//*** mismatch paramters
parameters ac0 = 2.2793E-02    
parameters cc0 = 1.1757 
parameters ar_c0 = ((lr*0.9)*(wr*0.9)*mr*1e12)  
parameters geo_fac=(1/sqrt(ar_c0))
parameters dmim15_mis_rf      = (ac0*pwr(geo_fac,cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//***  
parameters c0_a = 1.449
parameters cvc1  = 9.68e-6            
parameters cvc2 = 6.72e-6   
parameters ctc1 = 3.758E-05
parameters c0    = (c0_a*ar_c0)
parameters tcoef = (1.0+ctc1*(temp-25.0))  
parameters cf_rf = c0*(1+dmim15_shield_RF)*(1+dmim15_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
//* equivalent circuit
ls    (1 11)  inductor   l=max((0.1709-5.88E-06*(lr*0.9)*(wr*0.9)*1E12)*1E-9, 1E-13)    m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))    
rs    (11 22) resistor   r=max(189.3258/((lr*0.9)*(wr*0.9)*1E12)*(1.9845*pwr((lr*0.9)*(wr*0.9),0.02675)), 1E-6) m=mr
rsub1 (10 p)  resistor   r=max(3.0E+04-2.0*(lr*0.9)*(wr*0.9)*1E12, 1E-3) m=mr
csub1 (10 p)  capacitor  c=max((0.08*(lr*0.9)*1E6)*1E-15, 1E-18)   m=mr
cox1  (1 10)  capacitor  c=max((0.08*pwr(wr*lr*0.81*1e12,0.5)+0.02)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)   m=mr
rsub2 (20 p)  resistor   r=max((4.88E+03-6.495E-3*(lr*0.9)*(wr*0.9)*1E12)/(613044*pwr((lr*0.9)*(wr*0.9),0.38965)), 1E-3)    m=mr
csub2 (20 p)  capacitor  c=max((0.1*(lr*0.9)*1E6)*1E-15, 1E-18) m=mr
cox2  (2 20)  capacitor  c=max((6.38E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15+(0.105*(lr*0.9)*(wr*0.9)*1E12+0.9)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)  m=mr
ends mim15_shield_rf_3t

//*********************************
//* 0.11um 2.0fF/um^2 MIM Capacitor
//*********************************
//* 1=port1, 2=port2
subckt mim2_rf_2mask (1 2)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
// *** mismatch paramters 
parameters ac0 = 0.132900035    
parameters cc0 = 0.000206611
parameters dmim2_2mask_mis_rf = ((ac0/c0+cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//***
parameters  c0_a = 2.1  
parameters  cvc1 = -6.119607E-05 
parameters  cvc2 = 2.660293E-05  
parameters  ctc1 = 3.25876E-05  
parameters  ar_c0= (lr*0.9)*(wr*0.9)*mr*1e12  
parameters  c0   = c0_a*ar_c0
parameters  tcoef= 1.00+ctc1*(temp-25.00)
// *
parameters Ls_rf     = max((2.09*pwr((lr*0.9)*(wr*0.9)*1e12,-1.35)+4.1e-6*(lr*0.9)*(wr*0.9)*1e12+0.0061)*1e-9,1e-15)
parameters Cf_rf     = c0*(1+dmim2_RF_2mask)*(1+dmim2_2mask_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
parameters Rs_rf     = max(43.7*pwr((lr*0.9)*(wr*0.9)*1e12,-0.83)+0.00035*(lr*0.9)*(wr*0.9)*1e12,1e-6)
parameters Rsub1_rf  = max(31950*pwr((lr*0.9)*(wr*0.9)*1E12,-0.021), 1E-3)
parameters Csub1_rf  = max((0.08*sqrt((wr*0.9)*(lr*0.9)*1E12))*1E-15, 1E-18)
parameters Cox1_rf   = max((2.5E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)
parameters Rsub2_rf  = max(4929.7*pwr((lr*0.9)*(wr*0.9)*1E12,-0.0946), 1E-3)
parameters Csub2_rf  = max((0.1*sqrt((wr*0.9)*(lr*0.9)*1E12))*1E-15, 1E-18)
parameters Cox2_rf   = max((6.38E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)
//* equivalent circuit
ls    (1 11)  inductor   l=ls_rf      m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))
rs    (11 22) resistor   r=rs_rf      m=mr
rsub1 (10 0)  resistor   r=rsub1_rf   m=mr
csub1 (10 0)  capacitor  c=csub1_rf   m=mr
cox1  (1 10)  capacitor  c=cox1_rf    m=mr
rsub2 (20 0)  resistor   r=rsub2_rf   m=mr
csub2 (20 0)  capacitor  c=csub2_rf   m=mr
cox2  (2 20)  capacitor  c=cox2_rf    m=mr
ends mim2_rf_2mask

//******************************************************
//* 0.11um 2.0fF/um^2 MIM Capacitor with shielding layer
//******************************************************
//* 1=port1, 2=port2
subckt mim2_shield_rf_2mask (1 2)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
// *** mismatch paramters 
parameters ac0 = 0.132900035    
parameters cc0 = 0.000206611
parameters dmim2_2mask_mis_rf = ((ac0/c0+cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//***
parameters  c0_a = 2.1  
parameters  cvc1 = -6.119607E-05 
parameters  cvc2 = 2.660293E-05  
parameters  ctc1 = 3.25876E-05  
parameters ar_c0 = (lr*0.9)*(wr*0.9)*mr*1e12  
parameters c0    = c0_a*ar_c0
parameters tcoef = 1.00+ctc1*(temp-25.00)
// *
parameters Ls_rf     = max((1.23*pwr((lr*0.9)*(wr*0.9)*1e12,-1.25)+4.1e-6*(lr*0.9)*(wr*0.9)*1e12+0.0061)*1e-9,1e-15)
parameters Cf_rf     = c0*(1+dmim2_shield_RF_2mask)*(1+dmim2_2mask_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
parameters Rs_rf     = max(43.7*pwr((lr*0.9)*(wr*0.9)*1e12,-0.83)+0.00019*(lr*0.9)*(wr*0.9)*1e12,1e-6)
parameters Rsub1_rf  = max(31950*pwr((lr*0.9)*(wr*0.9)*1E12,-0.021), 1E-3)
parameters Csub1_rf  = max((0.08*sqrt((wr*0.9)*(lr*0.9)*1E12))*1E-15, 1E-18)
parameters Cox1_rf   = max((2.5E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)
parameters Rsub2_rf  = max(19.557*pwr((lr*0.9)*(wr*0.9)*1E12,-0.3473), 1E-3)
parameters Csub2_rf  = max((0.1*sqrt((wr*0.9)*(lr*0.9)*1E12))*1E-15, 1E-18)
parameters Cox2_rf   = max((2.9453*pwr((lr*0.9)*(wr*0.9)*1E12,0.87)+20.224)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)
//* equivalent circuit
ls    (1 11)  inductor   l=ls_rf      m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))
rs    (11 22) resistor   r=rs_rf      m=mr
rsub1 (10 0)  resistor   r=rsub1_rf   m=mr
csub1 (10 0)  capacitor  c=csub1_rf   m=mr
cox1  (1 10)  capacitor  c=cox1_rf    m=mr
rsub2 (20 0)  resistor   r=rsub2_rf   m=mr
csub2 (20 0)  capacitor  c=csub2_rf   m=mr
cox2  (2 20)  capacitor  c=cox2_rf    m=mr
ends mim2_shield_rf_2mask
//*
//******************************************************
//* 0.11um 2.0fF/um^2 MIM Capacitor with shielding layer (3-terminal)
//******************************************************
//* 1=port1, 2=port2
subckt mim2_shield_rf_2mask_3t (1 2 p)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
// *** mismatch paramters 
parameters ac0 = 0.132900035    
parameters cc0 = 0.000206611
parameters dmim2_2mask_mis_rf = ((ac0/c0+cc0)*sigma_mis_mim_rf*mismod_mim_rf)
//***
parameters  c0_a = 2.1  
parameters  cvc1 = -6.119607E-05 
parameters  cvc2 = 2.660293E-05  
parameters  ctc1 = 3.25876E-05  
parameters ar_c0 = (lr*0.9)*(wr*0.9)*mr*1e12  
parameters c0    = c0_a*ar_c0
parameters tcoef = 1.00+ctc1*(temp-25.00)
// *
parameters Ls_rf     = max((1.23*pwr((lr*0.9)*(wr*0.9)*1e12,-1.25)+4.1e-6*(lr*0.9)*(wr*0.9)*1e12+0.0061)*1e-9,1e-15)
parameters Cf_rf     = c0*(1+dmim2_shield_RF_2mask)*(1+dmim2_2mask_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
parameters Rs_rf     = max(43.7*pwr((lr*0.9)*(wr*0.9)*1e12,-0.83)+0.00019*(lr*0.9)*(wr*0.9)*1e12,1e-6)
parameters Rsub1_rf  = max(31950*pwr((lr*0.9)*(wr*0.9)*1E12,-0.021), 1E-3)
parameters Csub1_rf  = max((0.08*sqrt((wr*0.9)*(lr*0.9)*1E12))*1E-15, 1E-18)
parameters Cox1_rf   = max((2.5E-03*(lr*0.9)*(wr*0.9)*1E12)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18)
parameters Rsub2_rf  = max(19.557*pwr((lr*0.9)*(wr*0.9)*1E12,-0.3473), 1E-3)
parameters Csub2_rf  = max((0.1*sqrt((wr*0.9)*(lr*0.9)*1E12))*1E-15, 1E-18)
parameters Cox2_rf   = max((2.9453*pwr((lr*0.9)*(wr*0.9)*1E12,0.87)+20.224)*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18)
//* equivalent circuit
ls    (1 11)  inductor   l=ls_rf      m=mr
cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))
rs    (11 22) resistor   r=rs_rf      m=mr
rsub1 (10 p)  resistor   r=rsub1_rf   m=mr
csub1 (10 p)  capacitor  c=csub1_rf   m=mr
cox1  (1 10)  capacitor  c=cox1_rf    m=mr
rsub2 (20 p)  resistor   r=rsub2_rf   m=mr
csub2 (20 p)  capacitor  c=csub2_rf   m=mr
cox2  (2 20)  capacitor  c=cox2_rf    m=mr
ends mim2_shield_rf_2mask_3t
//*
//******************************************************************************** 
//            0.11um 3fF/um^2 stacked MIM Capacitor                              * 
//********************************************************************************
//* 1=port1, 2=port2
subckt mim3_rf (1 2)
//* mim capacitor scalable model parameters
parameters lr=l wr=w mr=m mismod_mim_rf=0 xm=8
// *** mismatch paramters
parameters  ac0 = 0.3305    
parameters  cc0 = 0.000152
parameters dmim3_mis_rf = ((ac0/c0+cc0)*sigma_mis_mim_rf*mismod_mim_rf)
// *** low frequency capacitor
parameters  c0_a = 3.01368807   
parameters  c0_p = 0.44926463
parameters  cvc1 = 2.37303251E-06  
parameters  cvc2 = 8.08656805E-06  
parameters  ctc1 = 3.92547475E-05  
parameters  ctc2 = 1.26746609E-07
parameters  ar_c0 = ((lr*0.9)*(wr*0.9)*mr*1e12 ) 
parameters  pe_c0 = (2*((lr*0.9)+(wr*0.9))*mr*1e6)
parameters  c0    = (c0_a*ar_c0+c0_p*pe_c0)
parameters  tcoef = (1.0+ctc1*(temp-25.0)+ctc2*(temp-25.0)*(temp-25.0))
//*
parameters cf_rf = c0*(1+dmim3_rf)*(1+dmim3_mis_rf)*1e-15*(1+(19.318*pwr(sqrt(wr*lr*1e12),-0.7578)*0.0001*(xm-8)))
//* equivalent circuit
ls    (1 11)  inductor   l=max((1.13*pwr((lr*0.9)*(wr*0.9)*1E12,-1.4)+0.005)*1E-9, 1E-12) m=mr
//cf    (22 2)  capacitor  c=cf_rf*tcoef*(1.0+v(22,2)*(cvc1+cvc2*v(22,2)))
cf    (22 2)  capacitor  c=c0*1e-15
rs    (11 22) resistor   r=max(65*pwr((lr*0.9)*(wr*0.9)*1E12,-1)+0.53, 1E-6) m=mr
rsub1 (10 0)  resistor   r=max(1887.8*pwr((lr*0.9)*(wr*0.9)*1E12,-0.3764), 1E-3) m=mr
csub1 (10 0)  capacitor  c=max(73.335*pwr((lr*0.9)*(wr*0.9)*1E12,-0.6825)*1E-15, 1E-18) m=mr
cox1  (1 10)  capacitor  c=max((0.0172*(lr*0.9)*(wr*0.9)*1E12+0.2275)*1E-15*(1-(0.0049*log(sqrt(wr*lr*1e12))+0.0201)*(xm-8)), 1E-18) m=mr
rsub2 (20 0)  resistor   r=max(1000, 1E-3) m=mr
csub2 (20 0)  capacitor  c=max(1*1E-15, 1E-18) m=mr
cox2  (2 20)  capacitor  c=max(0.0098*2*((lr*0.9)+(wr*0.9))*1E6*1E-15*(1-(0.0442*log(sqrt(wr*lr*1e12))-0.0019)*(xm-8)), 1E-18) m=mr
ends mim3_rf
//*
