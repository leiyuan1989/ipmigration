*  
* No part of this file can be released without the consent of SMIC. 
**************************************************************************************************** 
* SMIC 0.11um Radio Frequency 1P8M(1P7M, 1P6M, 1P5M) Top Metal SPICE Resistor model (for HSPICE only) * 
**************************************************************************************************** 
* 
* Release version    : 1.14
* 
* Release date       : 03/30/2016
* 
* Simulation tool    : Synopsys Star-HSPICE version 2006.9 
* 
*   Resistor         : 
*        *------------------------------------------*  
*        |       Resistor Type       | 		    |
*        |==========================================|         
*        |          Metal 8(TM2)     |    rtm2_rf   | 
*        |------------------------------------------| 
*        |          ALPA             |    ralpa_rf  | 
*        *------------------------------------------*  
*
*   The valid temperature range is from -40c to 125c
*
****************************************************************** 
*                         Resistor Model                         * 
******************************************************************  

****************************************************************** 
*                      Metal 8(TM2) resistance                   *  
****************************************************************** 
.subckt rtm2_rf n2 n1 sub l=lr w=wr   
.param  
+rsh       = '7E-03+DRSH_TM2_RF'       rtc1 = 3.69E-03     rtc2 = -1.80E-08   dw = '3.2167E-08+DDW_TM2_RF'
+jc1a      = -5.7371E-03               jc1b = 5.7922E-05
+jc2a      = 5.785E-05                 jc2b = 9.0221E-07
+rvc1      = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l'          
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+dl        = '3.2167E-08+DDW_TM2_RF'     weff = 'w*0.9-2*dw'     leff = 'l*0.9-2*dl' 
+cox       = '5.53E-06+DCOX_TM2_RF'               capsw    = '1.1540E-10+DCAPSW_TM2_RF'
C1 n2 sub 'cox*weff*leff/2+capsw*weff+capsw*leff'    
R1 n2 n1 'rsh*leff/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*leff/2+capsw*weff+capsw*leff'  
.ends rtm2_rf

****************************************************************** 
*                      ALPA resistance                           *  
****************************************************************** 
.subckt ralpa_rf n2 n1 sub l=lr w=wr   
.param  
+rsh       = '0.0231+DRSH_ALPA_RF'       rtc1 = 3.8865E-03   rtc2 = 5.5735E-08   dw = '-5.79E-08+DDW_ALPA_RF'
+jc1a      = 1.9362E-05              jc1b = -9.0694E-08
+jc2a      = 1.6459E-05              jc2b = 2.523E-07
+rvc1      = 'jc1a+jc1b/l'           rvc2   = '(jc2a+jc2b/l)/l'          
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+dl        = '-5.79E-08+DDW_ALPA_RF'     weff = 'w*0.9-2*dw'     leff = 'l*0.9-2*dl' 
+cox       = '3.53E-06+DCOX_ALPA_RF'               capsw    = '4.649E-11+DCAPSW_ALPA_RF'
C1 n2 sub 'cox*weff*leff/2+capsw*weff+capsw*leff'    
R1 n2 n1 'rsh*leff/weff*tcoef(temper)*min(1.0+rvc1*abs(v(n2,n1))+rvc2*v(n2,n1)*v(n2,n1), 1.1)'
C2 n1 sub 'cox*weff*leff/2+capsw*weff+capsw*leff'  
.ends ralpa_rf
