
.SUBCKT SDFFHQNX1MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net71 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net48 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 pm nmsi net60 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFHQNX2MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net71 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net48 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.6e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 pm nmsi net60 VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT SDFFHQNX4MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=2.9e-07
MXN2 net71 cn VSS VPW n12 l=1.3e-07 w=2.9e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.2e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=5e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net48 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP3 pm nmsi net60 VNW p12 l=1.3e-07 w=3.5e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=6.1e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFHQNX8MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=3.4e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3e-07
MXN3 net71 cn VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=5.4e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g2_MXNA1_2 s bm VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=4.2e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.8e-07
MXP4 net48 c cn VNW p12 l=1.3e-07 w=4.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.3e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=6.5e-07
MXP5 pm nmsi net60 VNW p12 l=1.3e-07 w=6.5e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.5e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=6e-07
mX_g2_MXPA1_2 s bm VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFHQX1MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.1e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=3.3e-07
MXN1 net54 cn VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.7e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net065 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.6e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=4e-07
MXP2 pm nmsi net71 VNW p12 l=1.3e-07 w=4e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.3e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
.ends


.SUBCKT SDFFHQX2MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=1.9e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=3.1e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=4.8e-07
MXN2 net54 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP3 net065 c cn VNW p12 l=1.3e-07 w=4.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP4 pm nmsi net71 VNW p12 l=1.3e-07 w=5.9e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
.ends


.SUBCKT SDFFHQX4MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=3.2e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.5e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.4e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=6.9e-07
MXN3 net54 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP5 net065 c cn VNW p12 l=1.3e-07 w=7.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=6.7e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP6 pm nmsi net71 VNW p12 l=1.3e-07 w=8e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT SDFFHQX8MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=5.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.5e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.4e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=6.9e-07
MXN3 net54 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.9e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP5 net065 c cn VNW p12 l=1.3e-07 w=7.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=6.7e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=5e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=8.3e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP6 pm nmsi net71 VNW p12 l=1.3e-07 w=8e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT SDFFHX1MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.3e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net0107 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 net104 cn VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 net079 c cn VNW p12 l=1.3e-07 w=4.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.8e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.8e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 nmsi SI net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP10 pm nmsi net087 VNW p12 l=1.3e-07 w=4.4e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.9e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=3e-07 nf=2
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
*mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFHX2MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=3.2e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net0107 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=5.1e-07
MXN7 net104 cn VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP13 net079 c cn VNW p12 l=1.3e-07 w=4.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.9e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 nmsi SI net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP12 pm nmsi net087 VNW p12 l=1.3e-07 w=6.2e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g6_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.1e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT SDFFHX4MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.4e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=2.9e-07
MXN8 net0107 SE VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=7e-07
MXN9 net104 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 net079 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=7e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP14 nmsi SI net76 VNW p12 l=1.3e-07 w=3.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 pm nmsi net087 VNW p12 l=1.3e-07 w=8.7e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g6_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT SDFFHX8MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.4e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=2.9e-07
MXN8 net0107 SE VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=7e-07
MXN9 net104 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 net079 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=7e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP14 nmsi SI net76 VNW p12 l=1.3e-07 w=3.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 pm nmsi net087 VNW p12 l=1.3e-07 w=8.7e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g6_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT SDFFNHX1MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmsi SI n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 n1 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=4.3e-07
MXN5 net58 cn VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=4e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP2 net87 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP8 p1 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmsi SI p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=6.8e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP10 pm nmsi net93 VNW p12 l=1.3e-07 w=3.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=4.8e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=3.1e-07 nf=2
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
*mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFNHX2MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmsi SI n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 n1 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=6.1e-07
MXN1 net58 cn VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP2 net87 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP8 p1 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmsi SI p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=8.4e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP5 pm nmsi net93 VNW p12 l=1.3e-07 w=4.6e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFNHX4MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.7e-07
MXN5 nmsi SI net058 VPW n12 l=1.3e-07 w=2.7e-07
MXN7 net058 SE VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=4.6e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=5.4e-07
MXN1 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MX_t3_2 pm nmsi net58 VPW n12 l=1.3e-07 w=5.4e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI59_MXNOE_2 nm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP10 net87 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.3e-07
MXP14 p1 nmse VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP9 nmsi SI p1 VNW p12 l=1.3e-07 w=3.3e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g10_MXPA1_2 cn net185 VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP13 pm nmsi net93 VNW p12 l=1.3e-07 w=6.9e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN_2 nm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g1_MXPA1_3 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFNHX8MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=4.7e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.1e-07
MXN7 nmsi SI n1 VPW n12 l=1.3e-07 w=5.1e-07
MXN6 n1 SE VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=5e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=7.4e-07
MXN1 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MX_t3_2 pm nmsi net58 VPW n12 l=1.3e-07 w=7.4e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI59_MXNOE_2 nm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP14 net87 cn c VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.5e-07
MXP8 p1 nmse VDD VNW p12 l=1.3e-07 w=3.4e-07
MXP15 nmsi SI p1 VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=7.2e-07
mX_g10_MXPA1_2 cn net185 VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP13 pm nmsi net93 VNW p12 l=1.3e-07 w=6.9e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.7e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN_2 nm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFNSRHX1MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net0207 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net0207 VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MX_t30 nmsi SI net172 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 net172 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS SN net163 VPW n12 l=1.3e-07 w=4.3e-07
MXN17 net163 cn net160 VPW n12 l=1.3e-07 w=4.3e-07
MX_t26 pm nmsi net160 VPW n12 l=1.3e-07 w=4.3e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 net0106 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t12 net0106 pm net166 VPW n12 l=1.3e-07 w=4.5e-07
MXN19 VSS RN net166 VPW n12 l=1.3e-07 w=4.5e-07
MXN20 net0106 nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE bm c net0106 VPW n12 l=1.3e-07 w=4e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net181 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net181 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 net0207 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net080 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net080 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn net0207 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP16 nmsi SI net117 VNW p12 l=1.3e-07 w=2.3e-07
MX_t32 net117 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP17 pm nmsi net0125 VNW p12 l=1.3e-07 w=3.3e-07
MX_t24 net0125 c VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI23_MXPA1 XI23_p1 net0106 VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 net0106 pm VDD VNW p12 l=1.3e-07 w=4.8e-07
MXP18 net111 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net0106 RN net111 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net0106 VNW p12 l=1.3e-07 w=4.8e-07
MXP21 bm nmset net126 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 net126 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP24 bm c net132 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net132 nmset net135 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net135 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT SDFFNSRHX2MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net261 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net261 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MX_t30 nmsi SI net168 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 net168 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN26 VSS SN net149 VPW n12 l=1.3e-07 w=6.1e-07
MXN25 net149 cn net153 VPW n12 l=1.3e-07 w=6.1e-07
MX_t26 pm nmsi net153 VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 net129 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN27 net129 pm net145 VPW n12 l=1.3e-07 w=6.3e-07
MXN28 VSS RN net145 VPW n12 l=1.3e-07 w=6.3e-07
MXN20 net129 nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE bm c net129 VPW n12 l=1.3e-07 w=5.5e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net261 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net109 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net109 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn net261 VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP16 nmsi SI net91 VNW p12 l=1.3e-07 w=2.3e-07
MX_t32 net91 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP25 pm nmsi net83 VNW p12 l=1.3e-07 w=4.6e-07
MX_t24 net83 c VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI23_MXPA1 XI23_p1 net129 VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 net129 pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP18 net103 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net129 RN net103 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net129 VNW p12 l=1.3e-07 w=6.7e-07
MXP28 bm nmset net79 VNW p12 l=1.3e-07 w=2.8e-07
MXP20 net79 RN VDD VNW p12 l=1.3e-07 w=2.8e-07
MXP24 bm c net123 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net123 nmset net119 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net119 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFNSRHX4MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net261 CKN VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net261 VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.7e-07
MX_t30 nmsi SI net168 VPW n12 l=1.3e-07 w=2.7e-07
MXN29 net168 SE VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN31 VSS SN net149 VPW n12 l=1.3e-07 w=7.6e-07
MXN30 net149 cn net153 VPW n12 l=1.3e-07 w=7.6e-07
MX_t26 pm nmsi net153 VPW n12 l=1.3e-07 w=7.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 net129 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN27 net129 pm net145 VPW n12 l=1.3e-07 w=8.4e-07
MXN32 VSS RN net145 VPW n12 l=1.3e-07 w=8.4e-07
MXN20 net129 nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI74_MXNOE bm c net129 VPW n12 l=1.3e-07 w=5.5e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net261 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net109 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP29 net109 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 cn net261 VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.2e-07
MXP30 nmsi SI net91 VNW p12 l=1.3e-07 w=3.3e-07
MX_t32 net91 nmse VDD VNW p12 l=1.3e-07 w=3.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP31 pm nmsi net83 VNW p12 l=1.3e-07 w=6.9e-07
MX_t24 net83 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI23_MXPA1 XI23_p1 net129 VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t10_2 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP18 net103 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net129 RN net103 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net129 VNW p12 l=1.3e-07 w=6.7e-07
MXP32 bm nmset net79 VNW p12 l=1.3e-07 w=3.6e-07
MXP20 net79 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP24 bm c net123 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net123 nmset net119 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net119 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFNSRHX8MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net261 CKN VSS VPW n12 l=1.3e-07 w=4.7e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net261 VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g10_MXNA1_2 cn net261 VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.4e-07
MX_t30 nmsi SI net168 VPW n12 l=1.3e-07 w=5.1e-07
MXN33 net168 SE VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN31 VSS SN net149 VPW n12 l=1.3e-07 w=7.6e-07
MXN30 net149 cn net153 VPW n12 l=1.3e-07 w=7.6e-07
MX_t26 pm nmsi net153 VPW n12 l=1.3e-07 w=7.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI23_MXNA1 XI23_n1 net129 VSS VPW n12 l=1.3e-07 w=2.5e-07
MXN27 net129 pm net145 VPW n12 l=1.3e-07 w=8.7e-07
MXN34 VSS RN net145 VPW n12 l=1.3e-07 w=8.7e-07
MXN20 net129 nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI74_MXNOE bm c net129 VPW n12 l=1.3e-07 w=5.5e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=3e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net261 CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MX_t4 net109 CKN VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP33 net109 cn c VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 cn net261 VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g10_MXPA1_2 cn net261 VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=1.03e-06
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=5.8e-07
MXP34 nmsi SI net91 VNW p12 l=1.3e-07 w=5.6e-07
MX_t32 net91 nmse VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=3.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP31 pm nmsi net83 VNW p12 l=1.3e-07 w=6.9e-07
MX_t24 net83 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI23_MXPA1 XI23_p1 net129 VDD VNW p12 l=1.3e-07 w=3.1e-07
MX_t10 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t10_2 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP18 net103 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net129 RN net103 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net129 VNW p12 l=1.3e-07 w=6.7e-07
MXP35 bm nmset net79 VNW p12 l=1.3e-07 w=3.5e-07
MXP20 net79 RN VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP24 bm c net123 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net123 nmset net119 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net119 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQNX1MTR QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net108 SE net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 VSS SI net108 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net111 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net129 D net111 VPW n12 l=1.3e-07 w=1.8e-07
MX_t1 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE pm c XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.7e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net69 nmse net65 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net65 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net68 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net69 D net68 VNW p12 l=1.3e-07 w=3.8e-07
MXP5 pm c net69 VNW p12 l=1.3e-07 w=3.8e-07
mXI1_MXPOEN pm cn XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFQNX2MTR QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net108 SE net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 VSS SI net108 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net111 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net129 D net111 VPW n12 l=1.3e-07 w=1.8e-07
MX_t1 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE pm c XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.7e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP6 net69 nmse net65 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net65 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net68 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net69 D net68 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 pm c net69 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN pm cn XI1_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQNX4MTR QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net108 SE net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 VSS SI net108 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net111 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net129 D net111 VPW n12 l=1.3e-07 w=1.8e-07
MX_t1 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE pm c XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.7e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP6 net69 nmse net65 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net65 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net68 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net69 D net68 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 pm c net69 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN pm cn XI1_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQX1MTR Q VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net064 SE net055 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 VSS SI net064 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net059 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net055 D net059 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm cn net055 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE pm c XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net105 m VSS VPW n12 l=1.3e-07 w=2.8e-07
MX_t12 ns c net105 VPW n12 l=1.3e-07 w=2.8e-07
mXI15_MXNOE ns cn XI15_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI15_MXNA1 XI15_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net076 nmse net070 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net070 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net074 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net076 D net074 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 pm c net076 VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN pm cn XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MX_t14 net80 m VDD VNW p12 l=1.3e-07 w=3.4e-07
MXP7 ns cn net80 VNW p12 l=1.3e-07 w=3.4e-07
mXI15_MXPOEN ns c XI15_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI15_MXPA1 XI15_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFQX2MTR Q VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net064 SE net055 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 VSS SI net064 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net059 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net055 D net059 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm cn net055 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE pm c XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net105 m VSS VPW n12 l=1.3e-07 w=3.9e-07
MX_t12 ns c net105 VPW n12 l=1.3e-07 w=3.9e-07
mXI15_MXNOE ns cn XI15_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI15_MXNA1 XI15_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net076 nmse net070 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net070 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net074 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net076 D net074 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 pm c net076 VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN pm cn XI16_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI16_MXPA1 XI16_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=4.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MX_t14 net80 m VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP8 ns cn net80 VNW p12 l=1.3e-07 w=4.9e-07
mXI15_MXPOEN ns c XI15_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI15_MXPA1 XI15_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQX4MTR Q VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net064 SE net055 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 VSS SI net064 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net059 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net055 D net059 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm cn net055 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE pm c XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net105 m VSS VPW n12 l=1.3e-07 w=4.4e-07
MX_t12 ns c net105 VPW n12 l=1.3e-07 w=4.4e-07
mXI15_MXNOE ns cn XI15_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI15_MXNA1 XI15_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net076 nmse net070 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net070 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net074 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net076 D net074 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 pm c net076 VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN pm cn XI16_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI16_MXPA1 XI16_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MX_t14 net80 m VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP9 ns cn net80 VNW p12 l=1.3e-07 w=6.4e-07
mXI15_MXPOEN ns c XI15_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI15_MXPA1 XI15_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRHQX1MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=3.5e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=3.5e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS RN net128 VPW n12 l=1.3e-07 w=4.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=4.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.7e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP8 net065 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=2.7e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP13 pm nmsi p1 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=6.6e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.3e-07
MX_t15 bm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 bm c net109 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=2.3e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFRHQX2MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS RN net128 VPW n12 l=1.3e-07 w=5.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=5.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP14 net065 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.9e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 pm nmsi p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
MX_t10_2 m pm VDD VNW p12 l=1.3e-07 w=5.1e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 bm RN VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP16 bm c net109 VNW p12 l=1.3e-07 w=1.5e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=1.5e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRHQX4MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS RN net128 VPW n12 l=1.3e-07 w=5.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=5.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP14 net065 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.9e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 pm nmsi p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
MX_t10_2 m pm VDD VNW p12 l=1.3e-07 w=5.1e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 bm RN VDD VNW p12 l=1.3e-07 w=3e-07
MXP16 bm c net109 VNW p12 l=1.3e-07 w=1.5e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=1.5e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRHQX8MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS RN net128 VPW n12 l=1.3e-07 w=5.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=5.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP14 net065 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.9e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 pm nmsi p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
MX_t10_2 m pm VDD VNW p12 l=1.3e-07 w=5.1e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 bm RN VDD VNW p12 l=1.3e-07 w=3e-07
MXP16 bm c net109 VNW p12 l=1.3e-07 w=1.5e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=1.5e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRQX1MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net130 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net130 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net138 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MX_t9 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN7 pm c net123 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net118 m net123 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net118 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE net76 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE net76 cn XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 s net76 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net97 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 nmrs SE net97 VNW p12 l=1.3e-07 w=3e-07
MXP1 nmrs nmse net105 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net105 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI74_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN net76 cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN net76 c XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s net76 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFRQX2MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net130 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net130 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net138 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MX_t9 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm c net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 net118 m net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN6 net118 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE net76 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE net76 cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1 s net76 XI1_n1 VPW n12 l=1.3e-07 w=2.7e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net97 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 nmrs SE net97 VNW p12 l=1.3e-07 w=3e-07
MXP1 nmrs nmse net105 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net105 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI74_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm cn net89 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD m net89 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN net76 cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN net76 c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s net76 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRQX4MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net130 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net130 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net138 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MX_t9 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm c net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 net118 m net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN6 net118 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE net76 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE net76 cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1 s net76 XI1_n1 VPW n12 l=1.3e-07 w=4.9e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net97 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 nmrs SE net97 VNW p12 l=1.3e-07 w=3e-07
MXP1 nmrs nmse net105 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net105 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI74_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm cn net89 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD m net89 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN net76 cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN net76 c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 s net76 VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRX1MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net104 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MXN9 nmrs nmse net104 VPW n12 l=1.3e-07 w=2.4e-07
MXN7 nmrs SE net77 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net77 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN12 pm c net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN13 net83 m net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net83 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNOE bm cn XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 s bm XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net139 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP10 nmrs SE net139 VNW p12 l=1.3e-07 w=3e-07
MXP8 nmrs nmse net115 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net115 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm cn net124 VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD m net124 VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPOEN bm c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFRX2MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net104 D net_clr_ VPW n12 l=1.3e-07 w=2.5e-07
MXN9 nmrs nmse net104 VPW n12 l=1.3e-07 w=2.5e-07
MXN7 nmrs SE net77 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net77 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.9e-07
MXN12 pm c net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN16 net83 m net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN17 net83 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.2e-07
mXI0_MXNOE bm cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1 s bm XI1_n1 VPW n12 l=1.3e-07 w=2.7e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net139 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP10 nmrs SE net139 VNW p12 l=1.3e-07 w=3e-07
MXP8 nmrs nmse net115 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net115 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP13 pm cn net124 VNW p12 l=1.3e-07 w=1.5e-07
MXP12 VDD m net124 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.4e-07
mXI0_MXPOEN bm c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRX4MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net104 D net_clr_ VPW n12 l=1.3e-07 w=4.9e-07
MXN9 nmrs nmse net104 VPW n12 l=1.3e-07 w=4.9e-07
MXN7 nmrs SE net77 VPW n12 l=1.3e-07 w=2.4e-07
MXN16 net77 SI net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MXN11 net_clr_ RN VSS VPW n12 l=1.3e-07 w=6.5e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=3.7e-07
MXN12 pm c net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN18 net83 m net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN19 net83 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=6.4e-07
mXI0_MXNOE bm cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1 s bm XI1_n1 VPW n12 l=1.3e-07 w=4.4e-07
mXI70_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI70_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net139 D VDD VNW p12 l=1.3e-07 w=6e-07
MXP14 nmrs SE net139 VNW p12 l=1.3e-07 w=6e-07
MXP13 nmrs nmse net115 VNW p12 l=1.3e-07 w=2.9e-07
MXP7 net115 SI VDD VNW p12 l=1.3e-07 w=2.9e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=3.9e-07
MXP15 pm cn net124 VNW p12 l=1.3e-07 w=1.5e-07
MXP12 VDD m net124 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.4e-07
mXI0_MXPOEN bm c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mXI70_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI70_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSHQX1MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net0112 SN VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN3 net169 cn net0112 VPW n12 l=1.3e-07 w=4.5e-07
MX_t11 pm nmsi net169 VPW n12 l=1.3e-07 w=4.5e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP3 net088 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=3e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm nmsi net56 VNW p12 l=1.3e-07 w=3.7e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT SDFFSHQX2MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.4e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net0104 SN VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN8 net169 cn net0104 VPW n12 l=1.3e-07 w=6.5e-07
MX_t11 pm nmsi net169 VPW n12 l=1.3e-07 w=6.5e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP8 net088 c cn VNW p12 l=1.3e-07 w=4.9e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=4.2e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=4.2e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=2.3e-07
MXP9 pm nmsi net56 VNW p12 l=1.3e-07 w=5.4e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.01e-06
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSHQX4MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net0104 SN VSS VPW n12 l=1.3e-07 w=7.4e-07
MXN10 net169 cn net0104 VPW n12 l=1.3e-07 w=7.4e-07
MX_t11 pm nmsi net169 VPW n12 l=1.3e-07 w=7.4e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.9e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP10 net088 c cn VNW p12 l=1.3e-07 w=5.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=3.8e-07
MXP11 pm nmsi net56 VNW p12 l=1.3e-07 w=6.9e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSHQX8MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net0104 SN VSS VPW n12 l=1.3e-07 w=7.5e-07
MXN12 net169 cn net0104 VPW n12 l=1.3e-07 w=7.5e-07
MXN13 pm nmsi net169 VPW n12 l=1.3e-07 w=7.5e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.9e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP10 net088 c cn VNW p12 l=1.3e-07 w=5.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=3.8e-07
MXP11 pm nmsi net56 VNW p12 l=1.3e-07 w=6.9e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSQX1MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmrs SE net150 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net150 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net123 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 nmrs nmse net123 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN11 bm cn net141 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 NSN s net141 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 nmrs SE net83 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net83 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 VDD SI net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net113 nmse nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 VDD pm m VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD SN m VNW p12 l=1.3e-07 w=2.3e-07
MXP13 VDD SN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP14 net107 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP15 net107 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSQX2MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmrs SE net150 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net150 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net123 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 nmrs nmse net123 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN11 bm cn net141 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 NSN s net141 VPW n12 l=1.3e-07 w=1.5e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 nmrs SE net83 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net83 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 VDD SI net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net113 nmse nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 VDD pm m VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD SN m VNW p12 l=1.3e-07 w=2.3e-07
MXP13 VDD SN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP16 net107 c bm VNW p12 l=1.3e-07 w=1.5e-07
MXP15 net107 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSQX4MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmrs SE net150 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net150 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net123 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 nmrs nmse net123 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN11 bm cn net141 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 NSN s net141 VPW n12 l=1.3e-07 w=1.5e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 nmrs SE net83 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net83 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 VDD SI net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net113 nmse nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 VDD pm m VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD SN m VNW p12 l=1.3e-07 w=2.3e-07
MXP13 VDD SN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP16 net107 c bm VNW p12 l=1.3e-07 w=1.5e-07
MXP15 net107 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRHQX1MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 net142 SN VSS VPW n12 l=1.3e-07 w=4.1e-07
MXN12 net166 cn net142 VPW n12 l=1.3e-07 w=4.1e-07
MX_t25 pm nmsi net166 VPW n12 l=1.3e-07 w=4.1e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=4.3e-07
MXN14 net170 RN VSS VPW n12 l=1.3e-07 w=4.3e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP12 net111 c cn VNW p12 l=1.3e-07 w=4.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmsi net131 VNW p12 l=1.3e-07 w=3.1e-07
MX_t28 net131 c VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 m RN net117 VNW p12 l=1.3e-07 w=2.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.6e-07
MXP21 bm nmset net93 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSRHQX2MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 net142 SN VSS VPW n12 l=1.3e-07 w=5.9e-07
MXN19 net166 cn net142 VPW n12 l=1.3e-07 w=5.9e-07
MXN20 pm nmsi net166 VPW n12 l=1.3e-07 w=5.9e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=6.1e-07
MXN21 net170 RN VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP12 net111 c cn VNW p12 l=1.3e-07 w=4.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmsi net131 VNW p12 l=1.3e-07 w=4.5e-07
MXP22 net131 c VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 m RN net117 VNW p12 l=1.3e-07 w=2.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP23 bm nmset net93 VNW p12 l=1.3e-07 w=2.7e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRHQX4MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN20 net142 SN VSS VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net166 cn net142 VPW n12 l=1.3e-07 w=7.5e-07
MX_t25 pm nmsi net166 VPW n12 l=1.3e-07 w=7.5e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=7.2e-07
MXN21 net170 RN VSS VPW n12 l=1.3e-07 w=7.2e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN22 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP22 net111 c cn VNW p12 l=1.3e-07 w=5.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.2e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.9e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP23 pm nmsi net131 VNW p12 l=1.3e-07 w=6.8e-07
MX_t28 net131 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP26 m RN net117 VNW p12 l=1.3e-07 w=3.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP27 bm nmset net93 VNW p12 l=1.3e-07 w=3.6e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRHQX8MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN20 net142 SN VSS VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net166 cn net142 VPW n12 l=1.3e-07 w=7.5e-07
MX_t25 pm nmsi net166 VPW n12 l=1.3e-07 w=7.5e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=7.2e-07
MXN21 net170 RN VSS VPW n12 l=1.3e-07 w=7.2e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN22 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP22 net111 c cn VNW p12 l=1.3e-07 w=5.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.2e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.9e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP23 pm nmsi net131 VNW p12 l=1.3e-07 w=6.8e-07
MX_t28 net131 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP26 m RN net117 VNW p12 l=1.3e-07 w=3.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP27 bm nmset net93 VNW p12 l=1.3e-07 w=3.6e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRX1MTR Q QN VDD VNW VPW VSS CK D RN SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE pm c XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MX_t15 NSN NRN m VPW n12 l=1.3e-07 w=1.9e-07
mXI60_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MXN5 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MX_t20 bm cn net75 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN s net75 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN pm cn XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 brn NRN VDD VNW p12 l=1.3e-07 w=4.9e-07
MX_t11 m pm brn VNW p12 l=1.3e-07 w=3.6e-07
MX_t12 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t16 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MXP6 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 brn s net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSRX2MTR Q QN VDD VNW VPW VSS CK D RN SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE pm c XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MX_t15 NSN NRN m VPW n12 l=1.3e-07 w=1.9e-07
mXI60_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MXN5 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MX_t20 bm cn net75 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN s net75 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN pm cn XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 brn NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP7 m pm brn VNW p12 l=1.3e-07 w=4.4e-07
MX_t12 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t16 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.4e-07
MXP6 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 brn s net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRX4MTR Q QN VDD VNW VPW VSS CK D RN SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=2.5e-07
mXI8_MXNOE pm c XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MX_t15 NSN NRN m VPW n12 l=1.3e-07 w=1.9e-07
mXI60_MXNOE bm c m VPW n12 l=1.3e-07 w=4.7e-07
MXN5 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MX_t20 bm cn net91 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN s net91 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=3e-07
mXI8_MXPOEN pm cn XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 brn NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP7 m pm brn VNW p12 l=1.3e-07 w=4.4e-07
MX_t12 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t16 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.7e-07
MXP6 bm c net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 brn s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSX1MTR Q QN VDD VNW VPW VSS CK D SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE pm c XI2_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNA1 XI2_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t11 m pm BSN VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MX_t19 bm cn net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 BSN s net138 VPW n12 l=1.3e-07 w=1.8e-07
MX_t33 BSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI33_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN pm cn XI2_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPA1 XI2_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MX_t24 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 bm c net104 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 VDD s net104 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI33_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSX2MTR Q QN VDD VNW VPW VSS CK D SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE pm c XI2_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNA1 XI2_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
MX_t11 m pm BSN VPW n12 l=1.3e-07 w=2.1e-07
MX_t11_2 m pm BSN VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MX_t19 bm cn net138 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN s net138 VPW n12 l=1.3e-07 w=1.5e-07
MX_t33 BSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN pm cn XI2_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPA1 XI2_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.4e-07
MX_t24 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm c net104 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD s net104 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI34_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSX4MTR Q QN VDD VNW VPW VSS CK D SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=2e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=2e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=2e-07
mXI2_MXNOE pm c XI2_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNA1 XI2_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.8e-07
MX_t11 m pm BSN VPW n12 l=1.3e-07 w=3.5e-07
MX_t11_2 m pm BSN VPW n12 l=1.3e-07 w=3.5e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.2e-07
MX_t19 bm cn net138 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN s net138 VPW n12 l=1.3e-07 w=1.5e-07
MX_t33 BSN SN VSS VPW n12 l=1.3e-07 w=1.08e-06
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI35_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI35_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=2.8e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=2.8e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.4e-07
mXI2_MXPOEN pm cn XI2_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPA1 XI2_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=7.8e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
MX_t24 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm c net104 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD s net104 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.9e-07
mXI35_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI35_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFTRX1MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net074 RN VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN5 net181 D net074 VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net181 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net193 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net193 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE bm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net96 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP7 nmrs SE net96 VNW p12 l=1.3e-07 w=3e-07
MXP6 nmrs nmse net114 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net114 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net105 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmrs RN net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI43_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI8_MXPOEN bm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFTRX2MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net074 RN VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN5 net181 D net074 VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net181 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net193 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net193 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mXI43_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI8_MXNOE bm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI47_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net96 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP7 nmrs SE net96 VNW p12 l=1.3e-07 w=3e-07
MXP6 nmrs nmse net114 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net114 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net105 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmrs RN net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI43_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI8_MXPOEN bm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFTRX4MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net074 RN VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN8 net181 D net074 VPW n12 l=1.3e-07 w=4.2e-07
MX_t7 nmrs nmse net181 VPW n12 l=1.3e-07 w=4.2e-07
MX_t3 nmrs SE net193 VPW n12 l=1.3e-07 w=2.3e-07
MXN7 net193 SI VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI43_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=3.4e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=8e-07
mXI8_MXNOE bm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI49_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI49_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net96 D VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP11 nmrs SE net96 VNW p12 l=1.3e-07 w=5.4e-07
MXP10 nmrs nmse net114 VNW p12 l=1.3e-07 w=2.7e-07
MX_t1 net114 SI VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP8 net105 SE VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP13 nmrs RN net105 VNW p12 l=1.3e-07 w=2.7e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI43_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=4.1e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_3 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_4 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI8_MXPOEN bm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=4.3e-07
mXI49_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI49_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFX1MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net137 SE net116 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net116 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net137 D net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 pm cn net137 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNOE pm c XI17_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 XI17_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI57_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI15_MXNOE sn c XI15_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI16_MXNOE sn cn XI16_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI16_MXNA1 XI16_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI58_MXNA1 Q sn VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 s sn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net77 nmse net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net73 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net76 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net77 D net76 VNW p12 l=1.3e-07 w=3.8e-07
MXP4 pm c net77 VNW p12 l=1.3e-07 w=3.8e-07
mXI17_MXPOEN pm cn XI17_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPA1 XI17_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI57_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI15_MXPOEN sn cn XI15_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI16_MXPOEN sn c XI16_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI16_MXPA1 XI16_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s sn VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPA1 Q sn VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFX2MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net137 SE net116 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net116 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net137 D net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 pm cn net137 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNOE pm c XI17_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 XI17_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI57_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI15_MXNOE sn c XI15_n1 VPW n12 l=1.3e-07 w=3.5e-07
mXI16_MXNOE sn cn XI16_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI16_MXNA1 XI16_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s sn VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI61_MXNA1 Q sn VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP5 net77 nmse net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net73 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net76 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net77 D net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm c net77 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPOEN pm cn XI17_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI17_MXPA1 XI17_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI57_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI15_MXPOEN sn cn XI15_p1 VNW p12 l=1.3e-07 w=4.9e-07
mXI16_MXPOEN sn c XI16_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI16_MXPA1 XI16_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s sn VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI61_MXPA1 Q sn VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT SDFFX4MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net137 SE net116 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net116 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net137 D net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 pm cn net137 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNOE pm c XI17_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 XI17_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI57_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=5.8e-07
mXI15_MXNOE sn c XI15_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI16_MXNOE sn cn XI16_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI16_MXNA1 XI16_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s sn VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI62_MXNA1 Q sn VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI62_MXNA1_2 Q sn VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP5 net77 nmse net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net73 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net76 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net77 D net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm c net77 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPOEN pm cn XI17_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI17_MXPA1 XI17_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=4.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI57_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI15_MXPOEN sn cn XI15_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI16_MXPOEN sn c XI16_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI16_MXPA1 XI16_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s sn VDD VNW p12 l=1.3e-07 w=4.2e-07
mXI62_MXPA1 Q sn VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI62_MXPA1_2 Q sn VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT SEDFFHQX1MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=2.3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=3.6e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.4e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=3e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP4 net079 c cn VNW p12 l=1.3e-07 w=4.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP5 pm nmsi net78 VNW p12 l=1.3e-07 w=4.4e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.4e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SEDFFHQX2MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=5.1e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=5.6e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=3.9e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP6 net079 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 pm nmsi net78 VNW p12 l=1.3e-07 w=6.2e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFHQX4MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=5.1e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=7e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.8e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 net079 c cn VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.8e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 pm nmsi net78 VNW p12 l=1.3e-07 w=6.2e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFHQX8MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=5.1e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=7e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.8e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 net079 c cn VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.8e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 pm nmsi net78 VNW p12 l=1.3e-07 w=6.2e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFTRX1MTR Q QN VDD VNW VPW VSS CK D E RN SE SI
MX_t9 nmrs RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmrs SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI44_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmsi SI VSS VPW n12 l=1.3e-07 w=1.7e-07
mXI38_MXNOE nmin_pass2 bse nmsi VPW n12 l=1.3e-07 w=1.8e-07
mXI39_MXNOE nmin_pass2 nmse nmin_pass1 VPW n12 l=1.3e-07 w=1.8e-07
mXI45_MXNA1 bse nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNOE nmin_pass1 be nmin VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE nmin_pass1 nmen s VPW n12 l=1.3e-07 w=1.8e-07
mX_g12_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 be nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net169 nmrs VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t5 net169 nmin_pass2 VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t4 pm cn net169 VPW n12 l=1.3e-07 w=2e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g18_MXNA1 nm m VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI59_MXNOE bnm c nm VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNOE bnm cn XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI46_MXNA1 QN bnm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP4 nmrs RN net108 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net108 SE VDD VNW p12 l=1.3e-07 w=3e-07
mXI44_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmsi SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI38_MXPOEN nmin_pass2 nmse nmsi VNW p12 l=1.3e-07 w=2.3e-07
mXI39_MXPOEN nmin_pass2 bse nmin_pass1 VNW p12 l=1.3e-07 w=2.3e-07
mXI45_MXPA1 bse nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPOEN nmin_pass1 nmen nmin VNW p12 l=1.3e-07 w=2.3e-07
mXI40_MXPOEN nmin_pass1 be s VNW p12 l=1.3e-07 w=2.3e-07
mX_g12_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 be nmen VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
MX_t1 net102 nmrs VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net111 nmin_pass2 net102 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 pm c net111 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g18_MXPA1 nm m VDD VNW p12 l=1.3e-07 w=4.1e-07
mXI59_MXPOEN bnm cn nm VNW p12 l=1.3e-07 w=4.1e-07
mXI1_MXPOEN bnm c XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI46_MXPA1 QN bnm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SEDFFTRX2MTR Q QN VDD VNW VPW VSS CK D E RN SE SI
MX_t9 nmrs RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmrs SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI44_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmsi SI VSS VPW n12 l=1.3e-07 w=1.7e-07
mXI38_MXNOE nmin_pass2 bse nmsi VPW n12 l=1.3e-07 w=1.8e-07
mXI39_MXNOE nmin_pass2 nmse nmin_pass1 VPW n12 l=1.3e-07 w=1.8e-07
mXI45_MXNA1 bse nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNOE nmin_pass1 be nmin VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE nmin_pass1 nmen s VPW n12 l=1.3e-07 w=1.8e-07
mX_g12_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 be nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN5 net169 nmrs VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t5 net169 nmin_pass2 VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t4 pm cn net169 VPW n12 l=1.3e-07 w=2e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g18_MXNA1 nm m VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE bnm c nm VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNOE bnm cn XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI47_MXNA1 QN bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmrs RN net108 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net108 SE VDD VNW p12 l=1.3e-07 w=3e-07
mXI44_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmsi SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI38_MXPOEN nmin_pass2 nmse nmsi VNW p12 l=1.3e-07 w=2.3e-07
mXI39_MXPOEN nmin_pass2 bse nmin_pass1 VNW p12 l=1.3e-07 w=2.3e-07
mXI45_MXPA1 bse nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPOEN nmin_pass1 nmen nmin VNW p12 l=1.3e-07 w=2.3e-07
mXI40_MXPOEN nmin_pass1 be s VNW p12 l=1.3e-07 w=2.3e-07
mX_g12_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 be nmen VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t1 net102 nmrs VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net111 nmin_pass2 net102 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 pm c net111 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g18_MXPA1 nm m VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI59_MXPOEN bnm cn nm VNW p12 l=1.3e-07 w=5.9e-07
mXI1_MXPOEN bnm c XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI47_MXPA1 QN bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFTRX4MTR Q QN VDD VNW VPW VSS CK D E RN SE SI
MX_t9 nmrs RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmrs SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI44_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmsi SI VSS VPW n12 l=1.3e-07 w=1.7e-07
mXI38_MXNOE nmin_pass2 bse nmsi VPW n12 l=1.3e-07 w=1.8e-07
mXI39_MXNOE nmin_pass2 nmse nmin_pass1 VPW n12 l=1.3e-07 w=1.8e-07
mXI45_MXNA1 bse nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNOE nmin_pass1 be nmin VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE nmin_pass1 nmen s VPW n12 l=1.3e-07 w=1.8e-07
mX_g12_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 be nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN5 net169 nmrs VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t5 net169 nmin_pass2 VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t4 pm cn net169 VPW n12 l=1.3e-07 w=2e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g18_MXNA1 nm m VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE bnm c nm VPW n12 l=1.3e-07 w=7.4e-07
mXI1_MXNOE bnm cn XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI48_MXNA1 QN bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI48_MXNA1_2 QN bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmrs RN net108 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net108 SE VDD VNW p12 l=1.3e-07 w=3e-07
mXI44_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmsi SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI38_MXPOEN nmin_pass2 nmse nmsi VNW p12 l=1.3e-07 w=2.3e-07
mXI39_MXPOEN nmin_pass2 bse nmin_pass1 VNW p12 l=1.3e-07 w=2.3e-07
mXI45_MXPA1 bse nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPOEN nmin_pass1 nmen nmin VNW p12 l=1.3e-07 w=2.3e-07
mXI40_MXPOEN nmin_pass1 be s VNW p12 l=1.3e-07 w=2.3e-07
mX_g12_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 be nmen VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t1 net102 nmrs VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net111 nmin_pass2 net102 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 pm c net111 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.9e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g18_MXPA1 nm m VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI59_MXPOEN bnm cn nm VNW p12 l=1.3e-07 w=8e-07
mXI1_MXPOEN bnm c XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI48_MXPA1 QN bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI48_MXPA1_2 QN bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFX1MTR Q QN VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net180 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net187 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net190 SE net187 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net190 D net181 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net181 E net180 VPW n12 l=1.3e-07 w=1.8e-07
MX_t16 net196 nmen net180 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net196 s net190 VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 pm cn net190 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI3_MXNOE nm c XI3_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI4_MXNOE nm cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI41_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t6 net85 SE VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t8 net97 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net96 nmse net97 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net96 D net91 VNW p12 l=1.3e-07 w=4.7e-07
MX_t5 net91 nmen net85 VNW p12 l=1.3e-07 w=4.7e-07
MXP9 net88 E net85 VNW p12 l=1.3e-07 w=4.7e-07
MXP10 net88 s net96 VNW p12 l=1.3e-07 w=4.7e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm c net96 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI40_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI3_MXPOEN nm cn XI3_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI4_MXPOEN nm c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.4e-07
mXI41_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SEDFFX2MTR Q QN VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net100 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net92 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net88 SE net92 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net88 D net76 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net76 E net100 VPW n12 l=1.3e-07 w=1.8e-07
MX_t16 net84 nmen net100 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net84 s net88 VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 pm cn net88 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI3_MXNOE nm c XI3_n1 VPW n12 l=1.3e-07 w=4.4e-07
mXI4_MXNOE nm cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI42_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t6 net127 SE VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t8 net111 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net113 nmse net111 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net113 D net131 VNW p12 l=1.3e-07 w=4.7e-07
MX_t5 net131 nmen net127 VNW p12 l=1.3e-07 w=4.7e-07
MXP9 net105 E net127 VNW p12 l=1.3e-07 w=4.7e-07
MXP10 net105 s net113 VNW p12 l=1.3e-07 w=4.7e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm c net113 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI40_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI3_MXPOEN nm cn XI3_p1 VNW p12 l=1.3e-07 w=5.4e-07
mXI4_MXPOEN nm c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI42_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFX4MTR Q QN VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net100 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net92 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net88 SE net92 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net88 D net76 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net76 E net100 VPW n12 l=1.3e-07 w=1.8e-07
MX_t16 net84 nmen net100 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net84 s net88 VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 pm cn net88 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI40_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI3_MXNOE nm c XI3_n1 VPW n12 l=1.3e-07 w=6.4e-07
mXI4_MXNOE nm cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI43_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI43_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 net127 SE VDD VNW p12 l=1.3e-07 w=2.4e-07
MXP14_2 net127 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net111 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net113 nmse net111 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net113 D net131 VNW p12 l=1.3e-07 w=4.7e-07
MX_t5 net131 nmen net127 VNW p12 l=1.3e-07 w=4.7e-07
MXP12 net105 E net127 VNW p12 l=1.3e-07 w=4.6e-07
MXP13 net105 s net113 VNW p12 l=1.3e-07 w=4.6e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm c net113 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI40_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI3_MXPOEN nm cn XI3_p1 VNW p12 l=1.3e-07 w=7.3e-07
mXI4_MXPOEN nm c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI43_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI43_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SMDFFHQX1MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=1.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=2.1e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN4 VSS cn net107 VPW n12 l=1.3e-07 w=3.3e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=3.3e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=3.7e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=2.6e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=2.6e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=3e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=3e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=4.2e-07
MXP0 cn c net085 VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=4e-07
MXP3 pm nmsi net060 VNW p12 l=1.3e-07 w=4e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=7.3e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SMDFFHQX2MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=1.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=3.1e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=3e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN5 VSS cn net107 VPW n12 l=1.3e-07 w=4.8e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=4.8e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=4.4e-07
MXP4 cn c net085 VNW p12 l=1.3e-07 w=4.4e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP5 pm nmsi net060 VNW p12 l=1.3e-07 w=5.9e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=9.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=9.8e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SMDFFHQX4MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=2.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=5e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN6 VSS cn net107 VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=5.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=3.4e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net085 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net060 VNW p12 l=1.3e-07 w=1.01e-06
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SMDFFHQX8MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=2.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=5e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN6 VSS cn net107 VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=5.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=3.4e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net085 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net060 VNW p12 l=1.3e-07 w=1.01e-06
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends

