* ---------------------------------------------------------------------------- 
* 
*     library Calibre-based CDL file 
* 
*     Date: Jan 31, 2012 7:10:22 PM IST 
* 
*     CellBuilder version 4.0.1 -- built on Nov 11, 2011 
*     Copyright (c) 2002-2011 ARM, Inc. 
*     The confidential and proprietary information contained in this file 
*     may only be used by a person authorised under and to the extent 
*     permitted by a subsisting licensing agreement from ARM Limited. 
*      
*     (C) COPYRIGHT 2004-2012 ARM Limited. 
*     ALL RIGHTS RESERVED 
*      
*     This entire notice must be reproduced on all copies of this file 
*     and copies of this file may only be made by a person if such person 
*     is permitted to do so under the terms of a subsisting license 
*     agreement from ARM Limited. 
* 
* ----------------------------------------------------------------------------

*.SCALE METER
*.OPTION SCALE 1e-6

.SUBCKT ADDFHX1MTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=130n w=530n
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=270n
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=6.3e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.9e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=6.3e-07
mXI5_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=3.9e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI11_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=3.7e-07
mXI12_MXNOE con xorab cin VPW n12 l=1.3e-07 w=3.7e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=3.7e-07
mXI10_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=3.7e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=7.7e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=7.7e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=7.7e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=5.8e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=7.7e-07
mXI5_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=6.8e-07
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI11_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=4.6e-07
mXI12_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=4.6e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=4.6e-07
mXI10_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=4.6e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT ADDFHX2MTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI15_MXNA1_2 ba na2 VSS VPW n12 l=1.3e-07 w=6e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=5.2e-07
mXI3_MXNOE_2 xnorab B ba VPW n12 l=1.3e-07 w=5.2e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNOE_2 xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=3.9e-07
mXI4_MXNOE_2 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI4_MXNOE_3 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI5_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=9.3e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI6_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI11_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=6.1e-07
mXI12_MXNOE con xorab cin VPW n12 l=1.3e-07 w=5.4e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI9_MXNOE_2 sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI10_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=5.5e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI7_MXNA1_2 cin CI VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI14_MXNA1_2 CO con VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI15_MXPA1_2 ba na2 VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=6.3e-07
mXI3_MXPOEN_2 xnorab nb ba VNW p12 l=1.3e-07 w=6.3e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPOEN_2 xnorab B na VNW p12 l=1.3e-07 w=5e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=6.3e-07
mXI4_MXPOEN_2 xorab nb na VNW p12 l=1.3e-07 w=6.3e-07
mXI5_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=1.22e-06
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI11_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=3.7e-07
mXI11_MXPOEN_2 con xorab nb VNW p12 l=1.3e-07 w=4.4e-07
mXI12_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=6e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=7.4e-07
mXI10_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=7.4e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=9.8e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI13_MXPA1_2 S sumn VDD VNW p12 l=1.3e-07 w=4.4e-07
.ends


.SUBCKT ADDFHX4MTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=8.6e-07
mXI15_MXNA1_2 ba na2 VSS VPW n12 l=1.3e-07 w=8.6e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=8.6e-07
mXI3_MXNOE_2 xnorab B ba VPW n12 l=1.3e-07 w=6.7e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNOE_2 xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=3.9e-07
mXI4_MXNOE_2 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI4_MXNOE_3 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI5_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=9.3e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=9.8e-07
mXI6_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=9.8e-07
mXI6_MXNA1_3 nb B VSS VPW n12 l=1.3e-07 w=9.8e-07
mXI11_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=6.1e-07
mXI12_MXNOE con xorab cin VPW n12 l=1.3e-07 w=5.4e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI9_MXNOE_2 sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI10_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=5.5e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI8_MXNA1_2 cib cin VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1_2 cin CI VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1_3 cin CI VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI14_MXNA1_2 CO con VSS VPW n12 l=1.3e-07 w=7e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI13_MXNA1_2 S sumn VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI15_MXPA1_2 ba na2 VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI15_MXPA1_3 ba na2 VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=6.7e-07
mXI3_MXPOEN_2 xnorab nb ba VNW p12 l=1.3e-07 w=6.7e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=5.5e-07
mXI1_MXPOEN_2 xnorab B na VNW p12 l=1.3e-07 w=5.5e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=8.6e-07
mXI4_MXPOEN_2 xorab nb na VNW p12 l=1.3e-07 w=1.01e-06
mXI5_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=1.2e-06
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_5 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_6 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_7 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI11_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=5.2e-07
mXI11_MXPOEN_2 con xorab nb VNW p12 l=1.3e-07 w=5.2e-07
mXI12_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=6e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=7.4e-07
mXI10_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=9.8e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=9.8e-07
mXI8_MXPA1_2 cib cin VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=9.8e-07
mXI7_MXPA1_2 cin CI VDD VNW p12 l=1.3e-07 w=9.8e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI14_MXPA1_2 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1_2 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT ADDFHX8MTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_4 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_5 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI2_MXNA1_2 na2 A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI2_MXNA1_3 na2 A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_2 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_3 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_4 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_5 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_6 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=6.9e-07
mXI3_MXNOE_2 xnorab B ba VPW n12 l=1.3e-07 w=6.7e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNOE_2 xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=3.7e-07
mXI4_MXNOE_2 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI4_MXNOE_3 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI5_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=6.7e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=9.9e-07
mXI6_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=9.9e-07
mXI11_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=6.1e-07
mXI12_MXNOE con xorab cin VPW n12 l=1.3e-07 w=5.4e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI9_MXNOE_2 sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI10_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=5.5e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI7_MXNA1_2 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI7_MXNA1_3 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI7_MXNA1_4 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI7_MXNA1_5 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI14_MXNA1_2 CO con VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI14_MXNA1_3 CO con VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI14_MXNA1_4 CO con VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNA1_2 S sumn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNA1_3 S sumn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNA1_4 S sumn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_4 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_5 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_6 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI2_MXPA1_2 na2 A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI2_MXPA1_3 na2 A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_2 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_3 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_4 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_5 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_6 ba na2 VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=6.7e-07
mXI3_MXPOEN_2 xnorab nb ba VNW p12 l=1.3e-07 w=6.7e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=5.5e-07
mXI1_MXPOEN_2 xnorab B na VNW p12 l=1.3e-07 w=5.5e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=8.6e-07
mXI4_MXPOEN_2 xorab nb na VNW p12 l=1.3e-07 w=1.01e-06
mXI5_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=1.22e-06
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI11_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=5.3e-07
mXI11_MXPOEN_2 con xorab nb VNW p12 l=1.3e-07 w=5.3e-07
mXI12_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=6e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=9.8e-07
mXI10_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=9.8e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI7_MXPA1_2 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI7_MXPA1_3 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI7_MXPA1_4 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI7_MXPA1_5 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI14_MXPA1_2 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI14_MXPA1_3 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI14_MXPA1_4 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI13_MXPA1_2 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1_3 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1_4 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT ADDFHXLMTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=3.5e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.5e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=3.5e-07
mXI25_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=3.5e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI23_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=2.1e-07
mXI24_MXNOE con xorab cin VPW n12 l=1.3e-07 w=2.1e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=2.1e-07
mXI22_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=2.1e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=4.3e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=4.3e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=4.3e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=4.3e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=4.3e-07
mXI25_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=4.3e-07
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI23_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=2.5e-07
mXI24_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=2.5e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=2.5e-07
mXI22_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=2.5e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT ADDFX1MTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT ADDFX2MTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.5e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.8e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDFX4MTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.5e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDFX8MTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 CO nco VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_3 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.5e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDFXLMTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT ADDHX1MTR CO S VDD VNW VPW VSS A B
mX_g3_MXNA1 ba na VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNOE S nb ba VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE S B na VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 na A VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g2_MXNA2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g2_MXNA1 nco B X_g2_n1 VPW n12 l=1.3e-07 w=2.3e-07
mX_g0_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 ba na VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPOEN S B ba VNW p12 l=1.3e-07 w=3.8e-07
mXI9_MXPOEN S nb na VNW p12 l=1.3e-07 w=3.8e-07
mX_g4_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g2_MXPA2 nco A VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 nco B VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT ADDHX2MTR CO S VDD VNW VPW VSS A B
mX_g1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g3_MXNA1 ba na VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI10_MXNOE S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE S B na VPW n12 l=1.3e-07 w=6e-07
mX_g2_MXNA1 nco B X_g2_n1 VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g4_MXNA1 na A VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g4_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g4_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=5.9e-07
mX_g0_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g3_MXPA1 ba na VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI10_MXPOEN S B ba VNW p12 l=1.3e-07 w=7.5e-07
mXI9_MXPOEN S nb na VNW p12 l=1.3e-07 w=7.5e-07
mX_g2_MXPA1 nco B VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA2 nco A VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g4_MXPA1 na A VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDHX4MTR CO S VDD VNW VPW VSS A B
mX_g3_MXNA1 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI10_MXNOE S nb ba VPW n12 l=1.3e-07 w=5.9e-07
mXI10_MXNOE_2 S nb ba VPW n12 l=1.3e-07 w=5.9e-07
mXI9_MXNOE S B na VPW n12 l=1.3e-07 w=5.9e-07
mXI9_MXNOE_2 S B na VPW n12 l=1.3e-07 w=5.9e-07
mX_g2_MXNA1 nco B X_g2_n1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1_4 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1_5 na A VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g0_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI10_MXPOEN S B ba VNW p12 l=1.3e-07 w=7.6e-07
mXI10_MXPOEN_2 S B ba VNW p12 l=1.3e-07 w=7.6e-07
mXI9_MXPOEN S nb na VNW p12 l=1.3e-07 w=7.6e-07
mXI9_MXPOEN_2 S nb na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 nco B VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g2_MXPA2 nco A VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g4_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g4_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g4_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g4_MXPA1_4 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g4_MXPA1_5 na A VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g0_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDHX8MTR CO S VDD VNW VPW VSS A B
mX_g3_MXNA1 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_3 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_4 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=5.7e-07
mX_g1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI10_MXNOE S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI10_MXNOE_2 S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI10_MXNOE_3 S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI10_MXNOE_4 S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE S B na VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE_2 S B na VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE_3 S B na VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE_4 S B na VPW n12 l=1.3e-07 w=6e-07
mX_g2_MXNA1 nco B X_g2_n1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nco B X_g2_n1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA2_2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g4_MXNA1_4 na A VSS VPW n12 l=1.3e-07 w=7e-07
mX_g4_MXNA1_5 na A VSS VPW n12 l=1.3e-07 w=7e-07
mX_g4_MXNA1_6 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_7 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_8 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_9 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_10 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI10_MXPOEN S B ba VNW p12 l=1.3e-07 w=6.1e-07
mXI10_MXPOEN_2 S B ba VNW p12 l=1.3e-07 w=6.1e-07
mXI10_MXPOEN_3 S B ba VNW p12 l=1.3e-07 w=6.1e-07
mXI10_MXPOEN_4 S B ba VNW p12 l=1.3e-07 w=6.1e-07
mXI9_MXPOEN S nb na VNW p12 l=1.3e-07 w=5.8e-07
mXI9_MXPOEN_2 S nb na VNW p12 l=1.3e-07 w=8.2e-07
mXI9_MXPOEN_3 S nb na VNW p12 l=1.3e-07 w=8.2e-07
mXI9_MXPOEN_4 S nb na VNW p12 l=1.3e-07 w=8.2e-07
mX_g2_MXPA1 nco B VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g2_MXPA1_2 nco B VDD VNW p12 l=1.3e-07 w=7.5e-07
mX_g2_MXPA2 nco A VDD VNW p12 l=1.3e-07 w=7.5e-07
mX_g2_MXPA2_2 nco A VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g4_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_4 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_5 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_6 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_7 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_8 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_9 na A VDD VNW p12 l=1.3e-07 w=8.6e-07
mX_g4_MXPA1_10 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND2X12MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA2_2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA2_3 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1_2 ny A XI0_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1_3 ny A XI0_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=6e-07
.ends


.SUBCKT AND2X1MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.1e-07
.ends


.SUBCKT AND2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND3X12MTR Y VDD VNW VPW VSS A B C
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A XI0_n2__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n2__3 B XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n1__3 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA3_3 ny C VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=5.9e-07
.ends


.SUBCKT AND3X1MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AND3X2MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND3X4MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND3X6MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_2 ny A XI0_n2__2 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND3X8MTR Y VDD VNW VPW VSS A B C
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 ny A XI0_n2__2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 ny A XI0_n2__3 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_3 XI0_n2__3 B XI0_n1__3 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3_3 XI0_n1__3 C VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3_3 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
.ends


.SUBCKT AND3XLMTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AND4X12MTR Y VDD VNW VPW VSS A B C D
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 ny A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA4_2 ny D VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA4_3 ny D VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA4_4 ny D VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA3_3 ny C VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA3_4 ny C VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA2_4 ny B VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=5e-07
.ends


.SUBCKT AND4X1MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=3.3e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=3.3e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=3.3e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AND4X2MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND4X4MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4_2 XI0_n1__2 D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3_2 XI0_n2__2 C XI0_n1__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_2 XI0_n3__2 B XI0_n2__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 ny A XI0_n3__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA4_2 ny D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND4X6MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA1_2 ny A XI0_n3 VPW n12 l=1.3e-07 w=6.5e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA4_2 ny D VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND4X8MTR Y VDD VNW VPW VSS A B C D
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 ny A XI0_n3 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 ny A XI0_n3 VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA4_2 ny D VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA4_3 ny D VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3_3 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
.ends


.SUBCKT AND4XLMTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends




.SUBCKT AO21X1MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AO21X2MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO21X4MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO21X8MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 ny A0 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 ny B0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO21XLMTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.4e-07
.ends


.SUBCKT AO22X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.1e-07
.ends


.SUBCKT AO22X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=4.4e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=4.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO22X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO22X8MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2_2 XI0_n1B__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 ny B0 XI0_n1B__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1A__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A0 XI0_n1A__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO22XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AO2B2BX1MTR Y VDD VNW VPW VSS A0 A1N B0 B1N
mXI2_MXNA1 b1 B1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN6 net34 b1 VSS VPW n12 l=1.3e-07 w=2.3e-07
MXNB0 ny B0 net34 VPW n12 l=1.3e-07 w=2.3e-07
MXN4 ny A0 net40 VPW n12 l=1.3e-07 w=2.3e-07
MXN5 net40 a1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI2_MXPA1 b1 B1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net46 b1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXPB0 net46 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 ny A0 net46 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 ny a1 net46 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AO2B2BX2MTR Y VDD VNW VPW VSS A0 A1N B0 B1N
mXI2_MXNA1 b1 B1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN9 net34 b1 VSS VPW n12 l=1.3e-07 w=3.7e-07
MXNB0 ny B0 net34 VPW n12 l=1.3e-07 w=3.7e-07
MXN7 ny A0 net40 VPW n12 l=1.3e-07 w=3.7e-07
MXN8 net40 a1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 b1 B1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net46 b1 VDD VNW p12 l=1.3e-07 w=4.4e-07
MXPB0 net46 B0 VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP7 ny A0 net46 VNW p12 l=1.3e-07 w=4.4e-07
MXP9 ny a1 net46 VNW p12 l=1.3e-07 w=4.4e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO2B2BX4MTR Y VDD VNW VPW VSS A0 A1N B0 B1N
mXI2_MXNA1 b1 B1N VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN12 net34 b1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 ny B0 net34 VPW n12 l=1.3e-07 w=7.1e-07
MXN10 ny A0 net40 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 net40 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 b1 B1N VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP10 net46 b1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPB0 net46 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12 ny A0 net46 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 ny a1 net46 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO2B2BXLMTR Y VDD VNW VPW VSS A0 A1N B0 B1N
mXI2_MXNA1 b1 B1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN15 net34 b1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNB0 ny B0 net34 VPW n12 l=1.3e-07 w=1.8e-07
MXN13 ny A0 net40 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net40 a1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXPA1 b1 B1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 net46 b1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 net46 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 ny A0 net46 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 ny a1 net46 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AO2B2X1MTR Y VDD VNW VPW VSS A0 A1N B0 B1
MXN8 net051 B1 VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN5 ny B0 net051 VPW n12 l=1.3e-07 w=2.3e-07
MXN6 ny A0 net35 VPW n12 l=1.3e-07 w=2.3e-07
MXN7 net35 a1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP5 net41 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net41 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 ny A0 net41 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 ny a1 net41 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AO2B2X2MTR Y VDD VNW VPW VSS A0 A1N B0 B1
MXN12 net051 B1 VSS VPW n12 l=1.3e-07 w=3.7e-07
MXN13 ny B0 net051 VPW n12 l=1.3e-07 w=3.7e-07
MXN10 ny A0 net35 VPW n12 l=1.3e-07 w=3.7e-07
MXN11 net35 a1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP9 net41 B1 VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP10 net41 B0 VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP11 ny A0 net41 VNW p12 l=1.3e-07 w=4.4e-07
MXP12 ny a1 net41 VNW p12 l=1.3e-07 w=4.4e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO2B2X4MTR Y VDD VNW VPW VSS A0 A1N B0 B1
MXN2 net051 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 ny B0 net051 VPW n12 l=1.3e-07 w=7.1e-07
MXN0 ny A0 net35 VPW n12 l=1.3e-07 w=7.1e-07
MXN1 net35 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP14 net41 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 net41 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16 ny A0 net41 VNW p12 l=1.3e-07 w=8.7e-07
MXP17 ny a1 net41 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO2B2XLMTR Y VDD VNW VPW VSS A0 A1N B0 B1
MXN7 net051 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 ny B0 net051 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 ny A0 net35 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net35 a1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP19 net41 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP20 net41 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP21 ny A0 net41 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 ny a1 net41 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI211X1MTR Y VDD VNW VPW VSS A0 A1 B0 C0
MXN5 Y A0 net17 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 net17 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN4 Y C0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNC0 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP6 p1 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXPA1 p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 net045 C0 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 Y B0 net045 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI211X2MTR Y VDD VNW VPW VSS A0 A1 B0 C0
MXN8 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y C0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNC0 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP9 p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA1 p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net045 C0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 Y B0 net045 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI211X4MTR Y VDD VNW VPW VSS A0 A1 B0 C0
MXN12_2 net17__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y A0 net17__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 Y C0 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN13 Y B0 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN13_2 Y B0 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN10_2 Y C0 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXPA1 p1 A1 VDD VNW p12 l=1.3e-07 w=8e-07
MXP12 p1 A0 VDD VNW p12 l=1.3e-07 w=8e-07
MXP12_2 p1 A0 VDD VNW p12 l=1.3e-07 w=8e-07
MXPA1_2 p1 A1 VDD VNW p12 l=1.3e-07 w=8e-07
MXP13_2 net045__2 C0 p1 VNW p12 l=1.3e-07 w=8e-07
MXP14_2 Y B0 net045__2 VNW p12 l=1.3e-07 w=8e-07
MXP14 Y B0 net045 VNW p12 l=1.3e-07 w=8e-07
MXP13 net045 C0 p1 VNW p12 l=1.3e-07 w=8e-07
.ends


.SUBCKT AOI211XLMTR Y VDD VNW VPW VSS A0 A1 B0 C0
MXN8 Y A0 net17 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net17 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 Y C0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNC0 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP9 p1 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXPA1 p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP10 net045 C0 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP11 Y B0 net045 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI21BX1MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=3e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI21BX2MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21BX4MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=3.4e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI2_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21BX8MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI1_MXNA2_2 XI1_n1__2 B0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 ny a0a1 XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1_2 ny a0a1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2_2 ny B0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI2_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI2_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI2_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21BXLMTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=3e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI21X1MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI21X2MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21X3MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB1_2 Y A0 XI0_n1__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT AOI21X4MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 Y A0 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21X6MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB1_2 Y A0 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_3 XI0_n1__3 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 Y A0 XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_3 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_3 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21X8MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 Y A0 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 Y A0 XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_3 XI0_n1__3 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_4 XI0_n1__4 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_4 Y A0 XI0_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_3 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_3 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_4 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_4 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21XLMTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI221X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN7 Y B0 net26 VPW n12 l=1.3e-07 w=3.6e-07
MXN10 net26 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN9 net17 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN8 Y A0 net17 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y C0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP5 p1 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP6 p1 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 p2 A1 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP9 p2 A0 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 Y C0 p2 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI221X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN14 net26 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B0 net26 VPW n12 l=1.3e-07 w=7.1e-07
MXN12 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXN13 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP10 p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5 p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12 p2 A0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 p2 A1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 Y C0 p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI221X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN18_2 net26__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 Y B0 net26__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN15 Y B0 net26 VPW n12 l=1.3e-07 w=7.1e-07
MXN18 net26 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN17_2 net17__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN16_2 Y A0 net17__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN16 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXN17 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y C0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP14 p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5 p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP14_2 p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 p2 A1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP16 p2 A0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 p2 A0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP15_2 p2 A1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP17 Y C0 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 Y C0 p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI221XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN12 Y B0 net26 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net26 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net17 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 Y A0 net17 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 Y C0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP10 p1 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP11 p1 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP12 p2 A1 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP13 p2 A0 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP14 Y C0 p2 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI222X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN6 Y C0 net29 VPW n12 l=1.3e-07 w=3.6e-07
MXN4 net29 C1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net26 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y B0 net26 VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y A0 net17 VPW n12 l=1.3e-07 w=3.6e-07
MXN2 net17 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP5 p1 C0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP6 p1 C1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 p2 B1 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 p2 B0 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP9 Y A0 p2 VNW p12 l=1.3e-07 w=6.2e-07
MXP10 Y A1 p2 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI222X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN10 net29 C1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 Y C0 net29 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y B0 net26 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net26 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXP11 p1 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12 p1 C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP13 p2 B0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 p2 B1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP15 Y A1 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP16 Y A0 p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI222X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN11_2 Y C0 net29__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN16_2 net29__2 C1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN16 net29 C1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y C0 net29 VPW n12 l=1.3e-07 w=7.1e-07
MXN12_2 Y B0 net26__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 net26__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15 net26 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 Y B0 net26 VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 Y A0 net17__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 net17__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXP5 p1 C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17 p1 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 p1 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 p1 C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP18 p2 B0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP19 p2 B1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_2 p2 B1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 p2 B0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP21 Y A0 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP20 Y A1 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 Y A1 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP21_2 Y A0 p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI222XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN11 Y C0 net29 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net29 C1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net26 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 Y B0 net26 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 Y A0 net17 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net17 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP12 p1 C0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP11 p1 C1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP14 p2 B1 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP13 p2 B0 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP16 Y A0 p2 VNW p12 l=1.3e-07 w=3.6e-07
MXP15 Y A1 p2 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI22X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 Y B0 XI0_n1B VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A0 XI0_n1A VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI22X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y B0 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI22X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB1_2 Y B0 XI0_n1B__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1B__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y B0 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A0 XI0_n1A__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1A__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI22XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 Y B0 XI0_n1B VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A0 XI0_n1A VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI2B1X1MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN3 net022 a1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=3.6e-07
MXN4 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net36 a1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP5 Y B0 net36 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI2B1X2MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=3e-07
MXN5 net022 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP8 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2B1X4MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN7_2 net022__2 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_2 Y A0 net022__2 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=7.1e-07
MXN7 net022 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP8 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0_2 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
MXP9_2 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2B1X8MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 net022__2 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_2 Y A0 net022__2 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_3 Y A0 net022__3 VPW n12 l=1.3e-07 w=7.1e-07
MXN9_3 net022__3 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_4 net022__4 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_4 Y A0 net022__4 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net022 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10_3 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10_4 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0_2 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10_2 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10_3 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0_3 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0_4 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10_4 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP11 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
MXP11_2 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
MXP11_3 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
MXP11_4 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2B1XLMTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN5 net022 a1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net36 a1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP7 Y B0 net36 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI2BB1X1MTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI2BB1X2MTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB1X4MTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA2_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2_2 XI24_p1__2 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_2 Y nmin XI24_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB1X8MTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNA1_2 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNA2_2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA2_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA2_3 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA2_4 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI23_MXPA2_2 XI23_p1__2 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI23_MXPA1_2 nmin A0N XI23_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2_2 XI24_p1__2 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_2 Y nmin XI24_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_3 Y nmin XI24_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2_3 XI24_p1__3 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2_4 XI24_p1__4 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_4 Y nmin XI24_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB1XLMTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=3e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=3e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI2BB2X1MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI2BB2X2MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB2X4MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2_2 XI27_n1__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1_2 Y B0 XI27_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1_2 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1_2 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2_2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB2X8MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI28_MXNA2_2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI28_MXNA1_2 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2_2 XI27_n1__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1_2 Y B0 XI27_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1_3 Y B0 XI27_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2_3 XI27_n1__3 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2_4 XI27_n1__4 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1_4 Y B0 XI27_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI28_MXPA1_2 nmin A0N XI28_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI28_MXPA2_2 XI28_p1__2 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1_2 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1_3 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1_4 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1_2 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2_2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2_3 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1_3 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1_4 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2_4 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB2XLMTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=3e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=3e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI31X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0
mXI0_MXNB3 XI0_n1 A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB2 XI0_n2 A1 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 Y A0 XI0_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI31X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0
mXI0_MXNB3 XI0_n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n2 A1 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI31X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0
mXI0_MXNB1_2 Y A0 XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n2__2 A1 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB3_2 XI0_n1__2 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB3 XI0_n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n2 A1 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB3_2 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI31XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0
mXI0_MXNB3 XI0_n1 A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB2 XI0_n2 A1 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 Y A0 XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI32X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
mXI0_MXNB3 XI0_n1B A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB2 XI0_n2B A1 XI0_n1B VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 Y A0 XI0_n2B VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 XI0_n1A VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 XI0_n1A B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI32X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
mXI0_MXNB3 XI0_n1B A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n2B A1 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n2B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI32X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
mXI0_MXNB1_2 Y A0 XI0_n2B__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n2B__2 A1 XI0_n1B__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB3_2 XI0_n1B__2 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB3 XI0_n1B A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n2B A1 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n2B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n1A__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1A__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB3_2 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI32XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
mXI0_MXNB3 XI0_n1B A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB2 XI0_n2B A1 XI0_n1B VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 Y A0 XI0_n2B VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 XI0_n1A VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1A B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI33X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN8 net55 B2 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN7 net49 B1 net55 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y B0 net49 VPW n12 l=1.3e-07 w=3.6e-07
MXNA0 Y A0 net43 VPW n12 l=1.3e-07 w=3.6e-07
MXN9 net43 A1 net40 VPW n12 l=1.3e-07 w=3.6e-07
MXN10 net40 A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP12 net057 B2 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 net057 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXPB0 net057 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 Y A0 net057 VNW p12 l=1.3e-07 w=6.2e-07
MXP14 Y A1 net057 VNW p12 l=1.3e-07 w=6.2e-07
MXP13 Y A2 net057 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI33X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN13 net55 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net49 B1 net55 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B0 net49 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net43 VPW n12 l=1.3e-07 w=7.1e-07
MXN15 net43 A1 net40 VPW n12 l=1.3e-07 w=7.1e-07
MXN14 net40 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP12 net057 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP11 net057 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPB0 net057 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 Y A0 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 Y A1 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 Y A2 net057 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI33X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN16_2 Y B0 net49__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN17_2 net49__2 B1 net55__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN18_2 net55__2 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN18 net55 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN17 net49 B1 net55 VPW n12 l=1.3e-07 w=7.1e-07
MXN16 Y B0 net49 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_2 Y A0 net43__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN20_2 net43__2 A1 net40__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN19_2 net40__2 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN19 net40 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN20 net43 A1 net40 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net43 VPW n12 l=1.3e-07 w=7.1e-07
MXPB0 net057 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16 net057 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17 net057 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net057 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 net057 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPB0_2 net057 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP20 Y A0 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP19 Y A1 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP18 Y A2 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A2 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_2 Y A1 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 Y A0 net057 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI33XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN13 net55 B2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net49 B1 net55 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 Y B0 net49 VPW n12 l=1.3e-07 w=1.8e-07
MXNA0 Y A0 net43 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net43 A1 net40 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net40 A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP17 net057 B2 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP16 net057 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXPB0 net057 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP20 Y A0 net057 VNW p12 l=1.3e-07 w=3.6e-07
MXP19 Y A1 net057 VNW p12 l=1.3e-07 w=3.6e-07
MXP18 Y A2 net057 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT BUFX10MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT BUFX12MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT BUFX14MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT BUFX16MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX18MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT BUFX20MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT BUFX24MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_5 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_11 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_12 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_5 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_11 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_12 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX2MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX32MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_5 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_6 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_7 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_11 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_12 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_13 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_14 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_15 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_16 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_5 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_6 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_7 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_11 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_12 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_13 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_14 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_15 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_16 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX3MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=7.2e-07
.ends


.SUBCKT BUFX4MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX5MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3.8e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=4.6e-07
.ends


.SUBCKT BUFX6MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX8MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKAND2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1_3 ny A XI0_n1__3 VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=1.05e-06
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=1.05e-06
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=1.05e-06
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=1.05e-06
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X16MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1_3 ny A XI0_n1__3 VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=5.55e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=5.55e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=5.55e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=5.55e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.32e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.5e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X3MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKAND2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=4e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=3.05e-07
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=3.05e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=3.05e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3.05e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=1.04e-06
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=1.04e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=5.45e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=5.45e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX12MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX16MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX1MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=5.1e-07
.ends


.SUBCKT CLKBUFX20MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX24MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=1.03e-06
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=1.03e-06
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKBUFX2MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX32MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_11 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_11 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_12 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX3MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT CLKBUFX40MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_11 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_12 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_13 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_14 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI0_MXPA1_5 ny A VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_11 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_12 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_13 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_14 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX4MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX6MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=2.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKBUFX8MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKINVX12MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX16MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX1MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=2.55e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=5e-07
.ends


.SUBCKT CLKINVX20MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX24MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=5.6e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=5.6e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=9.2e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=9.2e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=9.2e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=9.2e-07
.ends


.SUBCKT CLKINVX2MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX32MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=1.005e-06
mXI0_MXPA1_11 Y A VDD VNW p12 l=1.3e-07 w=1.005e-06
mXI0_MXPA1_12 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX3MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.4e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT CLKINVX40MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_10 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_11 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_12 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_13 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_14 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_15 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_16 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_17 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_11 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_12 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_13 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_14 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_15 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_16 Y A VDD VNW p12 l=1.3e-07 w=8.65e-07
mXI0_MXPA1_17 Y A VDD VNW p12 l=1.3e-07 w=8.65e-07
.ends


.SUBCKT CLKINVX4MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.85e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.85e-07
.ends


.SUBCKT CLKINVX6MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX8MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7.25e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.25e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7.25e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=7.25e-07
.ends


.SUBCKT CLKMX2X12MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g0_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g0_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g0_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X16MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=6.8e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X2MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=2.5e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=7e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X3MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=4.5e-07
.ends


.SUBCKT CLKMX2X4MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X6MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X8MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKNAND2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=6.5e-07
.ends


.SUBCKT CLKNAND2X16MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA2_4 XI0_n1__4 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_4 Y A XI0_n1__4 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_5 Y A XI0_n1__5 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_5 XI0_n1__5 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_6 XI0_n1__6 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_6 Y A XI0_n1__6 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_7 Y A XI0_n1__7 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_7 XI0_n1__7 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_8 XI0_n1__8 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_8 Y A XI0_n1__8 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_7 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_8 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
.ends


.SUBCKT CLKNAND2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8e-07
.ends


.SUBCKT CLKNAND2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.2e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.2e-07
.ends


.SUBCKT CLKNAND2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=7e-07
.ends


.SUBCKT CLKXOR2X12MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g3_MXNA1_2 nB B VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g3_MXNA1_3 nB B VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g2_MXNA1_2 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g2_MXNA1_3 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=3.8e-07
mXI6_MXNOE_2 ny A bB VPW n12 l=1.3e-07 w=3.8e-07
mXI6_MXNOE_3 ny A bB VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=3.8e-07
mXI5_MXNOE_2 ny nA nB VPW n12 l=1.3e-07 w=3.8e-07
mXI5_MXNOE_3 ny nA nB VPW n12 l=1.3e-07 w=4e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.65e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3e-07
mX_g0_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1_2 nB B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 nB B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 nB B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_5 nB B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=1.09e-06
mX_g2_MXPA1_2 bB nB VDD VNW p12 l=1.3e-07 w=1.09e-06
mX_g2_MXPA1_3 bB nB VDD VNW p12 l=1.3e-07 w=1.09e-06
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=8.1e-07
mXI6_MXPOEN_2 ny nA bB VNW p12 l=1.3e-07 w=8.3e-07
mXI6_MXPOEN_3 ny nA bB VNW p12 l=1.3e-07 w=8.3e-07
mXI6_MXPOEN_4 ny nA bB VNW p12 l=1.3e-07 w=8.3e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=8.3e-07
mXI5_MXPOEN_2 ny A nB VNW p12 l=1.3e-07 w=8.3e-07
mXI5_MXPOEN_3 ny A nB VNW p12 l=1.3e-07 w=8.3e-07
mXI5_MXPOEN_4 ny A nB VNW p12 l=1.3e-07 w=8.1e-07
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=1.04e-06
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.05e-06
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.05e-06
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.05e-06
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=3.4e-07
.ends


.SUBCKT CLKXOR2X16MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g3_MXNA1_2 nB B VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g3_MXNA1_3 nB B VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g3_MXNA1_4 nB B VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=5e-07
mX_g2_MXNA1_2 bB nB VSS VPW n12 l=1.3e-07 w=5e-07
mX_g2_MXNA1_3 bB nB VSS VPW n12 l=1.3e-07 w=5e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=5.2e-07
mXI6_MXNOE_2 ny A bB VPW n12 l=1.3e-07 w=5.2e-07
mXI6_MXNOE_3 ny A bB VPW n12 l=1.3e-07 w=5.2e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE_2 ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE_3 ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE_4 ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=1.6e-07
mX_g1_MXNA1_2 nA A VSS VPW n12 l=1.3e-07 w=1.6e-07
mX_g1_MXNA1_3 nA A VSS VPW n12 l=1.3e-07 w=1.6e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=5.45e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=5.45e-07
mX_g0_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g0_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g0_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g3_MXPA1_2 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_3 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_4 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_5 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_6 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_7 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=1.08e-06
mX_g2_MXPA1_2 bB nB VDD VNW p12 l=1.3e-07 w=1.08e-06
mX_g2_MXPA1_3 bB nB VDD VNW p12 l=1.3e-07 w=1.08e-06
mX_g2_MXPA1_4 bB nB VDD VNW p12 l=1.3e-07 w=1.08e-06
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=8.9e-07
mXI6_MXPOEN_2 ny nA bB VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN_3 ny nA bB VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN_4 ny nA bB VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN_5 ny nA bB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN_2 ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN_3 ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN_4 ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN_5 ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=1.33e-06
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.55e-07
.ends


.SUBCKT CLKXOR2X2MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=1.9e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.55e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=5.5e-07
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=4.5e-07
.ends


.SUBCKT CLKXOR2X4MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=5.9e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g3_MXPA1_2 nB B VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g2_MXPA1_2 bB nB VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPOEN_2 ny nA bB VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN_2 ny A nB VNW p12 l=1.3e-07 w=5.5e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=4.5e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=4.5e-07
.ends


.SUBCKT CLKXOR2X8MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=7e-07
mX_g3_MXNA1_2 nB B VSS VPW n12 l=1.3e-07 w=7e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g2_MXNA1_2 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=3.9e-07
mXI6_MXNOE_2 ny A bB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE_2 ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=6.85e-07
mX_g3_MXPA1_2 nB B VDD VNW p12 l=1.3e-07 w=6.85e-07
mX_g3_MXPA1_3 nB B VDD VNW p12 l=1.3e-07 w=6.85e-07
mX_g3_MXPA1_4 nB B VDD VNW p12 l=1.3e-07 w=6.85e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g2_MXPA1_2 bB nB VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN_2 ny nA bB VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN_3 ny nA bB VNW p12 l=1.3e-07 w=7.3e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=7.3e-07
mXI5_MXPOEN_2 ny A nB VNW p12 l=1.3e-07 w=7.3e-07
mXI5_MXPOEN_3 ny A nB VNW p12 l=1.3e-07 w=7.3e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=9.2e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.8e-07
.ends


.SUBCKT DFFHQNX1MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFHQNX2MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQNX4MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=6.1e-07
.ends


.SUBCKT DFFHQNX8MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_3 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_4 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_3 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_4 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQX1MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=3.4e-07
MXN3 net87 cn VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP4 net061 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm nmin net62 VNW p12 l=1.3e-07 w=4.1e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.4e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFHQX2MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=4.8e-07
MXN4 net87 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP6 net061 c cn VNW p12 l=1.3e-07 w=4.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP7 pm nmin net62 VNW p12 l=1.3e-07 w=5.9e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.4e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQX4MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net87 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP8 net061 c cn VNW p12 l=1.3e-07 w=7.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP9 pm nmin net62 VNW p12 l=1.3e-07 w=8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI36_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQX8MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=4.4e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net87 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=7.3e-07
MXP10 net061 c cn VNW p12 l=1.3e-07 w=7.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=8.5e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP9 pm nmin net62 VNW p12 l=1.3e-07 w=8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI36_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=7.3e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHX1MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net42 cn VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP5 net63 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP2 net53 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP6 pm nmin net53 VNW p12 l=1.3e-07 w=4.4e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.9e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFHX2MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=5.1e-07
MXN4 net42 cn VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP7 net63 c cn VNW p12 l=1.3e-07 w=4.6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8e-07
MXP8 net53 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP10 pm nmin net53 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI32_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.1e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT DFFHX4MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=7e-07
MXN5 net42 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP11 net63 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP8 net53 c VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP12 pm nmin net53 VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI32_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT DFFHX8MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=7e-07
MXN5 net42 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP11 net63 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP8 net53 c VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP12 pm nmin net53 VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI32_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT DFFNHX1MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=4.3e-07
MXN2 net67 cn VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net56 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=6.8e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP3 pm net150 net42 VNW p12 l=1.3e-07 w=3.3e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.8e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNHX2MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=6.1e-07
MXN3 net67 cn VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net56 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1_2 cn nckn VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP4 pm net150 net42 VNW p12 l=1.3e-07 w=4.6e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNHX4MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=5.4e-07
MXN3 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN3_2 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 pm net150 net67 VPW n12 l=1.3e-07 w=5.4e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI37_MXNOE_2 bm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP5 net56 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=6.6e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g10_MXPA1_2 cn nckn VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 pm net150 net42 VNW p12 l=1.3e-07 w=6.9e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI37_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mXI52_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNHX8MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=5e-07
mX_g13_MXNA1_2 net150 D VSS VPW n12 l=1.3e-07 w=5e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=7.4e-07
MXN3 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN3_2 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 pm net150 net67 VPW n12 l=1.3e-07 w=5.7e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI37_MXNOE_2 bm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP7 net56 cn c VNW p12 l=1.3e-07 w=6.4e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g13_MXPA1_2 net150 D VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g10_MXPA1_2 cn nckn VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 pm net150 net42 VNW p12 l=1.3e-07 w=6.9e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI37_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mXI52_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI52_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI52_MXPA1_5 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNSRHX1MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS SN net68 VPW n12 l=1.3e-07 w=4.3e-07
MXN11 net68 cn net72 VPW n12 l=1.3e-07 w=4.3e-07
MXN0 pm nmin net72 VPW n12 l=1.3e-07 w=4.3e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 m pm net80 VPW n12 l=1.3e-07 w=4.5e-07
MXN13 VSS RN net80 VPW n12 l=1.3e-07 w=4.5e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
MXN7 bm cn net91 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net91 RN net88 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net88 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net152 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP13 net152 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmin net118 VNW p12 l=1.3e-07 w=3.3e-07
MXP9 net118 c VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=4.8e-07
MXP1 net142 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net142 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.8e-07
MXP16 bm nmset net154 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net154 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP18 bm c net110 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net110 nmset net114 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net114 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT DFFNSRHX2MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS SN net70 VPW n12 l=1.3e-07 w=6e-07
MXN16 net70 cn net66 VPW n12 l=1.3e-07 w=6e-07
MXN0 pm nmin net66 VPW n12 l=1.3e-07 w=6e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 m pm net78 VPW n12 l=1.3e-07 w=6.3e-07
MXN18 VSS RN net78 VPW n12 l=1.3e-07 w=6.3e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.6e-07
MXN7 bm cn net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net89 RN net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net154 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP13 net154 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 pm nmin net120 VNW p12 l=1.3e-07 w=4.6e-07
MXP9 net120 c VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP1 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP20 bm nmset net104 VNW p12 l=1.3e-07 w=2.8e-07
MXP4 net104 RN VDD VNW p12 l=1.3e-07 w=2.8e-07
MXP18 bm c net112 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net112 nmset net116 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net116 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFNSRHX4MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=3e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN20 VSS SN net67 VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net67 cn net71 VPW n12 l=1.3e-07 w=7.5e-07
MXN0 pm nmin net71 VPW n12 l=1.3e-07 w=7.5e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 m pm net79 VPW n12 l=1.3e-07 w=8.4e-07
MXN21 VSS RN net79 VPW n12 l=1.3e-07 w=8.4e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN7 bm cn net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net90 RN net87 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net87 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net155 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP21 net155 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.6e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP22 pm nmin net121 VNW p12 l=1.3e-07 w=6.9e-07
MXP9 net121 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP11_2 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP1 net145 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net145 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP23 bm nmset net105 VNW p12 l=1.3e-07 w=3.6e-07
MXP4 net105 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP18 bm c net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net113 nmset net117 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net117 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFNSRHX8MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g10_MXNA1_2 cn nck VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN20 VSS SN net66 VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net66 cn net70 VPW n12 l=1.3e-07 w=7.5e-07
MXN0 pm nmin net70 VPW n12 l=1.3e-07 w=7.5e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=2.5e-07
MXN4 m pm net78 VPW n12 l=1.3e-07 w=8.7e-07
MXN22 VSS RN net78 VPW n12 l=1.3e-07 w=8.7e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN7 bm cn net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net89 RN net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=3e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP2 net154 CKN VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP24 net154 cn c VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g10_MXPA1_2 cn nck VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=1.03e-06
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP22 pm nmin net120 VNW p12 l=1.3e-07 w=6.9e-07
MXP9 net120 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP11_2 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP1 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP25 bm nmset net104 VNW p12 l=1.3e-07 w=3.5e-07
MXP4 net104 RN VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP18 bm c net112 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net112 nmset net116 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net116 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQNX1MTR QN VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE nm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE nm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN nm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN nm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFQNX2MTR QN VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE nm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE nm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN nm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN nm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQNX4MTR QN VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE nm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE nm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN nm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN nm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQX1MTR Q VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI6_MXNOE ns c XI6_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI7_MXNOE ns cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI6_MXPOEN ns cn XI6_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI7_MXPOEN ns c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFQX2MTR Q VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI6_MXNOE ns c XI6_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI7_MXNOE ns cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI6_MXPOEN ns cn XI6_p1 VNW p12 l=1.3e-07 w=4.9e-07
mXI7_MXPOEN ns c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g1_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQX4MTR Q VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI6_MXNOE ns c XI6_n1 VPW n12 l=1.3e-07 w=4.2e-07
mXI7_MXNOE ns cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI6_MXPOEN ns cn XI6_p1 VNW p12 l=1.3e-07 w=6.1e-07
mXI7_MXPOEN ns c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g1_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRHQX1MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net89 cn VSS VPW n12 l=1.3e-07 w=3.5e-07
MXN2 pm nmin net89 VPW n12 l=1.3e-07 w=3.5e-07
MXN3 pm c net66 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net66 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net73 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
MXN11 m pm net73 VPW n12 l=1.3e-07 w=4.9e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=3.7e-07
MXN7 bm cn net85 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net85 RN net82 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net82 VPW n12 l=1.3e-07 w=1.5e-07
mXI52_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net126 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP11 net126 c cn VNW p12 l=1.3e-07 w=4.2e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP2 net134 c VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP12 pm nmin net134 VNW p12 l=1.3e-07 w=4.2e-07
MXP14 pm cn net104 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 VDD m net104 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.3e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP16 bm c net120 VNW p12 l=1.3e-07 w=2.3e-07
MXP15 VDD s net120 VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFRHQX2MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net90 cn VSS VPW n12 l=1.3e-07 w=5.1e-07
MXN2 pm nmin net90 VPW n12 l=1.3e-07 w=5.1e-07
MXN3 pm c net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 net74 RN VSS VPW n12 l=1.3e-07 w=6.8e-07
MXN11 m pm net74 VPW n12 l=1.3e-07 w=6.8e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.4e-07
MXN7 bm cn net86 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net86 RN net83 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net83 VPW n12 l=1.3e-07 w=1.5e-07
mXI50_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI51_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net131 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP18 net131 c cn VNW p12 l=1.3e-07 w=4.5e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP19 pm nmin net105 VNW p12 l=1.3e-07 w=6.2e-07
MXP20 pm cn net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP5 VDD m net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=8.5e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.1e-07
mXI58_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=5.3e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=2.7e-07
MXP21 bm c net125 VNW p12 l=1.3e-07 w=1.5e-07
MXP15 VDD s net125 VNW p12 l=1.3e-07 w=1.5e-07
mXI50_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRHQX4MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MXN15 net90 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm nmin net90 VPW n12 l=1.3e-07 w=5.1e-07
MXN3 pm c net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net74 RN VSS VPW n12 l=1.3e-07 w=5.9e-07
MXN11 m pm net74 VPW n12 l=1.3e-07 w=5.9e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MXN7 bm cn net86 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net86 RN net83 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net83 VPW n12 l=1.3e-07 w=1.5e-07
mXI50_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net131 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP18 net131 c cn VNW p12 l=1.3e-07 w=4.5e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
MXP2 net105 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP19 pm nmin net105 VNW p12 l=1.3e-07 w=6.2e-07
MXP20 pm cn net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP5 VDD m net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP6_2 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI58_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=3e-07
MXP21 bm c net125 VNW p12 l=1.3e-07 w=1.5e-07
MXP15 VDD s net125 VNW p12 l=1.3e-07 w=1.5e-07
mXI50_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRHQX8MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MXN15 net90 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm nmin net90 VPW n12 l=1.3e-07 w=5.1e-07
MXN3 pm c net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net74 RN VSS VPW n12 l=1.3e-07 w=5.9e-07
MXN11 m pm net74 VPW n12 l=1.3e-07 w=5.9e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MXN7 bm cn net86 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net86 RN net83 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net83 VPW n12 l=1.3e-07 w=1.5e-07
mXI50_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net131 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP18 net131 c cn VNW p12 l=1.3e-07 w=4.5e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
MXP2 net105 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP19 pm nmin net105 VNW p12 l=1.3e-07 w=6.2e-07
MXP20 pm cn net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP5 VDD m net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP6_2 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI58_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=3e-07
MXP21 bm c net125 VNW p12 l=1.3e-07 w=1.5e-07
MXP15 VDD s net125 VNW p12 l=1.3e-07 w=1.5e-07
mXI50_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRQX1MTR Q VDD VNW VPW VSS CK D RN
MXN5 net86 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net78 D net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 pm cn net78 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 pm c net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net66 m net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net66 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI37_MXNOE net119 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE net119 cn XI4_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 s net119 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP4 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 D VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP6 pm c net105 VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI37_MXPOEN net119 cn m VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN net119 c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 s net119 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFRQX2MTR Q VDD VNW VPW VSS CK D RN
MXN5 net86 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net78 D net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 pm cn net78 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 pm c net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net66 m net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net66 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI37_MXNOE net119 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE net119 cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 s net119 XI0_n1 VPW n12 l=1.3e-07 w=2.7e-07
mXI0_MXNA2 XI0_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 D VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP6 pm c net105 VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3e-07
mXI37_MXPOEN net119 cn m VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN net119 c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 s net119 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRQX4MTR Q VDD VNW VPW VSS CK D RN
MXN5 net86 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net78 D net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 pm cn net78 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 pm c net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net66 m net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net66 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI37_MXNOE net119 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE net119 cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 s net119 XI0_n1 VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA2 XI0_n1 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 D VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP6 pm c net105 VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3e-07
mXI37_MXPOEN net119 cn m VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN net119 c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 s net119 VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRX1MTR Q QN VDD VNW VPW VSS CK D RN
MXN2 pm cn net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net45 D net53 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net53 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 pm c net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net61 m net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net61 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE bm cn XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 net90 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 net90 bm XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI45_MXNA1 Q net90 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP2 net68 D VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm c net68 VNW p12 l=1.3e-07 w=4.1e-07
MXP1 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MXP7 pm cn net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD m net72 VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI40_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI5_MXPOEN bm c XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 net90 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 net90 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 net90 bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI45_MXPA1 Q net90 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFRX2MTR Q QN VDD VNW VPW VSS CK D RN
MXN2 pm cn net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net45 D net53 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net53 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 pm c net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net61 m net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net61 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE bm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 net90 VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1 net90 bm XI1_n1 VPW n12 l=1.3e-07 w=2.7e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI45_MXNA1 Q net90 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP2 net68 D VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm c net68 VNW p12 l=1.3e-07 w=4.1e-07
MXP1 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 pm cn net72 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 VDD m net72 VNW p12 l=1.3e-07 w=2.2e-07
mXI43_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI40_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI5_MXPOEN bm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 net90 VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 net90 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 net90 bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI45_MXPA1 Q net90 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRX4MTR Q QN VDD VNW VPW VSS CK D RN
MXN2 pm cn net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net45 D net53 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net53 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 pm c net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net61 m net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net61 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE bm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 net90 VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1 net90 bm XI1_n1 VPW n12 l=1.3e-07 w=4.9e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI46_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI45_MXNA1 Q net90 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI45_MXNA1_2 Q net90 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP2 net68 D VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm c net68 VNW p12 l=1.3e-07 w=4.1e-07
MXP1 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 pm cn net72 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 VDD m net72 VNW p12 l=1.3e-07 w=2.2e-07
mXI43_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI40_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI5_MXPOEN bm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 net90 VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 net90 RN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 net90 bm VDD VNW p12 l=1.3e-07 w=3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI46_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI45_MXPA1 Q net90 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI45_MXPA1_2 Q net90 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSHQX1MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 VSS SN net92 VPW n12 l=1.3e-07 w=4.5e-07
MXN7 net92 cn net89 VPW n12 l=1.3e-07 w=4.5e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP7 net099 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 pm nmin net091 VNW p12 l=1.3e-07 w=3.7e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT DFFSHQX2MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS SN net92 VPW n12 l=1.3e-07 w=6.4e-07
MXN11 net92 cn net89 VPW n12 l=1.3e-07 w=6.4e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=6.4e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP13 net099 c cn VNW p12 l=1.3e-07 w=4.9e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmin net091 VNW p12 l=1.3e-07 w=5.4e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSHQX4MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN14 VSS SN net92 VPW n12 l=1.3e-07 w=7.5e-07
MXN13 net92 cn net89 VPW n12 l=1.3e-07 w=7.5e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=7.5e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP15 net099 c cn VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP16 pm nmin net091 VNW p12 l=1.3e-07 w=6.9e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSHQX8MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN14 VSS SN net92 VPW n12 l=1.3e-07 w=7.5e-07
MXN13 net92 cn net89 VPW n12 l=1.3e-07 w=7.5e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=7.5e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP15 net099 c cn VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP16 pm nmin net091 VNW p12 l=1.3e-07 w=6.9e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSQX1MTR Q VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN2 bm cn net84 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 NSN s net84 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI34_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm c net62 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD s net62 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSQX2MTR Q VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN2 bm cn net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 NSN s net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN1 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI34_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 bm c net53 VNW p12 l=1.3e-07 w=1.5e-07
MXP7 VDD s net53 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSQX4MTR Q VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN2 bm cn net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 NSN s net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN1 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI34_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 bm c net53 VNW p12 l=1.3e-07 w=1.5e-07
MXP7 VDD s net53 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRHQX1MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 VSS SN net62 VPW n12 l=1.3e-07 w=4.1e-07
MXN12 net62 cn net82 VPW n12 l=1.3e-07 w=4.1e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=4.1e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=4.3e-07
MXN14 VSS RN net70 VPW n12 l=1.3e-07 w=4.3e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net122 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 pm nmin net128 VNW p12 l=1.3e-07 w=3.1e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP17 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.6e-07
MXP23 bm nmset net112 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSRHQX2MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN21 VSS SN net62 VPW n12 l=1.3e-07 w=5.8e-07
MXN20 net62 cn net82 VPW n12 l=1.3e-07 w=5.8e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=5.8e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=6.1e-07
MXN22 VSS RN net70 VPW n12 l=1.3e-07 w=6.1e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net122 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP25 pm nmin net128 VNW p12 l=1.3e-07 w=4.5e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP17 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP27 bm nmset net112 VNW p12 l=1.3e-07 w=2.7e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRHQX4MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS SN net62 VPW n12 l=1.3e-07 w=7.5e-07
MXN23 net62 cn net82 VPW n12 l=1.3e-07 w=7.5e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=7.5e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN25 VSS RN net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP28 net122 c cn VNW p12 l=1.3e-07 w=6.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.03e-06
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP29 pm nmin net128 VNW p12 l=1.3e-07 w=6.8e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP30 m RN net144 VNW p12 l=1.3e-07 w=3.1e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP31 bm nmset net112 VNW p12 l=1.3e-07 w=3.6e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRHQX8MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS SN net62 VPW n12 l=1.3e-07 w=7.5e-07
MXN23 net62 cn net82 VPW n12 l=1.3e-07 w=7.5e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=7.5e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN25 VSS RN net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP28 net122 c cn VNW p12 l=1.3e-07 w=6.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.03e-06
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP29 pm nmin net128 VNW p12 l=1.3e-07 w=6.8e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP30 m RN net144 VNW p12 l=1.3e-07 w=3.1e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP31 bm nmset net112 VNW p12 l=1.3e-07 w=3.6e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRX1MTR Q QN VDD VNW VPW VSS CK D RN SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm c XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MXN2 m NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MXN3 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MXN8 bm cn net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 NSN s net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm cn XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net_NRN NRN VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP6 m pm net_NRN VNW p12 l=1.3e-07 w=3.6e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MXP7 bm c net75 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net_NRN s net75 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSRX2MTR Q QN VDD VNW VPW VSS CK D RN SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm c XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MXN2 m NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MXN3 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MXN4 bm cn net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 NSN s net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm cn XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net_NRN NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 m pm net_NRN VNW p12 l=1.3e-07 w=4.4e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.4e-07
MXP7 bm c net75 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net_NRN s net75 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRX4MTR Q QN VDD VNW VPW VSS CK D RN SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI4_MXNOE pm c XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MXN2 m NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=4.7e-07
MXN3 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MXN4 bm cn net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 NSN s net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN SN VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm cn XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net_NRN NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 m pm net_NRN VNW p12 l=1.3e-07 w=4.4e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.7e-07
MXP7 bm c net75 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net_NRN s net75 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSX1MTR Q QN VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm BSN VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MXN1 bm cn net134 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 BSN s net134 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 BSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net73 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSX2MTR Q QN VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN0 m pm BSN VPW n12 l=1.3e-07 w=2.1e-07
MXN0_2 m pm BSN VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MXN1 bm cn net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN4 BSN s net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.1e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm c net73 VNW p12 l=1.3e-07 w=1.5e-07
MXP6 VDD s net73 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSX4MTR Q QN VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=2e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=2e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 m pm BSN VPW n12 l=1.3e-07 w=3.3e-07
MXN0_2 m pm BSN VPW n12 l=1.3e-07 w=3.3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=5.2e-07
MXN1 bm cn net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN4 BSN s net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN SN VSS VPW n12 l=1.3e-07 w=1.08e-06
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=5.6e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.4e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.2e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm c net73 VNW p12 l=1.3e-07 w=1.5e-07
MXP6 VDD s net73 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFTRX1MTR Q QN VDD VNW VPW VSS CK D RN
MXN4 net129 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net132 D net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm cn net132 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
mXI4_MXNOE bm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g11_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP4 net62 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm c net62 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI4_MXPOEN bm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g11_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFTRX2MTR Q QN VDD VNW VPW VSS CK D RN
MXN6 net129 RN VSS VPW n12 l=1.3e-07 w=2.6e-07
MXN5 net132 D net129 VPW n12 l=1.3e-07 w=2.6e-07
MXN1 pm cn net132 VPW n12 l=1.3e-07 w=2.6e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI4_MXNOE bm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g11_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 net62 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP5 pm c net62 VNW p12 l=1.3e-07 w=2.6e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.7e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI4_MXPOEN bm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g11_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFTRX4MTR Q QN VDD VNW VPW VSS CK D RN
MXN8 net129 RN VSS VPW n12 l=1.3e-07 w=5e-07
MXN7 net132 D net129 VPW n12 l=1.3e-07 w=5e-07
MXN1 pm cn net132 VPW n12 l=1.3e-07 w=5e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=4e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=8e-07
mXI4_MXNOE bm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g11_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g11_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 net62 RN VDD VNW p12 l=1.3e-07 w=2.5e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP6 pm c net62 VNW p12 l=1.3e-07 w=5.1e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.6e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_3 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_4 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI47_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI4_MXPOEN bm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g11_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g11_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFX1MTR Q QN VDD VNW VPW VSS CK D
mXI14_MXNA1 XI14_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNOE pm cn XI14_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI12_MXNOE nm c XI12_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI11_MXNOE nm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI14_MXPA1 XI14_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI14_MXPOEN pm c XI14_p1 VNW p12 l=1.3e-07 w=3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI12_MXPOEN nm cn XI12_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI11_MXPOEN nm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFX2MTR Q QN VDD VNW VPW VSS CK D
mXI14_MXNA1 XI14_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNOE pm cn XI14_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=4e-07
mXI12_MXNOE nm c XI12_n1 VPW n12 l=1.3e-07 w=4e-07
mXI11_MXNOE nm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1 XI14_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI14_MXPOEN pm c XI14_p1 VNW p12 l=1.3e-07 w=3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=4.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI12_MXPOEN nm cn XI12_p1 VNW p12 l=1.3e-07 w=4.9e-07
mXI11_MXPOEN nm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFX4MTR Q QN VDD VNW VPW VSS CK D
mXI14_MXNA1 XI14_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNOE pm cn XI14_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=5.8e-07
mXI12_MXNOE nm c XI12_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI11_MXNOE nm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1 XI14_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI14_MXPOEN pm c XI14_p1 VNW p12 l=1.3e-07 w=3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g14_MXPA1_2 cn CK VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.7e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI12_MXPOEN nm cn XI12_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI11_MXPOEN nm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DLY1X1MTR Y VDD VNW VPW VSS A
mX_g1_MXNA1 nmin A VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 nmin1 nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 ny nmin1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 nmin A VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 nmin1 nmin VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 ny nmin1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=5.1e-07
.ends


.SUBCKT DLY1X4MTR Y VDD VNW VPW VSS A
mX_g1_MXNA1 nmin A VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN1 nmin1 nmin VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN3 ny nmin1 VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 nmin A VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP2 nmin1 nmin VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP3 ny nmin1 VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DLY2X1MTR Y VDD VNW VPW VSS A
mXI0_MXNOE ny A XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 A VSS VPW n12 l=1.3e-07 w=1.5e-07
MXN0 VSS ny VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN ny A XI0_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI0_MXPA1 XI0_p1 A VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP0 VDD ny VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DLY2X4MTR Y VDD VNW VPW VSS A
mXI0_MXNOE ny A XI0_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI0_MXNA1 XI0_n1 A VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN0 VSS ny VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPOEN ny A XI0_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA1 XI0_p1 A VDD VNW p12 l=1.3e-07 w=6.5e-07
MXP0 VDD ny VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DLY3X1MTR Y VDD VNW VPW VSS A
mX_g1_MXNA1 nmin A VSS VPW n12 l=1.3e-07 w=1.5e-07
MXN6 net64 nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net70 nmin net64 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 nmin1 nmin net70 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 ny nmin1 net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net67 nmin1 net61 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net61 nmin1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXPA1 nmin A VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP2 net51 nmin VDD VNW p12 l=1.3e-07 w=3.15e-07
MXP0 net36 nmin net51 VNW p12 l=1.3e-07 w=3.15e-07
MXP1 nmin1 nmin net36 VNW p12 l=1.3e-07 w=3.15e-07
MXP5 ny nmin1 net39 VNW p12 l=1.3e-07 w=3.15e-07
MXP4 net39 nmin1 net48 VNW p12 l=1.3e-07 w=3.15e-07
MXP3 net48 nmin1 VDD VNW p12 l=1.3e-07 w=3.15e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DLY3X4MTR Y VDD VNW VPW VSS A
mX_g1_MXNA1 nmin A VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN6 net64 nmin VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN0 net70 nmin net64 VPW n12 l=1.3e-07 w=4.2e-07
MXN1 nmin1 nmin net70 VPW n12 l=1.3e-07 w=4.2e-07
MXN3 ny nmin1 net67 VPW n12 l=1.3e-07 w=4.2e-07
MXN4 net67 nmin1 net61 VPW n12 l=1.3e-07 w=4.2e-07
MXN5 net61 nmin1 VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmin A VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP2 net51 nmin VDD VNW p12 l=1.3e-07 w=7.2e-07
MXP0 net36 nmin net51 VNW p12 l=1.3e-07 w=7.2e-07
MXP1 nmin1 nmin net36 VNW p12 l=1.3e-07 w=7.2e-07
MXP5 ny nmin1 net39 VNW p12 l=1.3e-07 w=7.2e-07
MXP4 net39 nmin1 net48 VNW p12 l=1.3e-07 w=7.2e-07
MXP3 net48 nmin1 VDD VNW p12 l=1.3e-07 w=7.2e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DLY4X1MTR Y VDD VNW VPW VSS A
mXI0_MXNOE na A XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 A VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 na VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNOE ba na XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNOE nba ba XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 ba VSS VPW n12 l=1.3e-07 w=1.5e-07
MXN0 VSS nba VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI3_MXNA1 Y nba VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN na A XI0_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI0_MXPA1 XI0_p1 A VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 na VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPOEN ba na XI1_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI2_MXPOEN nba ba XI2_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI2_MXPA1 XI2_p1 ba VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP0 VDD nba VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI3_MXPA1 Y nba VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DLY4X4MTR Y VDD VNW VPW VSS A
mXI0_MXNOE na A XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 A VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 na VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI1_MXNOE ba na XI1_n1 VPW n12 l=1.3e-07 w=2.2e-07
mXI2_MXNOE nba ba XI2_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI2_MXNA1 XI2_n1 ba VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN0 VSS nba VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI3_MXNA1 Y nba VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 Y nba VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPOEN na A XI0_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI0_MXPA1 XI0_p1 A VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 na VDD VNW p12 l=1.3e-07 w=3.75e-07
mXI1_MXPOEN ba na XI1_p1 VNW p12 l=1.3e-07 w=3.75e-07
mXI2_MXPOEN nba ba XI2_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI2_MXPA1 XI2_p1 ba VDD VNW p12 l=1.3e-07 w=6.5e-07
MXP0 VDD nba VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI3_MXPA1 Y nba VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 Y nba VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFHQX1MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 VSS s net104 VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=3.6e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=4e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=3e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 nmsi E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=4.5e-07
MXP0 cn c net053 VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP2 pm nmsi net047 VNW p12 l=1.3e-07 w=4.4e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=7.9e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT EDFFHQX2MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 VSS s net104 VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=5.1e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.2e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.6e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=3.9e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 nmsi E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=4.5e-07
MXP0 cn c net053 VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=8e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 pm nmsi net047 VNW p12 l=1.3e-07 w=6.2e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFHQX4MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=2.3e-07
MXN3 VSS s net104 VPW n12 l=1.3e-07 w=2.3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=5.1e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmsi E net73 VNW p12 l=1.3e-07 w=2.8e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=5e-07
MXP4 cn c net053 VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 pm nmsi net047 VNW p12 l=1.3e-07 w=6.2e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFHQX8MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=2.3e-07
MXN3 VSS s net104 VPW n12 l=1.3e-07 w=2.3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=5.1e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmsi E net73 VNW p12 l=1.3e-07 w=2.8e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=5e-07
MXP4 cn c net053 VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 pm nmsi net047 VNW p12 l=1.3e-07 w=6.2e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFTRX1MTR Q QN VDD VNW VPW VSS CK D E RN
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net122 s net140 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net122 nmen net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net107 E net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net140 D net107 VPW n12 l=1.3e-07 w=1.8e-07
MX_t3 net106 RN VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t19 pm cn net140 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI11_MXNOE bnm c XI11_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI5_MXNOE bnm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bnm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 net77 s net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 VDD nmen net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net76 D net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 VDD RN net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net77 c pm VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI11_MXPA1 XI11_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI11_MXPOEN bnm cn XI11_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI5_MXPOEN bnm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bnm VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT EDFFTRX2MTR Q QN VDD VNW VPW VSS CK D E RN
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net122 s net140 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net122 nmen net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net107 E net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net140 D net107 VPW n12 l=1.3e-07 w=1.8e-07
MX_t3 net106 RN VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t19 pm cn net140 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 m VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI11_MXNOE bnm c XI11_n1 VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE bnm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g1_MXNA1 Q bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 net77 s net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 VDD nmen net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net76 D net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 VDD RN net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net77 c pm VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI11_MXPA1 XI11_p1 m VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI11_MXPOEN bnm cn XI11_p1 VNW p12 l=1.3e-07 w=5.2e-07
mXI5_MXPOEN bnm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g1_MXPA1 Q bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFTRX4MTR Q QN VDD VNW VPW VSS CK D E RN
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net122 s net140 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net122 nmen net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net107 E net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net140 D net107 VPW n12 l=1.3e-07 w=1.8e-07
MX_t3 net106 RN VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t19 pm cn net140 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 m VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI11_MXNOE bnm c XI11_n1 VPW n12 l=1.3e-07 w=6.3e-07
mXI5_MXNOE bnm cn XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g1_MXNA1 Q bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 net77 s net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 VDD nmen net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net76 D net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 VDD RN net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net77 c pm VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI11_MXPA1 XI11_p1 m VDD VNW p12 l=1.3e-07 w=8.2e-07
mXI11_MXPOEN bnm cn XI11_p1 VNW p12 l=1.3e-07 w=8.2e-07
mXI5_MXPOEN bnm c XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g1_MXPA1 Q bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFX1MTR Q QN VDD VNW VPW VSS CK D E
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net120 s net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net120 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net123 E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net129 D net123 VPW n12 l=1.3e-07 w=1.8e-07
MX_t19 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI1_MXNOE nm c XI1_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net38 s net36 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 VDD E net36 VNW p12 l=1.3e-07 w=3.8e-07
MX_t5 VDD nmen net39 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net39 D net38 VNW p12 l=1.3e-07 w=3.8e-07
MXP2 net38 c pm VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI1_MXPOEN nm cn XI1_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT EDFFX2MTR Q QN VDD VNW VPW VSS CK D E
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net120 s net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net120 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net123 E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net129 D net123 VPW n12 l=1.3e-07 w=1.8e-07
MX_t19 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI1_MXNOE nm c XI1_n1 VPW n12 l=1.3e-07 w=4.3e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net38 s net36 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 VDD E net36 VNW p12 l=1.3e-07 w=3.8e-07
MX_t5 VDD nmen net39 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net39 D net38 VNW p12 l=1.3e-07 w=3.8e-07
MXP2 net38 c pm VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI1_MXPOEN nm cn XI1_p1 VNW p12 l=1.3e-07 w=5.2e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFX4MTR Q QN VDD VNW VPW VSS CK D E
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net120 s net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net120 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net123 E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net129 D net123 VPW n12 l=1.3e-07 w=1.8e-07
MX_t19 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI1_MXNOE nm c XI1_n1 VPW n12 l=1.3e-07 w=6.4e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net38 s net36 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 VDD E net36 VNW p12 l=1.3e-07 w=3.8e-07
MX_t5 VDD nmen net39 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net39 D net38 VNW p12 l=1.3e-07 w=3.8e-07
MXP2 net38 c pm VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.7e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI1_MXPOEN nm cn XI1_p1 VNW p12 l=1.3e-07 w=7.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=5e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends









.SUBCKT FILLCAP16MTR VDD VNW VPW VSS
MXN0 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_2 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_3 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_4 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_5 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_6 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_7 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_8 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_9 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_10 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_11 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXP0 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_2 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_3 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_4 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_5 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_6 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_7 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_8 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_9 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_10 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_11 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
.ends


.SUBCKT FILLCAP32MTR VDD VNW VPW VSS
MXN0 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_2 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_3 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_4 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_5 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_6 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_7 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_8 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_9 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_10 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_11 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_12 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_13 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_14 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_15 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_16 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_17 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_18 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_19 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_20 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_21 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_22 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_23 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXP0 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_2 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_3 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_4 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_5 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_6 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_7 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_8 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_9 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_10 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_11 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_12 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_13 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_14 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_15 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_16 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_17 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_18 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_19 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_20 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_21 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_22 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_23 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
.ends


.SUBCKT FILLCAP4MTR VDD VNW VPW VSS
MXN0 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_2 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXP0 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_2 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
.ends


.SUBCKT FILLCAP64MTR VDD VNW VPW VSS
MXN0 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_2 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_3 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_4 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_5 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_6 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_7 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_8 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_9 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_10 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_11 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_12 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_13 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_14 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_15 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_16 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_17 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_18 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_19 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_20 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_21 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_22 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_23 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_24 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_25 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_26 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_27 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_28 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_29 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_30 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_31 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_32 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_33 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_34 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_35 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_36 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_37 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_38 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_39 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_40 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_41 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_42 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_43 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_44 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_45 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_46 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_47 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXP0 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_2 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_3 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_4 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_5 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_6 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_7 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_8 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_9 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_10 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_11 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_12 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_13 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_14 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_15 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_16 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_17 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_18 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_19 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_20 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_21 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_22 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_23 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_24 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_25 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_26 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_27 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_28 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_29 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_30 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_31 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_32 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_33 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_34 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_35 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_36 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_37 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_38 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_39 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_40 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_41 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_42 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_43 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_44 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_45 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_46 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_47 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
.ends


.SUBCKT FILLCAP8MTR VDD VNW VPW VSS
MXN0 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_2 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_3 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_4 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXN0_5 VSS VDD VSS VPW n12 l=1.3e-07 w=5.85e-07
MXP0 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_2 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_3 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_4 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
MXP0_5 VDD VSS VDD VNW p12 l=1.3e-07 w=7.15e-07
.ends


.SUBCKT INVX10MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX12MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX14MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX16MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX18MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX1MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT INVX20MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_10 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX24MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_10 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_11 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_12 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_11 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_12 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX2MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX32MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_10 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_11 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_12 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_13 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_14 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_15 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_16 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_11 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_12 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_13 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_14 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_15 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_16 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX3MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT INVX4MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX5MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT INVX6MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX8MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVXLMTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MDFFHQX1MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=2.1e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 net135 cn VSS VPW n12 l=1.3e-07 w=3.3e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=3.3e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=3.7e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t9 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=2.6e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=3e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=3e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=4.2e-07
MXP0 cn c net50 VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=4e-07
MXP1 pm nmsi net61 VNW p12 l=1.3e-07 w=4e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=7.3e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MDFFHQX2MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=3.1e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=3e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN1 net135 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=4.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=4.4e-07
MXP2 cn c net50 VNW p12 l=1.3e-07 w=4.4e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=7.6e-07
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP5 pm nmsi net61 VNW p12 l=1.3e-07 w=5.9e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=9.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=9.8e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MDFFHQX4MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=5e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN2 net135 cn VSS VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=5.6e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net50 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net61 VNW p12 l=1.3e-07 w=1.01e-06
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MDFFHQX8MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=4.9e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN2 net135 cn VSS VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=5.6e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.3e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net50 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net61 VNW p12 l=1.3e-07 w=1.01e-06
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2X12MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=7.1e-07
MXN3 nmin nmsel net42 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_5 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_6 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=8.7e-07
MXP1 net42 S0 nmin VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_5 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2X1MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=3.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=3.7e-07
MXN0 nmin nmsel net38 VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 net38 A VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=4.6e-07
MXP0 net38 S0 nmin VNW p12 l=1.3e-07 w=4.6e-07
mX_g2_MXPA1 net38 A VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT MX2X2MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=4.1e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=5.9e-07
MXN0 nmin nmsel net38 VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1 net38 A VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=5.7e-07
MXP0 net38 S0 nmin VNW p12 l=1.3e-07 w=7.4e-07
mX_g2_MXPA1 net38 A VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2X3MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=6.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=6.7e-07
MXN1 nmin nmsel net42 VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net42 S0 nmin VNW p12 l=1.3e-07 w=8.6e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT MX2X4MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=6.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=6.7e-07
MXN1 nmin nmsel net42 VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net42 S0 nmin VNW p12 l=1.3e-07 w=8.6e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2X6MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=6.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=6.7e-07
MXN1 nmin nmsel net42 VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net42 S0 nmin VNW p12 l=1.3e-07 w=8.6e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2X8MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=6.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=6.7e-07
MXN1 nmin nmsel net42 VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net42 S0 nmin VNW p12 l=1.3e-07 w=8.6e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2XLMTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=2.1e-07
MXN1 nmin nmsel net38 VPW n12 l=1.3e-07 w=2.1e-07
mX_g2_MXNA1 net38 A VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=2.5e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=2.5e-07
MXP1 net38 S0 nmin VNW p12 l=1.3e-07 w=2.5e-07
mX_g2_MXPA1 net38 A VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MX3X1MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=4.1e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=4.7e-07
MX_t4 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=5.6e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=1.9e-07
MX_t0 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=4.5e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=3.7e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
MX_t5 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=6.8e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=2.4e-07
MX_t1 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=6.7e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=4.6e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MX3X2MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=5.8e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=6.4e-07
MX_t4 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=6.6e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t0 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=6.5e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=5.9e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=8.7e-07
MX_t5 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=8.8e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=3.4e-07
MX_t1 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=8.8e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=6.9e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX3X4MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=5.8e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=6.4e-07
MX_t4 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=6.6e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t0 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=6.6e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=6.6e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=8.7e-07
MX_t5 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=8.8e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MX_t1 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=8.8e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=7e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=7.6e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX3X8MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=5e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=6.4e-07
MX_t4 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=6.4e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t0 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=6.6e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=5.3e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=7.8e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=7.8e-07
MX_t5 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.6e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=8.6e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=8.6e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=8.6e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX3XLMTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=3.1e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=3.1e-07
MXN0 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=3.1e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=3.1e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=3e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=3.8e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=3.8e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=3.8e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=3e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MX4X1MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI17_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=5.6e-07
MXN0 nmin2in3 nmsel0 net100 VPW n12 l=1.3e-07 w=5.6e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=5.6e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g2_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI18_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=5.6e-07
MXN1 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=5.6e-07
MXN2 nmin0in1 nmsel0 net104 VPW n12 l=1.3e-07 w=5.6e-07
mXI19_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN4 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=5.6e-07
MXN3 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=5.6e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI17_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t9 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=5.9e-07
MX_t11 net98 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=6.8e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g2_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=5.8e-07
mXI18_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t7 net102 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=6.8e-07
mXI19_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=2.9e-07
MXP2 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=6.8e-07
MXP1 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=6.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MX4X2MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI17_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0 nmin2in3 nmsel0 net100 VPW n12 l=1.3e-07 w=7.1e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=6.8e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN1 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=6.8e-07
MXN2 nmin0in1 nmsel0 net104 VPW n12 l=1.3e-07 w=6.9e-07
mXI19_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MXN6 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=6.9e-07
MXN7 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI17_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t9 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=8.6e-07
MX_t11 net98 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI18_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t7 net102 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
MXP3 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.6e-07
mXI19_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP4 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=8.6e-07
MXP1 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=8.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX4X4MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI17_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0 nmin2in3 nmsel0 net100 VPW n12 l=1.3e-07 w=7.1e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=6.8e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN1 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=6.8e-07
MXN2 nmin0in1 nmsel0 net104 VPW n12 l=1.3e-07 w=6.9e-07
mXI19_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MXN7 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI17_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t9 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=8.6e-07
MX_t11 net98 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI18_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t7 net102 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
MXP3 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.6e-07
mXI19_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP4 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=8.6e-07
MXP1 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=8.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX4X8MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI17_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0 nmin2in3 nmsel0 net100 VPW n12 l=1.3e-07 w=7.1e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=6.8e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN1 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=6.8e-07
MXN2 nmin0in1 nmsel0 net104 VPW n12 l=1.3e-07 w=6.9e-07
mXI19_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MXN7 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI17_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t9 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=8.6e-07
MX_t11 net98 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI18_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t7 net102 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
MXP3 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.6e-07
mXI19_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP4 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=8.6e-07
MXP1 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=8.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX4XLMTR Y VDD VNW VPW VSS A B C D S0 S1
mXI20_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN5 nmin2in3 net0110 net100 VPW n12 l=1.3e-07 w=3.1e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=3.1e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 net0110 S0 VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI21_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN6 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=3.1e-07
MXN7 nmin0in1 net0110 net104 VPW n12 l=1.3e-07 w=3.1e-07
mXI22_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=3.1e-07
MXN8 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI20_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=3.8e-07
MX_t11 net98 net0110 nmin2in3 VNW p12 l=1.3e-07 w=3.8e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=3.8e-07
mX_g2_MXPA1 net0110 S0 VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI21_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net102 net0110 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
mXI22_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=3.8e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=3.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MXI2DX1MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=1.9e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=3.7e-07
MXN0 nmin nmsel A VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=4.6e-07
MXP0 A net31 nmin VNW p12 l=1.3e-07 w=4.6e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MXI2DX2MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=2.6e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MXN1 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=4.5e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=3.1e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MXP0 A net31 nmin VNW p12 l=1.3e-07 w=7.4e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2DX4MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=5.2e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MX_t2_2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MXN2 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
MXN2_2 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MX_t3_2 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MXP0 A net31 nmin VNW p12 l=1.3e-07 w=7.1e-07
MXP0_2 A net31 nmin VNW p12 l=1.3e-07 w=7.8e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2DX8MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 nmsel S0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g1_MXNA1_2 net31 nmsel VSS VPW n12 l=1.3e-07 w=5.7e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MX_t2_2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MX_t2_3 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MX_t2_4 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MXN3 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
MXN3_2 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
MXN3_3 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
MXN3_4 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 nmsel S0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g1_MXPA1_2 net31 nmsel VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MX_t3_2 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MX_t3_3 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MX_t3_4 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MXP0 A net31 nmin VNW p12 l=1.3e-07 w=7.2e-07
MXP0_2 A net31 nmin VNW p12 l=1.3e-07 w=7.7e-07
MXP0_3 A net31 nmin VNW p12 l=1.3e-07 w=7.7e-07
MXP0_4 A net31 nmin VNW p12 l=1.3e-07 w=7.3e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_3 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2DXLMTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=1.9e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=3e-07
MXN1 nmin nmsel A VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=3e-07
MXP1 A net31 nmin VNW p12 l=1.3e-07 w=3e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MXI2X12MTR Y VDD VNW VPW VSS A B S0
mXI16_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_3 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_4 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_5 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_6 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1_2 nmsel S0 VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g0_MXNA1_3 nmsel S0 VSS VPW n12 l=1.3e-07 w=5.8e-07
MXN5 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_3 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_4 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_5 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_6 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_3 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_4 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_5 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_6 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_3 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_4 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_5 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_6 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_3 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_4 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_5 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_6 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g0_MXPA1_2 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g0_MXPA1_3 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.5e-07
MXP4 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_3 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_4 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_5 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_6 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_4 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_5 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_6 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_3 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_4 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_5 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_6 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2X1MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y nmsel nmin0 VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=5.3e-07
MX_t1 nmin0 S0 Y VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MXI2X2MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7e-07
MXN0 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
mXI11_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.6e-07
MX_t1 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
mXI11_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2X3MTR Y VDD VNW VPW VSS A B S0
mXI12_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI12_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN1 Y nmsel nmin0 VPW n12 l=1.3e-07 w=5.4e-07
MXN1_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=5.4e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=5.4e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=5.4e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI12_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI12_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=5.6e-07
MXP0 nmin0 S0 Y VNW p12 l=1.3e-07 w=6.6e-07
MXP0_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=6.6e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=5.3e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=7.9e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=6.9e-07
.ends


.SUBCKT MXI2X4MTR Y VDD VNW VPW VSS A B S0
mXI13_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI13_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=6e-07
MXN2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN2_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI13_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI13_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP1 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP1_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2X6MTR Y VDD VNW VPW VSS A B S0
mXI14_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXNA1_3 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g0_MXNA1_2 nmsel S0 VSS VPW n12 l=1.3e-07 w=4.4e-07
MXN3 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN3_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN3_3 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_3 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_3 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI14_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI14_MXPA1_3 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g0_MXPA1_2 nmsel S0 VDD VNW p12 l=1.3e-07 w=5.6e-07
MXP2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP2_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP2_3 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_3 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2X8MTR Y VDD VNW VPW VSS A B S0
mXI15_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI15_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI15_MXNA1_3 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI15_MXNA1_4 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g0_MXNA1_2 nmsel S0 VSS VPW n12 l=1.3e-07 w=5.8e-07
MXN4 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN4_3 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN4_4 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_3 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_4 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_3 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_4 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI15_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI15_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI15_MXPA1_3 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI15_MXPA1_4 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g0_MXPA1_2 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.1e-07
MXP3 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP3_3 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP3_4 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_4 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_3 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_4 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2XLMTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 Y nmsel nmin0 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=3.6e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=3.6e-07
MXP0 nmin0 S0 Y VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MXI3X1MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=2.9e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=3.2e-07
MXN4 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=3.2e-07
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=3.7e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=3.7e-07
MXN5 net115 net104 net98 VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=3.9e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
MXP1 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=3.9e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=3.9e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=4.6e-07
MXP3 net98 S1 net115 VNW p12 l=1.3e-07 w=4.6e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT MXI3X2MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=4.7e-07
MXN0 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=5.1e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=4.7e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=6.1e-07
MXN1 net115 net104 net98 VPW n12 l=1.3e-07 w=4.1e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t5 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=6.2e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=2.7e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=7.2e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=7.2e-07
MXP0 net98 S1 net115 VNW p12 l=1.3e-07 w=7e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=6e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI3X4MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=4.7e-07
MXN0 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=6.1e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=4.7e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=6.1e-07
MXN1 net115 net104 net98 VPW n12 l=1.3e-07 w=4.1e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t5 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=7.4e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=8.1e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=8.1e-07
MXP0 net98 S1 net115 VNW p12 l=1.3e-07 w=7e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI3X8MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=4.7e-07
MXN0 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=6.1e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=4.7e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=6.1e-07
MXN1 net115 net104 net98 VPW n12 l=1.3e-07 w=4.3e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t5 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=7.4e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=8.2e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=7.1e-07
MXP0 net98 S1 net115 VNW p12 l=1.3e-07 w=7e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI3XLMTR Y VDD VNW VPW VSS A B C S0 S1
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=2.1e-07
MXN3 net115 net104 net98 VPW n12 l=1.3e-07 w=2.1e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=2.5e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=2.5e-07
MXP2 net98 S1 net115 VNW p12 l=1.3e-07 w=2.5e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT MXI4X1MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=3.2e-07
MXN2 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=3.2e-07
MXN1 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=3.2e-07
mXI18_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g4_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=3.2e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=3.2e-07
MXN0 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=3.2e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=3.7e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=3.7e-07
MXN3 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=3.7e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=3.9e-07
MXP2 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=3.9e-07
MXP1 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=3.9e-07
mXI18_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=3.9e-07
mX_g4_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=3.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=3.9e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=3.9e-07
MXP0 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=3.9e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=3.9e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=4.6e-07
MXP3 net112 S1 net99 VNW p12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MXI4X2MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=5.1e-07
MXN2 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=5.1e-07
MXN1 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=4.2e-07
mXI18_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=4.4e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=4e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=4.9e-07
MXN0 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=5.2e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=4.8e-07
MXN3 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=4.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP2 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=6.3e-07
MXP4 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mXI18_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g4_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=5.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=5.7e-07
MXP0 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=6.3e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=7.4e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=7.4e-07
MXP5 net112 S1 net99 VNW p12 l=1.3e-07 w=7.4e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI4X4MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN5 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=6.1e-07
MXN4 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=4e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=6.1e-07
MXN0 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=6.1e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=5e-07
MXN3 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=4.4e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP7 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=7.4e-07
MXP6 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mXI18_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=5.7e-07
MXP0 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=7.4e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=8.4e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=8.4e-07
MXP5 net112 S1 net99 VNW p12 l=1.3e-07 w=8.3e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI4X8MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN5 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=6.1e-07
MXN4 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=4e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=6.1e-07
MXN0 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=6.1e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=5e-07
MXN3 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=4.4e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP7 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=7.4e-07
MXP6 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mXI18_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=5.7e-07
MXP0 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=7.4e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=8.4e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=8.4e-07
MXP5 net112 S1 net99 VNW p12 l=1.3e-07 w=8.3e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI4XLMTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=3e-07
MXN6 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=3e-07
MXN5 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=1.8e-07
mXI21_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=2.1e-07
MXN7 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=2.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=3e-07
MXP6 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=2.3e-07
mXI21_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=3e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=2.5e-07
MXP7 net112 S1 net99 VNW p12 l=1.3e-07 w=2.5e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND2BX12MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_3 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2_2 XI1_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y a XI1_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 XI1_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 XI1_n1__4 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y a XI1_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y a XI1_n1__5 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_5 XI1_n1__5 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_6 XI1_n1__6 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y a XI1_n1__6 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_2 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_3 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2BX1MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND2BX2MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2BX4MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2_2 XI1_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2BX8MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2_2 XI1_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y a XI1_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 XI1_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 XI1_n1__4 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y a XI1_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_2 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2BXLMTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n1__4 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A XI0_n1__5 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 XI0_n1__5 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_6 XI0_n1__6 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A XI0_n1__6 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2X1MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2X3MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT NAND2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2X5MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_3 XI0_n1 B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 Y A XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 Y A XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7.3e-07
.ends


.SUBCKT NAND2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n1__4 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2XLMTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND3BX1MTR Y VDD VNW VPW VSS AN B C
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA3 XI1_n1 C VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA2 XI1_n2 B XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y a XI1_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND3BX2MTR Y VDD VNW VPW VSS AN B C
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA3 XI1_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n2 B XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3BX4MTR Y VDD VNW VPW VSS AN B C
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA3_2 XI1_n1__2 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 XI1_n2__2 B XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n2 B XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA3 XI1_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3BXLMTR Y VDD VNW VPW VSS AN B C
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA3 XI1_n1 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n2 B XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y a XI1_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND3X12MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_5 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_6 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_6 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_4 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_5 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_6 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3X1MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND3X2MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3X3MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y A XI0_n2__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT NAND3X4MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3X6MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n2__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n2__3 B XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n1__3 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3X8MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y A XI0_n2__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_3 Y A XI0_n2__3 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_3 XI0_n2__3 B XI0_n1__3 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3_3 XI0_n1__3 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3_4 XI0_n1__4 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_4 XI0_n2__4 B XI0_n1__4 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_4 Y A XI0_n2__4 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA3_4 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT NAND3XLMTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND4BBX1MTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net43 D VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net47 C net43 VPW n12 l=1.3e-07 w=3.6e-07
MXN0 net51 B net47 VPW n12 l=1.3e-07 w=3.6e-07
MXNA Y A net51 VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 Y D VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP1 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
MXPA Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT NAND4BBX2MTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=3e-07
MXN7 net43 D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN6 net47 C net43 VPW n12 l=1.3e-07 w=7.1e-07
MXN5 net51 B net47 VPW n12 l=1.3e-07 w=7.1e-07
MXNA Y A net51 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP5 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=3.7e-07
.ends


.SUBCKT NAND4BBX4MTR Y VDD VNW VPW VSS AN BN C D
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN11 net43 D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 net43 D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 net47 C net43 VPW n12 l=1.3e-07 w=7.1e-07
MXN10_2 net47 C net43 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net51 B net47 VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 net51 B net47 VPW n12 l=1.3e-07 w=7.1e-07
MXNA Y A net51 VPW n12 l=1.3e-07 w=7.1e-07
MXNA_2 Y A net51 VPW n12 l=1.3e-07 w=7.2e-07
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP5 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A VDD VNW p12 l=1.3e-07 w=8e-07
MXPA_2 Y A VDD VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT NAND4BBXLMTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN12 net43 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net47 C net43 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net51 B net47 VPW n12 l=1.3e-07 w=1.8e-07
MXNA Y A net51 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 Y D VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP9 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP8 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
MXPA Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT NAND4BX1MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA4 XI1_n1 D VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA3 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y a XI1_n3 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND4BX2MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA4 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA3 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4BX4MTR Y VDD VNW VPW VSS AN B C D
mXI1_MXNA4 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA4_2 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA3 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA3_2 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT NAND4BXLMTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA4 XI1_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA3 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y a XI1_n3 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND4X12MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_5 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_6 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_5 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_6 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_6 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_3 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_5 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_6 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_4 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_5 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_6 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4X1MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND4X2MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4X4MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4_2 XI0_n1__2 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2__2 C XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3__2 B XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n3__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4X6MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_3 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4X8MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_3 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_4 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4XLMTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR2BX12MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_3 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_5 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_6 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_2 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_3 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPA2_2 XI1_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y a XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y a XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y a XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y a XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2BX1MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NOR2BX2MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2BX4MTR Y VDD VNW VPW VSS AN B
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPA2_2 XI1_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT NOR2BX8MTR Y VDD VNW VPW VSS AN B
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPA2_2 XI1_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y a XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y a XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_2 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
.ends


.SUBCKT NOR2BXLMTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_6 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 XI0_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A XI0_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 XI0_p1__5 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_6 XI0_p1__6 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A XI0_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2X1MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NOR2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2X3MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT NOR2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2X5MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1_3 Y A XI0_p1__3 VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=7.3e-07
.ends


.SUBCKT NOR2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 XI0_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2XLMTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR3BX1MTR Y VDD VNW VPW VSS AN B C
mX_g0_MXNA1 net38 AN VSS VPW n12 l=1.3e-07 w=1.9e-07
MX_t5 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y net38 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 net38 AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t0 VDD C net33 VNW p12 l=1.3e-07 w=6.2e-07
MXP0 net33 B net30 VNW p12 l=1.3e-07 w=6.2e-07
MXP1 net30 net38 Y VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NOR3BX2MTR Y VDD VNW VPW VSS AN B C
mX_g0_MXNA1 net38 AN VSS VPW n12 l=1.3e-07 w=3e-07
MX_t5 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN3 Y net38 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 net38 AN VDD VNW p12 l=1.3e-07 w=3.7e-07
MX_t0 VDD C net33 VNW p12 l=1.3e-07 w=8.7e-07
MXP2 net33 B net30 VNW p12 l=1.3e-07 w=8.7e-07
MXP3 net30 net38 Y VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3BX4MTR Y VDD VNW VPW VSS AN B C
mX_g0_MXNA1 net38 AN VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t5 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 Y net38 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5_2 Y net38 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MX_t5_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 net38 AN VDD VNW p12 l=1.3e-07 w=7.4e-07
MX_t0_2 VDD C net33__2 VNW p12 l=1.3e-07 w=8.1e-07
MXP4_2 net33__2 B net30__2 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_2 net30__2 net38 Y VNW p12 l=1.3e-07 w=8.1e-07
MXP5 net30 net38 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net33 B net30 VNW p12 l=1.3e-07 w=8.7e-07
MX_t0 VDD C net33 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3BXLMTR Y VDD VNW VPW VSS AN B C
mX_g0_MXNA1 net38 AN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t5 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 Y net38 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXPA1 net38 AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t0 VDD C net33 VNW p12 l=1.3e-07 w=3.6e-07
MXP4 net33 B net30 VNW p12 l=1.3e-07 w=3.6e-07
MXP5 net30 net38 Y VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR3X12MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_5 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA2_6 Y B VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA3_6 Y C VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_2 Y A XI0_p2__2 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_3 Y A XI0_p2__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_3 XI0_p2__3 B XI0_p1__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_3 XI0_p1__3 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_4 XI0_p1__4 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_4 XI0_p2__4 B XI0_p1__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_4 Y A XI0_p2__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_5 Y A XI0_p2__5 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2_5 XI0_p2__5 B XI0_p1__5 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3_5 XI0_p1__5 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_6 XI0_p1__6 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_6 XI0_p2__6 B XI0_p1__6 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_6 Y A XI0_p2__6 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3X1MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NOR3X2MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3X4MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p2__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3X6MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p2__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A XI0_p2__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_3 XI0_p2__3 B XI0_p1__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_3 XI0_p1__3 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.1e-07
.ends


.SUBCKT NOR3X8MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_2 Y A XI0_p2__2 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_3 Y A XI0_p2__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_3 XI0_p2__3 B XI0_p1__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_3 XI0_p1__3 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_4 XI0_p1__4 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_4 XI0_p2__4 B XI0_p1__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_4 Y A XI0_p2__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3XLMTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR4BBX1MTR Y VDD VNW VPW VSS AN BN C D
MXN2 Y D VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=2.5e-07
MXPD net90 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0 net86 C net90 VNW p12 l=1.3e-07 w=8.7e-07
MXP1 net068 B net86 VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y A net068 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=3e-07
.ends


.SUBCKT NOR4BBX2MTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=4.9e-07
MXN5 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=6e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=6e-07
MXP5_2 Y A net068__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_2 net068__2 B net86__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 net86__2 C net90__2 VNW p12 l=1.3e-07 w=8.7e-07
MXPD_2 net90__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPD net90 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP3 net86 C net90 VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net068 B net86 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y A net068 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BBX4MTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_2 A AN VSS VPW n12 l=1.3e-07 w=5e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=5e-07
mXI1_MXNA1_2 B BN VSS VPW n12 l=1.3e-07 w=5e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN9 Y D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN9_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI0_MXPA1_2 A AN VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI1_MXPA1_2 B BN VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP5_2 Y A net068__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_2 net068__2 B net86__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP6_2 net86__2 C net90__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP7_2 net90__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7_3 net90__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6_3 net86__3 C net90__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_3 net068__3 B net86__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_3 Y A net068__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_4 Y A net068__4 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_4 net068__4 B net86__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP6_4 net86__4 C net90__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_4 net90__4 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7 net90 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6 net86 C net90 VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net068 B net86 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y A net068 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BBXLMTR Y VDD VNW VPW VSS AN BN C D
MXN5 Y D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=1.9e-07
MXP5 net90 D VDD VNW p12 l=1.3e-07 w=4.7e-07
MXP4 net86 C net90 VNW p12 l=1.3e-07 w=4.7e-07
MXP3 net068 B net86 VNW p12 l=1.3e-07 w=4.7e-07
MXP2 Y A net068 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT NOR4BX1MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=2.5e-07
MXN2 Y D VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=3e-07
MXPD net33 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0 net29 C net33 VNW p12 l=1.3e-07 w=8.7e-07
MXP1 net25 B net29 VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y A net25 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BX2MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=4.9e-07
MXN5 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=6e-07
MXPA_2 Y A net25__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 net25__2 B net29__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP1_2 net29__2 C net33__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP2_2 net33__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 net33 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP1 net29 C net33 VNW p12 l=1.3e-07 w=8.7e-07
MXP0 net25 B net29 VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A net25 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BX4MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_2 A AN VSS VPW n12 l=1.3e-07 w=5e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=6e-07
MXN6 Y D VSS VPW n12 l=1.3e-07 w=6e-07
MXN6_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI0_MXPA1_2 A AN VDD VNW p12 l=1.3e-07 w=6.1e-07
MXPA_2 Y A net25__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 net25__2 B net29__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_2 net29__2 C net33__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 net33__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5_3 net33__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4_3 net29__3 C net33__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_3 net25__3 B net29__3 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_3 Y A net25__3 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_4 Y A net25__4 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_4 net25__4 B net29__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP4_4 net29__4 C net33__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_4 net33__4 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP5 net33 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net29 C net33 VNW p12 l=1.3e-07 w=8.7e-07
MXP3 net25 B net29 VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A net25 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BXLMTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 Y D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net33 D VDD VNW p12 l=1.3e-07 w=4.7e-07
MXP10 net29 C net33 VNW p12 l=1.3e-07 w=4.7e-07
MXP9 net25 B net29 VNW p12 l=1.3e-07 w=4.7e-07
MXP8 Y A net25 VNW p12 l=1.3e-07 w=4.7e-07
.ends


.SUBCKT NOR4X12MTR Y VDD VNW VPW VSS A B C D
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNC Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNC_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB_2 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_3 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNB_3 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNC_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_3 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_4 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNC_4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB_4 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_4 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_5 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNB_5 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNC_5 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_5 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_6 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNC_6 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB_6 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_3 Y A net37__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_3 net37__3 B net40__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP7_3 net40__3 C net43__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net43__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net43__4 D VDD VNW p12 l=1.3e-07 w=7.8e-07
MXP7_4 net40__4 C net43__4 VNW p12 l=1.3e-07 w=7.8e-07
MXP5_4 net37__4 B net40__4 VNW p12 l=1.3e-07 w=7.8e-07
MXPA_4 Y A net37__4 VNW p12 l=1.3e-07 w=7.8e-07
MXPA_5 Y A net37__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_5 net37__5 B net40__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_5 net40__5 C net43__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_5 net43__5 D VDD VNW p12 l=1.3e-07 w=7.8e-07
MXP8_6 net43__6 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7_6 net40__6 C net43__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_6 net37__6 B net40__6 VNW p12 l=1.3e-07 w=8.1e-07
MXPA_6 Y A net37__6 VNW p12 l=1.3e-07 w=8.1e-07
MXPA_7 Y A net37__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_7 net37__7 B net40__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_7 net40__7 C net43__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_7 net43__7 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP8_8 net43__8 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7_8 net40__8 C net43__8 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_8 net37__8 B net40__8 VNW p12 l=1.3e-07 w=8.1e-07
MXPA_8 Y A net37__8 VNW p12 l=1.3e-07 w=8.1e-07
MXPA_9 Y A net37__9 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_9 net37__9 B net40__9 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_9 net40__9 C net43__9 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_9 net43__9 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP8_10 net43__10 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7_10 net40__10 C net43__10 VNW p12 l=1.3e-07 w=7.8e-07
MXP5_10 net37__10 B net40__10 VNW p12 l=1.3e-07 w=7.8e-07
MXPA_10 Y A net37__10 VNW p12 l=1.3e-07 w=7.8e-07
MXPA_11 Y A net37__11 VNW p12 l=1.3e-07 w=7.8e-07
MXP5_11 net37__11 B net40__11 VNW p12 l=1.3e-07 w=7.8e-07
MXP7_11 net40__11 C net43__11 VNW p12 l=1.3e-07 w=7.8e-07
MXP8_11 net43__11 D VDD VNW p12 l=1.3e-07 w=7.8e-07
MXP8_12 net43__12 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7_12 net40__12 C net43__12 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_12 net37__12 B net40__12 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_12 Y A net37__12 VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP7 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4X1MTR Y VDD VNW VPW VSS A B C D
MXN7 Y D VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN5 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4X2MTR Y VDD VNW VPW VSS A B C D
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP13_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4X4MTR Y VDD VNW VPW VSS A B C D
MXN14 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13 Y B VSS VPW n12 l=1.3e-07 w=6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=6e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_3 Y A net37__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_3 net37__3 B net40__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP12_3 net40__3 C net43__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net43__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net43__4 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_4 net40__4 C net43__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP17_4 net37__4 B net40__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP18_4 Y A net37__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP18 Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
MXP17 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4X6MTR Y VDD VNW VPW VSS A B C D
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_3 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_3 Y A net37__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_3 net37__3 B net40__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP12_3 net40__3 C net43__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net43__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net43__4 D VDD VNW p12 l=1.3e-07 w=7.8e-07
MXP12_4 net40__4 C net43__4 VNW p12 l=1.3e-07 w=7.8e-07
MXP17_4 net37__4 B net40__4 VNW p12 l=1.3e-07 w=7.8e-07
MXP18_4 Y A net37__4 VNW p12 l=1.3e-07 w=7.8e-07
MXP18_5 Y A net37__5 VNW p12 l=1.3e-07 w=8.2e-07
MXP17_5 net37__5 B net40__5 VNW p12 l=1.3e-07 w=8.2e-07
MXP12_5 net40__5 C net43__5 VNW p12 l=1.3e-07 w=8.2e-07
MXP8_5 net43__5 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_6 net43__6 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_6 net40__6 C net43__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP17_6 net37__6 B net40__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP18_6 Y A net37__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP18 Y A net37 VNW p12 l=1.3e-07 w=8.1e-07
MXP17 net37 B net40 VNW p12 l=1.3e-07 w=8.1e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=8.1e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.1e-07
.ends


.SUBCKT NOR4X8MTR Y VDD VNW VPW VSS A B C D
MXN14 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B VSS VPW n12 l=1.3e-07 w=6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=6e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXN9_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_3 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_3 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA_4 Y A VSS VPW n12 l=1.3e-07 w=6e-07
MXN11_4 Y B VSS VPW n12 l=1.3e-07 w=6e-07
MXN9_4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_4 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_3 Y A net37__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_3 net37__3 B net40__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP12_3 net40__3 C net43__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net43__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net43__4 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_4 net40__4 C net43__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP19_4 net37__4 B net40__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP20_4 Y A net37__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP20_5 Y A net37__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP19_5 net37__5 B net40__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP12_5 net40__5 C net43__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_5 net43__5 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_6 net43__6 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_6 net40__6 C net43__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP19_6 net37__6 B net40__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP20_6 Y A net37__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP20_7 Y A net37__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP19_7 net37__7 B net40__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP12_7 net40__7 C net43__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_7 net43__7 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_8 net43__8 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_8 net40__8 C net43__8 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_8 net37__8 B net40__8 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_8 Y A net37__8 VNW p12 l=1.3e-07 w=8.7e-07
MXP20 Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
MXP19 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4XLMTR Y VDD VNW VPW VSS A B C D
MXN10 Y D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=4.7e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=4.7e-07
MXP13 net37 B net40 VNW p12 l=1.3e-07 w=4.7e-07
MXP14 Y A net37 VNW p12 l=1.3e-07 w=4.7e-07
.ends


.SUBCKT OA21X1MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OA21X2MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA21X4MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA21X8MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPB1_2 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 ny B0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA21XLMTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OA22X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 ny A1 net48 VPW n12 l=1.3e-07 w=2.3e-07
MXN3 ny A0 net48 VPW n12 l=1.3e-07 w=2.3e-07
MXN4 net48 B0 VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN5 net48 B1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP6 net67 A1 VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP5 ny A0 net67 VNW p12 l=1.3e-07 w=3.1e-07
MXP4 ny B0 net73 VNW p12 l=1.3e-07 w=3.1e-07
MXP8 net73 B1 VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OA22X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 ny A1 net45 VPW n12 l=1.3e-07 w=3.6e-07
MXN7 ny A0 net45 VPW n12 l=1.3e-07 w=3.6e-07
MXN8 net45 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN9 net45 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP7 net60 A1 VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP9 ny A0 net60 VNW p12 l=1.3e-07 w=5.1e-07
MXP10 ny B0 net66 VNW p12 l=1.3e-07 w=5.1e-07
MXP8 net66 B1 VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA22X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 ny A1 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN10 ny A0 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 net45 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net45 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP11 net60 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12 ny A0 net60 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 ny B0 net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net66 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA22X8MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN13 ny A0 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 ny A1 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 ny A1 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 ny A0 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN14 net45 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15 net45 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 net45 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 net45 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP15_2 ny A0 net60__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14_2 net60__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP14 net60 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 ny A0 net60 VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 ny B0 net66__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net66__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net66 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16 ny B0 net66 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA22XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 ny A1 net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 ny A0 net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net45 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net45 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP7 net60 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 ny A0 net60 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 ny B0 net66 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net66 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI211X1MTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI211X2MTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI211X4MTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n2__2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPC1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPB1_2 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI211X8MTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC1_3 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2_3 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2_4 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC1_4 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n2__2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 XI0_n2__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 XI0_n2__3 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_4 XI0_n2__4 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y B0 XI0_n2__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPC1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2_3 XI0_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC1_3 Y A0 XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC1_4 Y A0 XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2_4 XI0_p1__4 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPB1_2 Y C0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPB1_3 Y C0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_3 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_4 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPB1_4 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI211XLMTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI21BX1MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT OAI21BX2MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=3.7e-07
.ends


.SUBCKT OAI21BX4MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPB2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT OAI21BX8MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_3 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_3 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_4 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_4 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXPB2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_3 Y A0 XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_3 XI1_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_4 XI1_p1__4 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_4 Y A0 XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21BXLMTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT OAI21X1MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI21X2MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21X3MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPB2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT OAI21X4MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21X6MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_3 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_3 Y A0 XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_3 XI0_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21X8MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_3 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_4 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_4 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_3 Y A0 XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_3 XI0_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_4 XI0_p1__4 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_4 Y A0 XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21XLMTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI221X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN2 net33 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net33 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 net25 A1 net33 VPW n12 l=1.3e-07 w=3.6e-07
MXN1 net25 A0 net33 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y C0 net25 VPW n12 l=1.3e-07 w=3.6e-07
MXP0 Y B0 net46 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 net46 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP2 net58 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP1 Y A0 net58 VNW p12 l=1.3e-07 w=6.2e-07
MXP3 Y C0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI221X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN7 net33 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 net33 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 net25 A1 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN8 net25 A0 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 net25 VPW n12 l=1.3e-07 w=7.1e-07
MXP5 Y B0 net073 VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net073 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6 net059 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7 Y A0 net059 VNW p12 l=1.3e-07 w=8.7e-07
MXP3 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI221X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN11 net33 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 net33 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10_2 net33 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 net33 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net25 A0 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net25 A1 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 net25 A1 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN12_2 net25 A0 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 net25 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y C0 net25 VPW n12 l=1.3e-07 w=7.1e-07
MXP9_2 Y B0 net077__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net077__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net077 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y B0 net077 VNW p12 l=1.3e-07 w=8.7e-07
MXP11_2 Y A0 net069__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP10_2 net069__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net069 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP11 Y A0 net069 VNW p12 l=1.3e-07 w=8.7e-07
MXP3 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI221XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN10 net33 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net33 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net25 A1 net33 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net25 A0 net33 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 Y C0 net25 VPW n12 l=1.3e-07 w=1.8e-07
MXP5 Y B0 net069 VNW p12 l=1.3e-07 w=3.6e-07
MXP4 net069 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP7 net077 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP6 Y A0 net077 VNW p12 l=1.3e-07 w=3.6e-07
MXP3 Y C0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI222X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN2 net28 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 net28 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 net24 A1 net28 VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net24 A0 net28 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y C0 net24 VPW n12 l=1.3e-07 w=3.6e-07
MXN4 Y C1 net24 VPW n12 l=1.3e-07 w=3.6e-07
MXP6 Y B0 net089 VNW p12 l=1.3e-07 w=6.2e-07
MXP5 net089 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP9 net083 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP10 Y A0 net083 VNW p12 l=1.3e-07 w=6.2e-07
MXP7 Y C0 net59 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 net59 C1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI222X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN8 net28 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 net28 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net24 A1 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN7 net24 A0 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXN5 Y C1 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXP12 Y B0 net094 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 net094 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP14 net088 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 Y A0 net088 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 Y C0 net59 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net59 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI222X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN13 net28 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15 net28 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 net28 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 net28 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net24 A0 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN14 net24 A1 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 net24 A1 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN12_2 net24 A0 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y C1 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y C1 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y C0 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXP19_2 Y B0 net082__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 net082__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16 net082 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP19 Y B0 net082 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A0 net092__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net092__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17 net092 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP18 Y A0 net092 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 Y C0 net59__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net59__2 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net59 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP20 Y C0 net59 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI222XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN2 net28 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net28 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net24 A1 net28 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net24 A0 net28 VPW n12 l=1.3e-07 w=3e-07
MXN6 Y C0 net24 VPW n12 l=1.3e-07 w=3e-07
MXN4 Y C1 net24 VPW n12 l=1.3e-07 w=3e-07
MXP14 Y B0 net082 VNW p12 l=1.3e-07 w=3.6e-07
MXP11 net082 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP12 net086 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP13 Y A0 net086 VNW p12 l=1.3e-07 w=3.6e-07
MXP15 Y C0 net59 VNW p12 l=1.3e-07 w=3.6e-07
MXP8 net59 C1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI22X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y A0 net072 VPW n12 l=1.3e-07 w=3.6e-07
MXN1 net072 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN2 net072 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP0 net22 A1 VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP1 Y A0 net22 VNW p12 l=1.3e-07 w=5.9e-07
MXP2 Y B0 net32 VNW p12 l=1.3e-07 w=5.9e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=5.9e-07
.ends


.SUBCKT OAI22X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN3 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN4 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP3 net22 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 Y A0 net22 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y B0 net32 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI22X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN3 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN3_2 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN4 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5_2 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4_2 Y A0 net22__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 net22__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP3 net22 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 Y A0 net22 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 Y B0 net32__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net32__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y B0 net32 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI22X8MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN8 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_2 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_3 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_3 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_4 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_4 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN7_2 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN7_3 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_3 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_4 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN7_4 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXP9_2 Y B0 net32__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net32__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net32__3 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9_3 Y B0 net32__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP9_4 Y B0 net32__4 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net32__4 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y B0 net32 VNW p12 l=1.3e-07 w=8.7e-07
MXP7_2 Y A0 net22__2 VNW p12 l=1.3e-07 w=8.1e-07
MXP6_2 net22__2 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP6_3 net22__3 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7_3 Y A0 net22__3 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_4 Y A0 net22__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP6_4 net22__4 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP6 net22 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7 Y A0 net22 VNW p12 l=1.3e-07 w=8.1e-07
.ends


.SUBCKT OAI22XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 Y A0 net072 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net072 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net072 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP3 net22 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP4 Y A0 net22 VNW p12 l=1.3e-07 w=3.6e-07
MXP5 Y B0 net32 VNW p12 l=1.3e-07 w=3.6e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2B11X1MTR Y VDD VNW VPW VSS A0 A1N B0 C0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNC2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNC1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y B0 XI1_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB1 XI1_n2 C0 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPC2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPC1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2B11X2MTR Y VDD VNW VPW VSS A0 A1N B0 C0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNC2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNC1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n2 C0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPC2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPC1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B11X4MTR Y VDD VNW VPW VSS A0 A1N B0 C0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNC2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNC1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNC1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNC2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n2__2 C0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y B0 XI1_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n2 C0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPC2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPC1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPC1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPC2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B11XLMTR Y VDD VNW VPW VSS A0 A1N B0 C0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNC2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNC1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y B0 XI1_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n2 C0 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPC2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPC1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2B1X1MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2B1X2MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B1X4MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPB2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B1X8MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_3 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_3 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_4 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_4 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPB2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_3 Y A0 XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_3 XI1_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_4 XI1_p1__4 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_4 Y A0 XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B1XLMTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2B2X1MTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2B2X2MTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B2X4MTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2_2 XI1_p1A__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y A0 XI1_p1A__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_2 XI1_p1B__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y B0 XI1_p1B__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B2X8MTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_3 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_3 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_4 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_4 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2_2 XI1_p1A__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y A0 XI1_p1A__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y A0 XI1_p1A__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI1_MXPA2_3 XI1_p1A__3 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI1_MXPA2_4 XI1_p1A__4 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI1_MXPA1_4 Y A0 XI1_p1A__4 VNW p12 l=1.3e-07 w=8.1e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_2 XI1_p1B__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y B0 XI1_p1B__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_3 Y B0 XI1_p1B__3 VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPB2_3 XI1_p1B__3 B1 VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPB2_4 XI1_p1B__4 B1 VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPB1_4 Y B0 XI1_p1B__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B2XLMTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2BB1X1MTR Y VDD VNW VPW VSS A0N A1N B0
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2BB1X2MTR Y VDD VNW VPW VSS A0N A1N B0
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI1_MXPA2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB1X4MTR Y VDD VNW VPW VSS A0N A1N B0
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPA2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB1XLMTR Y VDD VNW VPW VSS A0N A1N B0
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2BB2X1MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2BB2X2MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB2X4MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_2 XI1_p1__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y B0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB2X8MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA1_2 nmin1 A1N XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1__2 A0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_3 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_3 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_4 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_4 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA2_2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 nmin1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_2 XI1_p1__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y B0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_3 Y B0 XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_3 XI1_p1__3 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_4 XI1_p1__4 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_4 Y B0 XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB2XLMTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=3e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI31X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0
MXN3 n1 A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN2 n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXPA2 net42 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP1 net039 A1 net42 VNW p12 l=1.3e-07 w=6.2e-07
MXP2 Y A0 net039 VNW p12 l=1.3e-07 w=6.2e-07
MXP3 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI31X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0
MXN6 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXPA2 net42 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net039 A1 net42 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y A0 net039 VNW p12 l=1.3e-07 w=8.7e-07
MXP6 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI31X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0
MXN9 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7_2 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_2 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXNB0_2 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXPA2_2 net42__2 A2 VDD VNW p12 l=1.3e-07 w=8.2e-07
MXP10_2 net039__2 A1 net42__2 VNW p12 l=1.3e-07 w=8.2e-07
MXP11_2 Y A0 net039__2 VNW p12 l=1.3e-07 w=8.2e-07
MXP11 Y A0 net039 VNW p12 l=1.3e-07 w=8.2e-07
MXP10 net039 A1 net42 VNW p12 l=1.3e-07 w=8.2e-07
MXPA2 net42 A2 VDD VNW p12 l=1.3e-07 w=8.2e-07
MXP9 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI31XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0
MXN6 n1 A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXPA2 net42 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP4 net039 A1 net42 VNW p12 l=1.3e-07 w=3.6e-07
MXP5 Y A0 net039 VNW p12 l=1.3e-07 w=3.6e-07
MXP6 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI32X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
MXN3 n1 A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN4 n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN5 n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y B0 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXN2 Y B1 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXP1 net59 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP4 net67 A1 net59 VNW p12 l=1.3e-07 w=6.2e-07
MXP5 Y A0 net67 VNW p12 l=1.3e-07 w=6.2e-07
MXP3 Y B0 net55 VNW p12 l=1.3e-07 w=6.2e-07
MXP2 net55 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI32X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
MXN7 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y B1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXPA2 net59 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net67 A1 net59 VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y A0 net67 VNW p12 l=1.3e-07 w=8.7e-07
MXP7 Y B0 net55 VNW p12 l=1.3e-07 w=8.7e-07
MXP6 net55 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI32X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
MXN12 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12_2 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN10 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN10_2 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y B1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXP10_2 net59__2 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP13_2 net67__2 A1 net59__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14_2 Y A0 net67__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 Y A0 net67 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 net67 A1 net59 VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net59 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP11_2 net55__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 Y B0 net55__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 Y B0 net55 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 net55 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI32XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
MXN16 n1 A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN17 n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN18 n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 Y B1 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXPA2 net59 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP17 net67 A1 net59 VNW p12 l=1.3e-07 w=3.6e-07
MXP18 Y A0 net67 VNW p12 l=1.3e-07 w=3.6e-07
MXP16 Y B0 net55 VNW p12 l=1.3e-07 w=3.6e-07
MXP15 net55 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI33X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN4 VSS B2 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXN5 VSS B1 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 VSS B0 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXN2 n1 A0 Y VPW n12 l=1.3e-07 w=3.6e-07
MXN1 n1 A1 Y VPW n12 l=1.3e-07 w=3.6e-07
MXN3 n1 A2 Y VPW n12 l=1.3e-07 w=3.6e-07
MXP1 net77 B2 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 net73 B1 net77 VNW p12 l=1.3e-07 w=6.2e-07
MXP4 Y B0 net73 VNW p12 l=1.3e-07 w=6.2e-07
MXP6 Y A0 net89 VNW p12 l=1.3e-07 w=6.2e-07
MXP5 net89 A1 net81 VNW p12 l=1.3e-07 w=6.2e-07
MXP2 net81 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI33X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN10 n1 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 Y A0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y A1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN8 Y A2 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXP7 net77 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 net73 B1 net77 VNW p12 l=1.3e-07 w=8.7e-07
MXP10 Y B0 net73 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 Y A0 net89 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 net89 A1 net81 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net81 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI33X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN16 n1 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN17 n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN18 n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN18_2 n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN17_2 n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN16_2 n1 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15 Y A2 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN13 Y A1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN14 Y A0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 Y A0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 Y A1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 Y A2 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXP14_2 net77__2 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15_2 net73__2 B1 net77__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 Y B0 net73__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP16 Y B0 net73 VNW p12 l=1.3e-07 w=8.7e-07
MXP15 net73 B1 net77 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 net77 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP13_2 net81__2 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net89__2 A1 net81__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A0 net89__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18 Y A0 net89 VNW p12 l=1.3e-07 w=8.1e-07
MXP17 net89 A1 net81 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 net81 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI33XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN9 n1 B2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 n1 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 n1 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN18 Y A0 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 Y A1 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 Y A2 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXP7 net77 B2 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP8 net73 B1 net77 VNW p12 l=1.3e-07 w=3.6e-07
MXP9 Y B0 net73 VNW p12 l=1.3e-07 w=3.6e-07
MXP11 Y A0 net89 VNW p12 l=1.3e-07 w=3.6e-07
MXP10 net89 A1 net81 VNW p12 l=1.3e-07 w=3.6e-07
MXPA2 net81 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OR2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 XI0_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 ny A XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR2X1MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OR2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X12MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2_3 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3_2 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3_3 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_4 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_5 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X1MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=4.8e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=4.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OR3X2MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X4MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_2 ny A XI0_p2__2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X6MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_2 ny A XI0_p2__2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X8MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3_2 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X12MTR Y VDD VNW VPW VSS A B C D
MXN14 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN14_2 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN14_3 net43 D VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN14_4 net43 D VSS VPW n12 l=1.3e-07 w=3e-07
MXN13 net43 C VSS VPW n12 l=1.3e-07 w=3e-07
MXN13_2 net43 C VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN13_3 net43 C VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN13_4 net43 C VSS VPW n12 l=1.3e-07 w=3e-07
MXN13_5 net43 C VSS VPW n12 l=1.3e-07 w=3e-07
MXN13_6 net43 C VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN12 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN12_2 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN12_3 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA_2 net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA_3 net43 A VSS VPW n12 l=1.3e-07 w=3.1e-07
MXNA_4 net43 A VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI0_MXNA1_2 Y net43 VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI0_MXNA1_3 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 net62 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_3 net62 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_4 net62 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_5 net62 D VDD VNW p12 l=1.3e-07 w=1.23e-06
MXP20 net66 C net62 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 net66 C net62 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_3 net66 C net62 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_4 net66 C net62 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_5 net66 C net62 VNW p12 l=1.3e-07 w=1.23e-06
MXP21 net70 B net66 VNW p12 l=1.3e-07 w=1.23e-06
MXP21_2 net70 B net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP21_3 net70 B net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP21_4 net70 B net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP21_5 net70 B net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP22 net43 A net70 VNW p12 l=1.3e-07 w=8.7e-07
MXP22_2 net43 A net70 VNW p12 l=1.3e-07 w=8.7e-07
MXP22_3 net43 A net70 VNW p12 l=1.3e-07 w=8.7e-07
MXP22_4 net43 A net70 VNW p12 l=1.3e-07 w=8.7e-07
MXP22_5 net43 A net70 VNW p12 l=1.3e-07 w=1.23e-06
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X1MTR Y VDD VNW VPW VSS A B C D
MXNA net43 A VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN0 net43 B VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN1 net43 C VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN2 net43 D VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP7 net43 A net70 VNW p12 l=1.3e-07 w=4.9e-07
MXP6 net70 B net66 VNW p12 l=1.3e-07 w=4.9e-07
MXP5 net66 C net62 VNW p12 l=1.3e-07 w=4.9e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OR4X2MTR Y VDD VNW VPW VSS A B C D
MXNA net43 A VSS VPW n12 l=1.3e-07 w=3e-07
MXN3 net43 B VSS VPW n12 l=1.3e-07 w=3e-07
MXN4 net43 C VSS VPW n12 l=1.3e-07 w=3e-07
MXN5 net43 D VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP10 net43 A net70 VNW p12 l=1.3e-07 w=7.9e-07
MXP9 net70 B net66 VNW p12 l=1.3e-07 w=7.9e-07
MXP8 net66 C net62 VNW p12 l=1.3e-07 w=7.9e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X4MTR Y VDD VNW VPW VSS A B C D
MXN8 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN7 net43 C VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN6 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_2 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP11 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP11_2 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP12 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP12_2 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP13 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP13_2 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X6MTR Y VDD VNW VPW VSS A B C D
MXNA net43 A VSS VPW n12 l=1.3e-07 w=4.6e-07
MXNA_2 net43 A VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN9 net43 B VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN9_2 net43 B VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN10 net43 C VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN10_2 net43 C VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN11 net43 D VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN11_2 net43 D VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP16 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP16_2 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP16_3 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP15 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP15_2 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP15_3 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP14 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP14_2 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP14_3 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_2 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_3 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X8MTR Y VDD VNW VPW VSS A B C D
MXN14 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN14_2 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN13 net43 C VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN13_2 net43 C VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN12 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN12_2 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA_2 net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_2 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_3 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_4 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP17 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP17_2 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP17_3 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP17_4 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP18 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP18_2 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP18_3 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP18_4 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP19 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP19_2 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP19_3 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP19_4 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFHQNX1MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net71 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net48 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 pm nmsi net60 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFHQNX2MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net71 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net48 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.6e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 pm nmsi net60 VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT SDFFHQNX4MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=2.9e-07
MXN2 net71 cn VSS VPW n12 l=1.3e-07 w=2.9e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.2e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=5e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net48 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP3 pm nmsi net60 VNW p12 l=1.3e-07 w=3.5e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=6.1e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFHQNX8MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=3.4e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3e-07
MXN3 net71 cn VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=5.4e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g2_MXNA1_2 s bm VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=4.2e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.8e-07
MXP4 net48 c cn VNW p12 l=1.3e-07 w=4.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.3e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=6.5e-07
MXP5 pm nmsi net60 VNW p12 l=1.3e-07 w=6.5e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.5e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=6e-07
mX_g2_MXPA1_2 s bm VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFHQX1MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.1e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=3.3e-07
MXN1 net54 cn VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.7e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net065 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.6e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=4e-07
MXP2 pm nmsi net71 VNW p12 l=1.3e-07 w=4e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.3e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
.ends


.SUBCKT SDFFHQX2MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=1.9e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=3.1e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=4.8e-07
MXN2 net54 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP3 net065 c cn VNW p12 l=1.3e-07 w=4.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP4 pm nmsi net71 VNW p12 l=1.3e-07 w=5.9e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
.ends


.SUBCKT SDFFHQX4MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=3.2e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.5e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.4e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=6.9e-07
MXN3 net54 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP5 net065 c cn VNW p12 l=1.3e-07 w=7.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=6.7e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP6 pm nmsi net71 VNW p12 l=1.3e-07 w=8e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT SDFFHQX8MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=5.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.5e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.4e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=6.9e-07
MXN3 net54 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.9e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP5 net065 c cn VNW p12 l=1.3e-07 w=7.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=6.7e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=5e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=8.3e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP6 pm nmsi net71 VNW p12 l=1.3e-07 w=8e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT SDFFHX1MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.3e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net0107 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 net104 cn VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 net079 c cn VNW p12 l=1.3e-07 w=4.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.8e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.8e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 nmsi SI net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP10 pm nmsi net087 VNW p12 l=1.3e-07 w=4.4e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.9e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFHX2MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=3.2e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net0107 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=5.1e-07
MXN7 net104 cn VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP13 net079 c cn VNW p12 l=1.3e-07 w=4.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.9e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 nmsi SI net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP12 pm nmsi net087 VNW p12 l=1.3e-07 w=6.2e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g6_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.1e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT SDFFHX4MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.4e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=2.9e-07
MXN8 net0107 SE VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=7e-07
MXN9 net104 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 net079 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=7e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP14 nmsi SI net76 VNW p12 l=1.3e-07 w=3.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 pm nmsi net087 VNW p12 l=1.3e-07 w=8.7e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g6_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT SDFFHX8MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.4e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=2.9e-07
MXN8 net0107 SE VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=7e-07
MXN9 net104 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 net079 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=7e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP14 nmsi SI net76 VNW p12 l=1.3e-07 w=3.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 pm nmsi net087 VNW p12 l=1.3e-07 w=8.7e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g6_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT SDFFNHX1MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmsi SI n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 n1 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=4.3e-07
MXN5 net58 cn VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=4e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP2 net87 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP8 p1 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmsi SI p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=6.8e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP10 pm nmsi net93 VNW p12 l=1.3e-07 w=3.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=4.8e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFNHX2MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmsi SI n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 n1 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=6.1e-07
MXN1 net58 cn VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP2 net87 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP8 p1 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmsi SI p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=8.4e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP5 pm nmsi net93 VNW p12 l=1.3e-07 w=4.6e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFNHX4MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.7e-07
MXN5 nmsi SI net058 VPW n12 l=1.3e-07 w=2.7e-07
MXN7 net058 SE VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=4.6e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=5.4e-07
MXN1 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MX_t3_2 pm nmsi net58 VPW n12 l=1.3e-07 w=5.4e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI59_MXNOE_2 nm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP10 net87 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.3e-07
MXP14 p1 nmse VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP9 nmsi SI p1 VNW p12 l=1.3e-07 w=3.3e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g10_MXPA1_2 cn net185 VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP13 pm nmsi net93 VNW p12 l=1.3e-07 w=6.9e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN_2 nm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g1_MXPA1_3 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFNHX8MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=4.7e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.1e-07
MXN7 nmsi SI n1 VPW n12 l=1.3e-07 w=5.1e-07
MXN6 n1 SE VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=5e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=7.4e-07
MXN1 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MX_t3_2 pm nmsi net58 VPW n12 l=1.3e-07 w=7.4e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI59_MXNOE_2 nm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP14 net87 cn c VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.5e-07
MXP8 p1 nmse VDD VNW p12 l=1.3e-07 w=3.4e-07
MXP15 nmsi SI p1 VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=7.2e-07
mX_g10_MXPA1_2 cn net185 VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP13 pm nmsi net93 VNW p12 l=1.3e-07 w=6.9e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.7e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN_2 nm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFNSRHX1MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net0207 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net0207 VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MX_t30 nmsi SI net172 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 net172 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS SN net163 VPW n12 l=1.3e-07 w=4.3e-07
MXN17 net163 cn net160 VPW n12 l=1.3e-07 w=4.3e-07
MX_t26 pm nmsi net160 VPW n12 l=1.3e-07 w=4.3e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 net0106 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t12 net0106 pm net166 VPW n12 l=1.3e-07 w=4.5e-07
MXN19 VSS RN net166 VPW n12 l=1.3e-07 w=4.5e-07
MXN20 net0106 nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE bm c net0106 VPW n12 l=1.3e-07 w=4e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net181 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net181 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 net0207 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net080 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net080 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn net0207 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP16 nmsi SI net117 VNW p12 l=1.3e-07 w=2.3e-07
MX_t32 net117 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP17 pm nmsi net0125 VNW p12 l=1.3e-07 w=3.3e-07
MX_t24 net0125 c VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI23_MXPA1 XI23_p1 net0106 VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 net0106 pm VDD VNW p12 l=1.3e-07 w=4.8e-07
MXP18 net111 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net0106 RN net111 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net0106 VNW p12 l=1.3e-07 w=4.8e-07
MXP21 bm nmset net126 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 net126 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP24 bm c net132 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net132 nmset net135 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net135 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT SDFFNSRHX2MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net261 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net261 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MX_t30 nmsi SI net168 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 net168 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN26 VSS SN net149 VPW n12 l=1.3e-07 w=6.1e-07
MXN25 net149 cn net153 VPW n12 l=1.3e-07 w=6.1e-07
MX_t26 pm nmsi net153 VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 net129 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN27 net129 pm net145 VPW n12 l=1.3e-07 w=6.3e-07
MXN28 VSS RN net145 VPW n12 l=1.3e-07 w=6.3e-07
MXN20 net129 nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE bm c net129 VPW n12 l=1.3e-07 w=5.5e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net261 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net109 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net109 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn net261 VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP16 nmsi SI net91 VNW p12 l=1.3e-07 w=2.3e-07
MX_t32 net91 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP25 pm nmsi net83 VNW p12 l=1.3e-07 w=4.6e-07
MX_t24 net83 c VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI23_MXPA1 XI23_p1 net129 VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 net129 pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP18 net103 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net129 RN net103 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net129 VNW p12 l=1.3e-07 w=6.7e-07
MXP28 bm nmset net79 VNW p12 l=1.3e-07 w=2.8e-07
MXP20 net79 RN VDD VNW p12 l=1.3e-07 w=2.8e-07
MXP24 bm c net123 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net123 nmset net119 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net119 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFNSRHX4MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net261 CKN VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net261 VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.7e-07
MX_t30 nmsi SI net168 VPW n12 l=1.3e-07 w=2.7e-07
MXN29 net168 SE VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN31 VSS SN net149 VPW n12 l=1.3e-07 w=7.6e-07
MXN30 net149 cn net153 VPW n12 l=1.3e-07 w=7.6e-07
MX_t26 pm nmsi net153 VPW n12 l=1.3e-07 w=7.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 net129 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN27 net129 pm net145 VPW n12 l=1.3e-07 w=8.4e-07
MXN32 VSS RN net145 VPW n12 l=1.3e-07 w=8.4e-07
MXN20 net129 nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI74_MXNOE bm c net129 VPW n12 l=1.3e-07 w=5.5e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net261 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net109 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP29 net109 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 cn net261 VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.2e-07
MXP30 nmsi SI net91 VNW p12 l=1.3e-07 w=3.3e-07
MX_t32 net91 nmse VDD VNW p12 l=1.3e-07 w=3.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP31 pm nmsi net83 VNW p12 l=1.3e-07 w=6.9e-07
MX_t24 net83 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI23_MXPA1 XI23_p1 net129 VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t10_2 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP18 net103 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net129 RN net103 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net129 VNW p12 l=1.3e-07 w=6.7e-07
MXP32 bm nmset net79 VNW p12 l=1.3e-07 w=3.6e-07
MXP20 net79 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP24 bm c net123 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net123 nmset net119 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net119 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFNSRHX8MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net261 CKN VSS VPW n12 l=1.3e-07 w=4.7e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net261 VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g10_MXNA1_2 cn net261 VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.4e-07
MX_t30 nmsi SI net168 VPW n12 l=1.3e-07 w=5.1e-07
MXN33 net168 SE VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN31 VSS SN net149 VPW n12 l=1.3e-07 w=7.6e-07
MXN30 net149 cn net153 VPW n12 l=1.3e-07 w=7.6e-07
MX_t26 pm nmsi net153 VPW n12 l=1.3e-07 w=7.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI23_MXNA1 XI23_n1 net129 VSS VPW n12 l=1.3e-07 w=2.5e-07
MXN27 net129 pm net145 VPW n12 l=1.3e-07 w=8.7e-07
MXN34 VSS RN net145 VPW n12 l=1.3e-07 w=8.7e-07
MXN20 net129 nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI74_MXNOE bm c net129 VPW n12 l=1.3e-07 w=5.5e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=3e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net261 CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MX_t4 net109 CKN VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP33 net109 cn c VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 cn net261 VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g10_MXPA1_2 cn net261 VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=1.03e-06
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=5.8e-07
MXP34 nmsi SI net91 VNW p12 l=1.3e-07 w=5.6e-07
MX_t32 net91 nmse VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=3.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP31 pm nmsi net83 VNW p12 l=1.3e-07 w=6.9e-07
MX_t24 net83 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI23_MXPA1 XI23_p1 net129 VDD VNW p12 l=1.3e-07 w=3.1e-07
MX_t10 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t10_2 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP18 net103 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net129 RN net103 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net129 VNW p12 l=1.3e-07 w=6.7e-07
MXP35 bm nmset net79 VNW p12 l=1.3e-07 w=3.5e-07
MXP20 net79 RN VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP24 bm c net123 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net123 nmset net119 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net119 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQNX1MTR QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net108 SE net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 VSS SI net108 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net111 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net129 D net111 VPW n12 l=1.3e-07 w=1.8e-07
MX_t1 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE pm c XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.7e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net69 nmse net65 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net65 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net68 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net69 D net68 VNW p12 l=1.3e-07 w=3.8e-07
MXP5 pm c net69 VNW p12 l=1.3e-07 w=3.8e-07
mXI1_MXPOEN pm cn XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFQNX2MTR QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net108 SE net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 VSS SI net108 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net111 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net129 D net111 VPW n12 l=1.3e-07 w=1.8e-07
MX_t1 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE pm c XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.7e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP6 net69 nmse net65 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net65 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net68 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net69 D net68 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 pm c net69 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN pm cn XI1_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQNX4MTR QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net108 SE net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 VSS SI net108 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net111 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net129 D net111 VPW n12 l=1.3e-07 w=1.8e-07
MX_t1 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE pm c XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.7e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP6 net69 nmse net65 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net65 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net68 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net69 D net68 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 pm c net69 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN pm cn XI1_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQX1MTR Q VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net064 SE net055 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 VSS SI net064 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net059 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net055 D net059 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm cn net055 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE pm c XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net105 m VSS VPW n12 l=1.3e-07 w=2.8e-07
MX_t12 ns c net105 VPW n12 l=1.3e-07 w=2.8e-07
mXI15_MXNOE ns cn XI15_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI15_MXNA1 XI15_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net076 nmse net070 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net070 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net074 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net076 D net074 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 pm c net076 VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN pm cn XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MX_t14 net80 m VDD VNW p12 l=1.3e-07 w=3.4e-07
MXP7 ns cn net80 VNW p12 l=1.3e-07 w=3.4e-07
mXI15_MXPOEN ns c XI15_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI15_MXPA1 XI15_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFQX2MTR Q VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net064 SE net055 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 VSS SI net064 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net059 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net055 D net059 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm cn net055 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE pm c XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net105 m VSS VPW n12 l=1.3e-07 w=3.9e-07
MX_t12 ns c net105 VPW n12 l=1.3e-07 w=3.9e-07
mXI15_MXNOE ns cn XI15_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI15_MXNA1 XI15_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net076 nmse net070 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net070 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net074 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net076 D net074 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 pm c net076 VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN pm cn XI16_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI16_MXPA1 XI16_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=4.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MX_t14 net80 m VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP8 ns cn net80 VNW p12 l=1.3e-07 w=4.9e-07
mXI15_MXPOEN ns c XI15_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI15_MXPA1 XI15_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQX4MTR Q VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net064 SE net055 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 VSS SI net064 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net059 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net055 D net059 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm cn net055 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE pm c XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net105 m VSS VPW n12 l=1.3e-07 w=4.4e-07
MX_t12 ns c net105 VPW n12 l=1.3e-07 w=4.4e-07
mXI15_MXNOE ns cn XI15_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI15_MXNA1 XI15_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net076 nmse net070 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net070 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net074 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net076 D net074 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 pm c net076 VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN pm cn XI16_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI16_MXPA1 XI16_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MX_t14 net80 m VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP9 ns cn net80 VNW p12 l=1.3e-07 w=6.4e-07
mXI15_MXPOEN ns c XI15_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI15_MXPA1 XI15_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRHQX1MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=3.5e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=3.5e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS RN net128 VPW n12 l=1.3e-07 w=4.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=4.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.7e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP8 net065 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=2.7e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP13 pm nmsi p1 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=6.6e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.3e-07
MX_t15 bm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 bm c net109 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=2.3e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFRHQX2MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS RN net128 VPW n12 l=1.3e-07 w=5.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=5.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP14 net065 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.9e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 pm nmsi p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
MX_t10_2 m pm VDD VNW p12 l=1.3e-07 w=5.1e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 bm RN VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP16 bm c net109 VNW p12 l=1.3e-07 w=1.5e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=1.5e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRHQX4MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS RN net128 VPW n12 l=1.3e-07 w=5.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=5.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP14 net065 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.9e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 pm nmsi p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
MX_t10_2 m pm VDD VNW p12 l=1.3e-07 w=5.1e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 bm RN VDD VNW p12 l=1.3e-07 w=3e-07
MXP16 bm c net109 VNW p12 l=1.3e-07 w=1.5e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=1.5e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRHQX8MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS RN net128 VPW n12 l=1.3e-07 w=5.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=5.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP14 net065 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.9e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 pm nmsi p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
MX_t10_2 m pm VDD VNW p12 l=1.3e-07 w=5.1e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 bm RN VDD VNW p12 l=1.3e-07 w=3e-07
MXP16 bm c net109 VNW p12 l=1.3e-07 w=1.5e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=1.5e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRQX1MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net130 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net130 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net138 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MX_t9 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN7 pm c net123 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net118 m net123 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net118 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE net76 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE net76 cn XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 s net76 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net97 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 nmrs SE net97 VNW p12 l=1.3e-07 w=3e-07
MXP1 nmrs nmse net105 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net105 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI74_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN net76 cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN net76 c XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s net76 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFRQX2MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net130 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net130 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net138 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MX_t9 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm c net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 net118 m net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN6 net118 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE net76 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE net76 cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1 s net76 XI1_n1 VPW n12 l=1.3e-07 w=2.7e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net97 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 nmrs SE net97 VNW p12 l=1.3e-07 w=3e-07
MXP1 nmrs nmse net105 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net105 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI74_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm cn net89 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD m net89 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN net76 cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN net76 c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s net76 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRQX4MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net130 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net130 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net138 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MX_t9 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm c net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 net118 m net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN6 net118 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE net76 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE net76 cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1 s net76 XI1_n1 VPW n12 l=1.3e-07 w=4.9e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net97 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 nmrs SE net97 VNW p12 l=1.3e-07 w=3e-07
MXP1 nmrs nmse net105 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net105 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI74_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm cn net89 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD m net89 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN net76 cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN net76 c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 s net76 VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRX1MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net104 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MXN9 nmrs nmse net104 VPW n12 l=1.3e-07 w=2.4e-07
MXN7 nmrs SE net77 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net77 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN12 pm c net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN13 net83 m net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net83 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNOE bm cn XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 s bm XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net139 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP10 nmrs SE net139 VNW p12 l=1.3e-07 w=3e-07
MXP8 nmrs nmse net115 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net115 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm cn net124 VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD m net124 VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPOEN bm c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFRX2MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net104 D net_clr_ VPW n12 l=1.3e-07 w=2.5e-07
MXN9 nmrs nmse net104 VPW n12 l=1.3e-07 w=2.5e-07
MXN7 nmrs SE net77 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net77 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.9e-07
MXN12 pm c net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN16 net83 m net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN17 net83 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.2e-07
mXI0_MXNOE bm cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1 s bm XI1_n1 VPW n12 l=1.3e-07 w=2.7e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net139 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP10 nmrs SE net139 VNW p12 l=1.3e-07 w=3e-07
MXP8 nmrs nmse net115 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net115 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP13 pm cn net124 VNW p12 l=1.3e-07 w=1.5e-07
MXP12 VDD m net124 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.4e-07
mXI0_MXPOEN bm c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRX4MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net104 D net_clr_ VPW n12 l=1.3e-07 w=4.9e-07
MXN9 nmrs nmse net104 VPW n12 l=1.3e-07 w=4.9e-07
MXN7 nmrs SE net77 VPW n12 l=1.3e-07 w=2.4e-07
MXN16 net77 SI net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MXN11 net_clr_ RN VSS VPW n12 l=1.3e-07 w=6.5e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=3.7e-07
MXN12 pm c net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN18 net83 m net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN19 net83 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=6.4e-07
mXI0_MXNOE bm cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1 s bm XI1_n1 VPW n12 l=1.3e-07 w=4.4e-07
mXI70_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI70_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net139 D VDD VNW p12 l=1.3e-07 w=6e-07
MXP14 nmrs SE net139 VNW p12 l=1.3e-07 w=6e-07
MXP13 nmrs nmse net115 VNW p12 l=1.3e-07 w=2.9e-07
MXP7 net115 SI VDD VNW p12 l=1.3e-07 w=2.9e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=3.9e-07
MXP15 pm cn net124 VNW p12 l=1.3e-07 w=1.5e-07
MXP12 VDD m net124 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.4e-07
mXI0_MXPOEN bm c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mXI70_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI70_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSHQX1MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net0112 SN VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN3 net169 cn net0112 VPW n12 l=1.3e-07 w=4.5e-07
MX_t11 pm nmsi net169 VPW n12 l=1.3e-07 w=4.5e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP3 net088 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=3e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm nmsi net56 VNW p12 l=1.3e-07 w=3.7e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT SDFFSHQX2MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.4e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net0104 SN VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN8 net169 cn net0104 VPW n12 l=1.3e-07 w=6.5e-07
MX_t11 pm nmsi net169 VPW n12 l=1.3e-07 w=6.5e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP8 net088 c cn VNW p12 l=1.3e-07 w=4.9e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=4.2e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=4.2e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=2.3e-07
MXP9 pm nmsi net56 VNW p12 l=1.3e-07 w=5.4e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.01e-06
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSHQX4MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net0104 SN VSS VPW n12 l=1.3e-07 w=7.4e-07
MXN10 net169 cn net0104 VPW n12 l=1.3e-07 w=7.4e-07
MX_t11 pm nmsi net169 VPW n12 l=1.3e-07 w=7.4e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.9e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP10 net088 c cn VNW p12 l=1.3e-07 w=5.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=3.8e-07
MXP11 pm nmsi net56 VNW p12 l=1.3e-07 w=6.9e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSHQX8MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net0104 SN VSS VPW n12 l=1.3e-07 w=7.5e-07
MXN12 net169 cn net0104 VPW n12 l=1.3e-07 w=7.5e-07
MXN13 pm nmsi net169 VPW n12 l=1.3e-07 w=7.5e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.9e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP10 net088 c cn VNW p12 l=1.3e-07 w=5.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=3.8e-07
MXP11 pm nmsi net56 VNW p12 l=1.3e-07 w=6.9e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSQX1MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmrs SE net150 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net150 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net123 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 nmrs nmse net123 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN11 bm cn net141 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 NSN s net141 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 nmrs SE net83 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net83 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 VDD SI net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net113 nmse nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 VDD pm m VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD SN m VNW p12 l=1.3e-07 w=2.3e-07
MXP13 VDD SN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP14 net107 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP15 net107 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSQX2MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmrs SE net150 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net150 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net123 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 nmrs nmse net123 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN11 bm cn net141 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 NSN s net141 VPW n12 l=1.3e-07 w=1.5e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 nmrs SE net83 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net83 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 VDD SI net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net113 nmse nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 VDD pm m VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD SN m VNW p12 l=1.3e-07 w=2.3e-07
MXP13 VDD SN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP16 net107 c bm VNW p12 l=1.3e-07 w=1.5e-07
MXP15 net107 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSQX4MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmrs SE net150 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net150 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net123 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 nmrs nmse net123 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN11 bm cn net141 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 NSN s net141 VPW n12 l=1.3e-07 w=1.5e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 nmrs SE net83 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net83 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 VDD SI net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net113 nmse nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 VDD pm m VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD SN m VNW p12 l=1.3e-07 w=2.3e-07
MXP13 VDD SN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP16 net107 c bm VNW p12 l=1.3e-07 w=1.5e-07
MXP15 net107 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRHQX1MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 net142 SN VSS VPW n12 l=1.3e-07 w=4.1e-07
MXN12 net166 cn net142 VPW n12 l=1.3e-07 w=4.1e-07
MX_t25 pm nmsi net166 VPW n12 l=1.3e-07 w=4.1e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=4.3e-07
MXN14 net170 RN VSS VPW n12 l=1.3e-07 w=4.3e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP12 net111 c cn VNW p12 l=1.3e-07 w=4.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmsi net131 VNW p12 l=1.3e-07 w=3.1e-07
MX_t28 net131 c VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 m RN net117 VNW p12 l=1.3e-07 w=2.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.6e-07
MXP21 bm nmset net93 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSRHQX2MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 net142 SN VSS VPW n12 l=1.3e-07 w=5.9e-07
MXN19 net166 cn net142 VPW n12 l=1.3e-07 w=5.9e-07
MXN20 pm nmsi net166 VPW n12 l=1.3e-07 w=5.9e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=6.1e-07
MXN21 net170 RN VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP12 net111 c cn VNW p12 l=1.3e-07 w=4.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmsi net131 VNW p12 l=1.3e-07 w=4.5e-07
MXP22 net131 c VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 m RN net117 VNW p12 l=1.3e-07 w=2.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP23 bm nmset net93 VNW p12 l=1.3e-07 w=2.7e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRHQX4MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN20 net142 SN VSS VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net166 cn net142 VPW n12 l=1.3e-07 w=7.5e-07
MX_t25 pm nmsi net166 VPW n12 l=1.3e-07 w=7.5e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=7.2e-07
MXN21 net170 RN VSS VPW n12 l=1.3e-07 w=7.2e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN22 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP22 net111 c cn VNW p12 l=1.3e-07 w=5.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.2e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.9e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP23 pm nmsi net131 VNW p12 l=1.3e-07 w=6.8e-07
MX_t28 net131 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP26 m RN net117 VNW p12 l=1.3e-07 w=3.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP27 bm nmset net93 VNW p12 l=1.3e-07 w=3.6e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRHQX8MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN20 net142 SN VSS VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net166 cn net142 VPW n12 l=1.3e-07 w=7.5e-07
MX_t25 pm nmsi net166 VPW n12 l=1.3e-07 w=7.5e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=7.2e-07
MXN21 net170 RN VSS VPW n12 l=1.3e-07 w=7.2e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN22 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP22 net111 c cn VNW p12 l=1.3e-07 w=5.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.2e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.9e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP23 pm nmsi net131 VNW p12 l=1.3e-07 w=6.8e-07
MX_t28 net131 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP26 m RN net117 VNW p12 l=1.3e-07 w=3.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP27 bm nmset net93 VNW p12 l=1.3e-07 w=3.6e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRX1MTR Q QN VDD VNW VPW VSS CK D RN SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE pm c XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MX_t15 NSN NRN m VPW n12 l=1.3e-07 w=1.9e-07
mXI60_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MXN5 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MX_t20 bm cn net75 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN s net75 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN pm cn XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 brn NRN VDD VNW p12 l=1.3e-07 w=4.9e-07
MX_t11 m pm brn VNW p12 l=1.3e-07 w=3.6e-07
MX_t12 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t16 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MXP6 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 brn s net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSRX2MTR Q QN VDD VNW VPW VSS CK D RN SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE pm c XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MX_t15 NSN NRN m VPW n12 l=1.3e-07 w=1.9e-07
mXI60_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MXN5 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MX_t20 bm cn net75 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN s net75 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN pm cn XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 brn NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP7 m pm brn VNW p12 l=1.3e-07 w=4.4e-07
MX_t12 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t16 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.4e-07
MXP6 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 brn s net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRX4MTR Q QN VDD VNW VPW VSS CK D RN SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=2.5e-07
mXI8_MXNOE pm c XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MX_t15 NSN NRN m VPW n12 l=1.3e-07 w=1.9e-07
mXI60_MXNOE bm c m VPW n12 l=1.3e-07 w=4.7e-07
MXN5 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MX_t20 bm cn net91 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN s net91 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=3e-07
mXI8_MXPOEN pm cn XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 brn NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP7 m pm brn VNW p12 l=1.3e-07 w=4.4e-07
MX_t12 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t16 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.7e-07
MXP6 bm c net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 brn s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSX1MTR Q QN VDD VNW VPW VSS CK D SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE pm c XI2_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNA1 XI2_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t11 m pm BSN VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MX_t19 bm cn net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 BSN s net138 VPW n12 l=1.3e-07 w=1.8e-07
MX_t33 BSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI33_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN pm cn XI2_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPA1 XI2_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MX_t24 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 bm c net104 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 VDD s net104 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI33_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSX2MTR Q QN VDD VNW VPW VSS CK D SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE pm c XI2_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNA1 XI2_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
MX_t11 m pm BSN VPW n12 l=1.3e-07 w=2.1e-07
MX_t11_2 m pm BSN VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MX_t19 bm cn net138 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN s net138 VPW n12 l=1.3e-07 w=1.5e-07
MX_t33 BSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN pm cn XI2_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPA1 XI2_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.4e-07
MX_t24 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm c net104 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD s net104 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI34_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSX4MTR Q QN VDD VNW VPW VSS CK D SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=2e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=2e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=2e-07
mXI2_MXNOE pm c XI2_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNA1 XI2_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.8e-07
MX_t11 m pm BSN VPW n12 l=1.3e-07 w=3.5e-07
MX_t11_2 m pm BSN VPW n12 l=1.3e-07 w=3.5e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.2e-07
MX_t19 bm cn net138 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN s net138 VPW n12 l=1.3e-07 w=1.5e-07
MX_t33 BSN SN VSS VPW n12 l=1.3e-07 w=1.08e-06
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI35_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI35_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=2.8e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=2.8e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.4e-07
mXI2_MXPOEN pm cn XI2_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPA1 XI2_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=7.8e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
MX_t24 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm c net104 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD s net104 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.9e-07
mXI35_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI35_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFTRX1MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net074 RN VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN5 net181 D net074 VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net181 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net193 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net193 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE bm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net96 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP7 nmrs SE net96 VNW p12 l=1.3e-07 w=3e-07
MXP6 nmrs nmse net114 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net114 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net105 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmrs RN net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI43_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI8_MXPOEN bm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFTRX2MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net074 RN VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN5 net181 D net074 VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net181 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net193 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net193 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mXI43_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI8_MXNOE bm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI47_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net96 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP7 nmrs SE net96 VNW p12 l=1.3e-07 w=3e-07
MXP6 nmrs nmse net114 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net114 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net105 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmrs RN net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI43_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI8_MXPOEN bm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFTRX4MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net074 RN VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN8 net181 D net074 VPW n12 l=1.3e-07 w=4.2e-07
MX_t7 nmrs nmse net181 VPW n12 l=1.3e-07 w=4.2e-07
MX_t3 nmrs SE net193 VPW n12 l=1.3e-07 w=2.3e-07
MXN7 net193 SI VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI43_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=3.4e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=8e-07
mXI8_MXNOE bm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI49_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI49_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net96 D VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP11 nmrs SE net96 VNW p12 l=1.3e-07 w=5.4e-07
MXP10 nmrs nmse net114 VNW p12 l=1.3e-07 w=2.7e-07
MX_t1 net114 SI VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP8 net105 SE VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP13 nmrs RN net105 VNW p12 l=1.3e-07 w=2.7e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI43_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=4.1e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_3 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_4 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI8_MXPOEN bm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=4.3e-07
mXI49_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI49_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFX1MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net137 SE net116 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net116 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net137 D net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 pm cn net137 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNOE pm c XI17_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 XI17_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI57_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI15_MXNOE sn c XI15_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI16_MXNOE sn cn XI16_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI16_MXNA1 XI16_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI58_MXNA1 Q sn VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 s sn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net77 nmse net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net73 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net76 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net77 D net76 VNW p12 l=1.3e-07 w=3.8e-07
MXP4 pm c net77 VNW p12 l=1.3e-07 w=3.8e-07
mXI17_MXPOEN pm cn XI17_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPA1 XI17_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI57_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI15_MXPOEN sn cn XI15_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI16_MXPOEN sn c XI16_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI16_MXPA1 XI16_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s sn VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPA1 Q sn VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFX2MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net137 SE net116 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net116 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net137 D net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 pm cn net137 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNOE pm c XI17_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 XI17_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI57_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI15_MXNOE sn c XI15_n1 VPW n12 l=1.3e-07 w=3.5e-07
mXI16_MXNOE sn cn XI16_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI16_MXNA1 XI16_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s sn VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI61_MXNA1 Q sn VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP5 net77 nmse net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net73 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net76 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net77 D net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm c net77 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPOEN pm cn XI17_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI17_MXPA1 XI17_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI57_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI15_MXPOEN sn cn XI15_p1 VNW p12 l=1.3e-07 w=4.9e-07
mXI16_MXPOEN sn c XI16_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI16_MXPA1 XI16_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s sn VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI61_MXPA1 Q sn VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT SDFFX4MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net137 SE net116 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net116 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net137 D net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 pm cn net137 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNOE pm c XI17_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 XI17_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI57_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=5.8e-07
mXI15_MXNOE sn c XI15_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI16_MXNOE sn cn XI16_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI16_MXNA1 XI16_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s sn VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI62_MXNA1 Q sn VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI62_MXNA1_2 Q sn VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP5 net77 nmse net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net73 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net76 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net77 D net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm c net77 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPOEN pm cn XI17_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI17_MXPA1 XI17_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=4.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI57_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI15_MXPOEN sn cn XI15_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI16_MXPOEN sn c XI16_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI16_MXPA1 XI16_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s sn VDD VNW p12 l=1.3e-07 w=4.2e-07
mXI62_MXPA1 Q sn VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI62_MXPA1_2 Q sn VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT SEDFFHQX1MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=2.3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=3.6e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.4e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=3e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP4 net079 c cn VNW p12 l=1.3e-07 w=4.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP5 pm nmsi net78 VNW p12 l=1.3e-07 w=4.4e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.4e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SEDFFHQX2MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=5.1e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=5.6e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=3.9e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP6 net079 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 pm nmsi net78 VNW p12 l=1.3e-07 w=6.2e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFHQX4MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=5.1e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=7e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.8e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 net079 c cn VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.8e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 pm nmsi net78 VNW p12 l=1.3e-07 w=6.2e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFHQX8MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=5.1e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=7e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.8e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 net079 c cn VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.8e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 pm nmsi net78 VNW p12 l=1.3e-07 w=6.2e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFTRX1MTR Q QN VDD VNW VPW VSS CK D E RN SE SI
MX_t9 nmrs RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmrs SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI44_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmsi SI VSS VPW n12 l=1.3e-07 w=1.7e-07
mXI38_MXNOE nmin_pass2 bse nmsi VPW n12 l=1.3e-07 w=1.8e-07
mXI39_MXNOE nmin_pass2 nmse nmin_pass1 VPW n12 l=1.3e-07 w=1.8e-07
mXI45_MXNA1 bse nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNOE nmin_pass1 be nmin VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE nmin_pass1 nmen s VPW n12 l=1.3e-07 w=1.8e-07
mX_g12_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 be nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net169 nmrs VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t5 net169 nmin_pass2 VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t4 pm cn net169 VPW n12 l=1.3e-07 w=2e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g18_MXNA1 nm m VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI59_MXNOE bnm c nm VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNOE bnm cn XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI46_MXNA1 QN bnm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP4 nmrs RN net108 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net108 SE VDD VNW p12 l=1.3e-07 w=3e-07
mXI44_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmsi SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI38_MXPOEN nmin_pass2 nmse nmsi VNW p12 l=1.3e-07 w=2.3e-07
mXI39_MXPOEN nmin_pass2 bse nmin_pass1 VNW p12 l=1.3e-07 w=2.3e-07
mXI45_MXPA1 bse nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPOEN nmin_pass1 nmen nmin VNW p12 l=1.3e-07 w=2.3e-07
mXI40_MXPOEN nmin_pass1 be s VNW p12 l=1.3e-07 w=2.3e-07
mX_g12_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 be nmen VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
MX_t1 net102 nmrs VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net111 nmin_pass2 net102 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 pm c net111 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g18_MXPA1 nm m VDD VNW p12 l=1.3e-07 w=4.1e-07
mXI59_MXPOEN bnm cn nm VNW p12 l=1.3e-07 w=4.1e-07
mXI1_MXPOEN bnm c XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI46_MXPA1 QN bnm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SEDFFTRX2MTR Q QN VDD VNW VPW VSS CK D E RN SE SI
MX_t9 nmrs RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmrs SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI44_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmsi SI VSS VPW n12 l=1.3e-07 w=1.7e-07
mXI38_MXNOE nmin_pass2 bse nmsi VPW n12 l=1.3e-07 w=1.8e-07
mXI39_MXNOE nmin_pass2 nmse nmin_pass1 VPW n12 l=1.3e-07 w=1.8e-07
mXI45_MXNA1 bse nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNOE nmin_pass1 be nmin VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE nmin_pass1 nmen s VPW n12 l=1.3e-07 w=1.8e-07
mX_g12_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 be nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN5 net169 nmrs VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t5 net169 nmin_pass2 VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t4 pm cn net169 VPW n12 l=1.3e-07 w=2e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g18_MXNA1 nm m VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE bnm c nm VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNOE bnm cn XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI47_MXNA1 QN bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmrs RN net108 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net108 SE VDD VNW p12 l=1.3e-07 w=3e-07
mXI44_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmsi SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI38_MXPOEN nmin_pass2 nmse nmsi VNW p12 l=1.3e-07 w=2.3e-07
mXI39_MXPOEN nmin_pass2 bse nmin_pass1 VNW p12 l=1.3e-07 w=2.3e-07
mXI45_MXPA1 bse nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPOEN nmin_pass1 nmen nmin VNW p12 l=1.3e-07 w=2.3e-07
mXI40_MXPOEN nmin_pass1 be s VNW p12 l=1.3e-07 w=2.3e-07
mX_g12_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 be nmen VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t1 net102 nmrs VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net111 nmin_pass2 net102 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 pm c net111 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g18_MXPA1 nm m VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI59_MXPOEN bnm cn nm VNW p12 l=1.3e-07 w=5.9e-07
mXI1_MXPOEN bnm c XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI47_MXPA1 QN bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFTRX4MTR Q QN VDD VNW VPW VSS CK D E RN SE SI
MX_t9 nmrs RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmrs SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI44_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmsi SI VSS VPW n12 l=1.3e-07 w=1.7e-07
mXI38_MXNOE nmin_pass2 bse nmsi VPW n12 l=1.3e-07 w=1.8e-07
mXI39_MXNOE nmin_pass2 nmse nmin_pass1 VPW n12 l=1.3e-07 w=1.8e-07
mXI45_MXNA1 bse nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNOE nmin_pass1 be nmin VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE nmin_pass1 nmen s VPW n12 l=1.3e-07 w=1.8e-07
mX_g12_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 be nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN5 net169 nmrs VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t5 net169 nmin_pass2 VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t4 pm cn net169 VPW n12 l=1.3e-07 w=2e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g18_MXNA1 nm m VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE bnm c nm VPW n12 l=1.3e-07 w=7.4e-07
mXI1_MXNOE bnm cn XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI48_MXNA1 QN bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI48_MXNA1_2 QN bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmrs RN net108 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net108 SE VDD VNW p12 l=1.3e-07 w=3e-07
mXI44_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmsi SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI38_MXPOEN nmin_pass2 nmse nmsi VNW p12 l=1.3e-07 w=2.3e-07
mXI39_MXPOEN nmin_pass2 bse nmin_pass1 VNW p12 l=1.3e-07 w=2.3e-07
mXI45_MXPA1 bse nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPOEN nmin_pass1 nmen nmin VNW p12 l=1.3e-07 w=2.3e-07
mXI40_MXPOEN nmin_pass1 be s VNW p12 l=1.3e-07 w=2.3e-07
mX_g12_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 be nmen VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t1 net102 nmrs VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net111 nmin_pass2 net102 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 pm c net111 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.9e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g18_MXPA1 nm m VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI59_MXPOEN bnm cn nm VNW p12 l=1.3e-07 w=8e-07
mXI1_MXPOEN bnm c XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI48_MXPA1 QN bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI48_MXPA1_2 QN bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFX1MTR Q QN VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net180 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net187 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net190 SE net187 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net190 D net181 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net181 E net180 VPW n12 l=1.3e-07 w=1.8e-07
MX_t16 net196 nmen net180 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net196 s net190 VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 pm cn net190 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI3_MXNOE nm c XI3_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI4_MXNOE nm cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI41_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t6 net85 SE VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t8 net97 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net96 nmse net97 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net96 D net91 VNW p12 l=1.3e-07 w=4.7e-07
MX_t5 net91 nmen net85 VNW p12 l=1.3e-07 w=4.7e-07
MXP9 net88 E net85 VNW p12 l=1.3e-07 w=4.7e-07
MXP10 net88 s net96 VNW p12 l=1.3e-07 w=4.7e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm c net96 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI40_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI3_MXPOEN nm cn XI3_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI4_MXPOEN nm c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.4e-07
mXI41_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SEDFFX2MTR Q QN VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net100 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net92 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net88 SE net92 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net88 D net76 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net76 E net100 VPW n12 l=1.3e-07 w=1.8e-07
MX_t16 net84 nmen net100 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net84 s net88 VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 pm cn net88 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI3_MXNOE nm c XI3_n1 VPW n12 l=1.3e-07 w=4.4e-07
mXI4_MXNOE nm cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI42_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t6 net127 SE VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t8 net111 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net113 nmse net111 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net113 D net131 VNW p12 l=1.3e-07 w=4.7e-07
MX_t5 net131 nmen net127 VNW p12 l=1.3e-07 w=4.7e-07
MXP9 net105 E net127 VNW p12 l=1.3e-07 w=4.7e-07
MXP10 net105 s net113 VNW p12 l=1.3e-07 w=4.7e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm c net113 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI40_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI3_MXPOEN nm cn XI3_p1 VNW p12 l=1.3e-07 w=5.4e-07
mXI4_MXPOEN nm c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI42_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFX4MTR Q QN VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net100 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net92 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net88 SE net92 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net88 D net76 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net76 E net100 VPW n12 l=1.3e-07 w=1.8e-07
MX_t16 net84 nmen net100 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net84 s net88 VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 pm cn net88 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI40_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI3_MXNOE nm c XI3_n1 VPW n12 l=1.3e-07 w=6.4e-07
mXI4_MXNOE nm cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI43_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI43_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 net127 SE VDD VNW p12 l=1.3e-07 w=2.4e-07
MXP14_2 net127 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net111 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net113 nmse net111 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net113 D net131 VNW p12 l=1.3e-07 w=4.7e-07
MX_t5 net131 nmen net127 VNW p12 l=1.3e-07 w=4.7e-07
MXP12 net105 E net127 VNW p12 l=1.3e-07 w=4.6e-07
MXP13 net105 s net113 VNW p12 l=1.3e-07 w=4.6e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm c net113 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI40_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI3_MXPOEN nm cn XI3_p1 VNW p12 l=1.3e-07 w=7.3e-07
mXI4_MXPOEN nm c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI43_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI43_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SMDFFHQX1MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=1.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=2.1e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN4 VSS cn net107 VPW n12 l=1.3e-07 w=3.3e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=3.3e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=3.7e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=2.6e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=2.6e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=3e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=3e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=4.2e-07
MXP0 cn c net085 VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=4e-07
MXP3 pm nmsi net060 VNW p12 l=1.3e-07 w=4e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=7.3e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SMDFFHQX2MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=1.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=3.1e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=3e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN5 VSS cn net107 VPW n12 l=1.3e-07 w=4.8e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=4.8e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=4.4e-07
MXP4 cn c net085 VNW p12 l=1.3e-07 w=4.4e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP5 pm nmsi net060 VNW p12 l=1.3e-07 w=5.9e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=9.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=9.8e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SMDFFHQX4MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=2.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=5e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN6 VSS cn net107 VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=5.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=3.4e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net085 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net060 VNW p12 l=1.3e-07 w=1.01e-06
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SMDFFHQX8MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=2.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=5e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN6 VSS cn net107 VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=5.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=3.4e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net085 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net060 VNW p12 l=1.3e-07 w=1.01e-06
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX12MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=3.2e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=5e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=4.5e-07
MXN3_2 nmin OE net31 VPW n12 l=1.3e-07 w=4.5e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN0_3 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_5 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_6 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=3.9e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=6.5e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=3e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=8e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP0_3 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_5 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX16MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=4.1e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN3_2 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN0_3 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_5 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_6 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_7 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_8 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=8e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=5.2e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=8.6e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_3 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_5 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_7 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_8 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX1MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TBUFX20MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=5.2e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=4.4e-07
MXN4_2 net31 nmen VSS VPW n12 l=1.3e-07 w=4.4e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=6.5e-07
MXN3_2 nmin OE net31 VPW n12 l=1.3e-07 w=6.5e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_3 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_4 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_5 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_6 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_7 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_8 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_9 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_10 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP4_2 nmin OE VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=8e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=8e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_3 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_4 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_5 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_7 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_8 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_9 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_10 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX24MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=6.3e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=5.2e-07
MXN4_2 net31 nmen VSS VPW n12 l=1.3e-07 w=5.2e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN3_2 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN3_3 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_3 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_4 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_5 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_5 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_6 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_7 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_8 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_9 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_10 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_11 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_12 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=7.7e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP5_3 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP5_4 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=6.6e-07
MXP4_2 nmin OE VDD VNW p12 l=1.3e-07 w=6.6e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_3 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_4 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_5 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_5 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_7 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_8 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_9 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_10 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_11 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_12 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX2MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=3e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=7e-07
.ends


.SUBCKT TBUFX3MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=2.3e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=3e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=6.6e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT TBUFX4MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=3e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=3.6e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
.ends


.SUBCKT TBUFX6MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=3e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=3.7e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
.ends


.SUBCKT TBUFX8MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=3e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=6.4e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=3e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=5e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TIEHIMTR Y VDD VNW VPW VSS
MXNhi lo hi VSS VPW n12 l=1.3e-07 w=1.5e-07
MXNlo lo lo VSS VPW n12 l=1.3e-07 w=1.5e-07
MXPlo1 hi lo VDD VNW p12 l=1.3e-07 w=1.5e-07
MXPlo2 Y lo VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TIELOMTR Y VDD VNW VPW VSS
MXNhi1 lo hi VSS VPW n12 l=1.3e-07 w=1.5e-07
MXNhi2 Y hi VSS VPW n12 l=1.3e-07 w=3.6e-07
MXPlo hi lo VDD VNW p12 l=1.3e-07 w=1.5e-07
MXPhi hi hi VDD VNW p12 l=1.3e-07 w=1.5e-07
.ends


.SUBCKT TLATNCAX12MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_3 XI14_n1__3 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_3 nmin c XI14_n1__3 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_4 nmin c XI14_n1__4 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_4 XI14_n1__4 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_5 XI14_n1__5 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_5 nmin c XI14_n1__5 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=2.9e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=2.9e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_2 ECK nmin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_3 ECK nmin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=7.9e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_3 XI14_p1__3 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPOEN_3 nmin cn XI14_p1__3 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPOEN_4 nmin cn XI14_p1__4 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_4 XI14_p1__4 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_5 XI14_p1__5 E VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPOEN_5 nmin cn XI14_p1__5 VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK nmin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK nmin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK nmin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX16MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_3 XI14_n1__3 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_3 nmin c XI14_n1__3 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_4 nmin c XI14_n1__4 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_4 XI14_n1__4 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_5 XI14_n1__5 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_5 nmin c XI14_n1__5 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_2 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_3 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=8.1e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_3 XI14_p1__3 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPOEN_3 nmin cn XI14_p1__3 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPOEN_4 nmin cn XI14_p1__4 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_4 XI14_p1__4 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_5 XI14_p1__5 E VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPOEN_5 nmin cn XI14_p1__5 VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK nmin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK nmin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK nmin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 ECK nmin XI1_p1__7 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_7 XI1_p1__7 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_8 XI1_p1__8 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 ECK nmin XI1_p1__8 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX20MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_3 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_4 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_5 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1_3 XI14_n1__3 E VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNOE_3 nmin c XI14_n1__3 VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNOE_4 nmin c XI14_n1__4 VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1_4 XI14_n1__4 E VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1_5 XI14_n1__5 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_5 nmin c XI14_n1__5 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_6 nmin c XI14_n1__6 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_6 XI14_n1__6 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_7 XI14_n1__7 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_7 nmin c XI14_n1__7 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_2 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_3 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA2_4 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_4 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_4 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_5 c CK VDD VNW p12 l=1.3e-07 w=8.1e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPA1_3 XI14_p1__3 E VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPOEN_3 nmin cn XI14_p1__3 VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPOEN_4 nmin cn XI14_p1__4 VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPA1_4 XI14_p1__4 E VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPA1_5 XI14_p1__5 E VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI14_MXPOEN_5 nmin cn XI14_p1__5 VNW p12 l=1.3e-07 w=7.1e-07
mXI14_MXPOEN_6 nmin cn XI14_p1__6 VNW p12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1_6 XI14_p1__6 E VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1_7 XI14_p1__7 E VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI14_MXPOEN_7 nmin cn XI14_p1__7 VNW p12 l=1.3e-07 w=6.8e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.8e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK nmin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK nmin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK nmin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 ECK nmin XI1_p1__7 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_7 XI1_p1__7 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_8 XI1_p1__8 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 ECK nmin XI1_p1__8 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_9 ECK nmin XI1_p1__9 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_9 XI1_p1__9 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_10 XI1_p1__10 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_10 ECK nmin XI1_p1__10 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX2MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX3MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.8e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX4MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=3e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=4.3e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=4.3e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=5.9e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=5.9e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX6MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=5.6e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX8MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_2 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK nmin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNSRX1MTR Q QN VDD VNW VPW VSS D GN RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=4e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=3.7e-07
MXN7 net048 D VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN6 net052 RN net048 VPW n12 l=1.3e-07 w=5.3e-07
MX_t13 pm c net052 VPW n12 l=1.3e-07 w=5.3e-07
MX_t2 pm cn net98 VPW n12 l=1.3e-07 w=2.8e-07
MXN8 net98 RN net101 VPW n12 l=1.3e-07 w=2.8e-07
MXN9 VSS m net101 VPW n12 l=1.3e-07 w=2.8e-07
mX_g4_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 c GN VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI47_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI46_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP11 pm nms net61 VNW p12 l=1.3e-07 w=6.3e-07
MX_t14 net61 RN VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t9 net083 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP9 net075 nms net083 VNW p12 l=1.3e-07 w=6.4e-07
MXP10 pm cn net075 VNW p12 l=1.3e-07 w=6.4e-07
MXP13 pm c net70 VNW p12 l=1.3e-07 w=3.2e-07
MXP12 net70 nms net67 VNW p12 l=1.3e-07 w=3.2e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3.2e-07
mX_g4_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 c GN VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI47_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI46_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TLATNSRX2MTR Q QN VDD VNW VPW VSS D GN RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=6.2e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN7_2 net048__2 D VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN6_2 net052__2 RN net048__2 VPW n12 l=1.3e-07 w=5.3e-07
MX_t13_2 pm c net052__2 VPW n12 l=1.3e-07 w=5e-07
MX_t13 pm c net052 VPW n12 l=1.3e-07 w=4.1e-07
MXN6 net052 RN net048 VPW n12 l=1.3e-07 w=2.6e-07
MXN7 net048 D VSS VPW n12 l=1.3e-07 w=3.7e-07
MX_t2 pm cn net98 VPW n12 l=1.3e-07 w=2.8e-07
MXN8 net98 RN net101 VPW n12 l=1.3e-07 w=2.8e-07
MXN9 VSS m net101 VPW n12 l=1.3e-07 w=2.8e-07
mX_g4_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g5_MXNA1 c GN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI48_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI46_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=7.5e-07
MXP18 pm nms net61 VNW p12 l=1.3e-07 w=8.8e-07
MX_t14 net61 RN VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t9_2 net083__2 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP16_2 net075__2 nms net083__2 VNW p12 l=1.3e-07 w=6.4e-07
MXP17_2 pm cn net075__2 VNW p12 l=1.3e-07 w=6.4e-07
MXP17 pm cn net075 VNW p12 l=1.3e-07 w=6.4e-07
MXP16 net075 nms net083 VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 net083 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 pm c net70 VNW p12 l=1.3e-07 w=3.2e-07
MXP12 net70 nms net67 VNW p12 l=1.3e-07 w=3.2e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3.2e-07
mX_g4_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g5_MXPA1 c GN VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.4e-07
mXI48_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI46_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNSRX4MTR Q QN VDD VNW VPW VSS D GN RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=5.9e-07
mX_g3_MXNA1_2 nms SN VSS VPW n12 l=1.3e-07 w=5.8e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t6_2 pm nms VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN7_2 net048__2 D VSS VPW n12 l=1.3e-07 w=5.1e-07
MXN6_2 net052__2 RN net048__2 VPW n12 l=1.3e-07 w=5.1e-07
MX_t13_2 pm c net052__2 VPW n12 l=1.3e-07 w=5e-07
MX_t13 pm c net052 VPW n12 l=1.3e-07 w=4.1e-07
MXN6 net052 RN net048 VPW n12 l=1.3e-07 w=2.6e-07
MXN7 net048 D VSS VPW n12 l=1.3e-07 w=3.9e-07
MX_t2 pm cn net98 VPW n12 l=1.3e-07 w=2.8e-07
MXN8 net98 RN net101 VPW n12 l=1.3e-07 w=2.8e-07
MXN9 VSS m net101 VPW n12 l=1.3e-07 w=2.8e-07
mX_g4_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g5_MXNA1 c GN VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI50_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI50_MXNA1_2 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI49_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI49_MXNA1_2 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1_2 nms SN VDD VNW p12 l=1.3e-07 w=7.2e-07
MXP18 pm nms net61 VNW p12 l=1.3e-07 w=8.8e-07
MX_t14 net61 RN VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t9_2 net083__2 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP16_2 net075__2 nms net083__2 VNW p12 l=1.3e-07 w=6.4e-07
MXP17_2 pm cn net075__2 VNW p12 l=1.3e-07 w=6.4e-07
MXP17 pm cn net075 VNW p12 l=1.3e-07 w=6.4e-07
MXP16 net075 nms net083 VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 net083 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 pm c net70 VNW p12 l=1.3e-07 w=3.2e-07
MXP12 net70 nms net67 VNW p12 l=1.3e-07 w=3.2e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3.2e-07
mX_g4_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g5_MXPA1 c GN VDD VNW p12 l=1.3e-07 w=8.2e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI50_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI50_MXPA1_2 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI49_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI49_MXPA1_2 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX12MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g6_MXNA1_3 c CK VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g6_MXNA1_4 c CK VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g7_MXNA1_2 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_4 X_g3_n1__4 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_4 csetin c X_g3_n1__4 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_5 csetin c X_g3_n1__5 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_5 X_g3_n1__5 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_6 X_g3_n1__6 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_6 csetin c X_g3_n1__6 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1_4 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=7.9e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=8.7e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g7_MXPA1_2 setin nmsetin VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1_4 X_g3_p1__4 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_4 csetin cn X_g3_p1__4 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_5 csetin cn X_g3_p1__5 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1_5 X_g3_p1__5 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1_6 X_g3_p1__6 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_6 csetin cn X_g3_p1__6 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK csetin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK csetin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX16MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_3 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_4 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_5 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g5_MXNA1_2 cn c VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g8_MXNA1_2 nmsetin E VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g8_MXNA2_2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g7_MXNA1_2 setin nmsetin VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g7_MXNA1_3 setin nmsetin VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=4.95e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=4.95e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=4.95e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=4.95e-07
mX_g3_MXNA1_4 X_g3_n1__4 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_4 csetin c X_g3_n1__4 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_5 csetin c X_g3_n1__5 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1_5 X_g3_n1__5 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1_6 X_g3_n1__6 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_6 csetin c X_g3_n1__6 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_7 csetin c X_g3_n1__7 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1_7 X_g3_n1__7 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1_8 X_g3_n1__8 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_8 csetin c X_g3_n1__8 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=5e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_3 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_4 ECK csetin VSS VPW n12 l=1.3e-07 w=2e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g6_MXPA1_4 c CK VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g6_MXPA1_5 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g5_MXPA1_2 cn c VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g8_MXPA2_2 X_g8_p1__2 SE VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1_2 nmsetin E X_g8_p1__2 VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g7_MXPA1_2 setin nmsetin VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g7_MXPA1_3 setin nmsetin VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=4.65e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=4.65e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=4.65e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=4.65e-07
mX_g3_MXPA1_4 X_g3_p1__4 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_4 csetin cn X_g3_p1__4 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_5 csetin cn X_g3_p1__5 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1_5 X_g3_p1__5 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1_6 X_g3_p1__6 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_6 csetin cn X_g3_p1__6 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_7 csetin cn X_g3_p1__7 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1_7 X_g3_p1__7 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1_8 X_g3_p1__8 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_8 csetin cn X_g3_p1__8 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK csetin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK csetin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK csetin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 ECK csetin XI1_p1__7 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_7 XI1_p1__7 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX20MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_3 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_4 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_5 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g5_MXNA1_2 cn c VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g8_MXNA1_2 nmsetin E VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g8_MXNA2_2 nmsetin SE VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g7_MXNA1_2 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g7_MXNA1_3 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=7.2e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=7.2e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNOE_4 csetin c X_g3_n1__4 VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_4 X_g3_n1__4 setin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_5 X_g3_n1__5 setin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNOE_5 csetin c X_g3_n1__5 VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNOE_6 csetin c X_g3_n1__6 VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_6 X_g3_n1__6 setin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_7 X_g3_n1__7 setin VSS VPW n12 l=1.3e-07 w=4.4e-07
mX_g3_MXNOE_7 csetin c X_g3_n1__7 VPW n12 l=1.3e-07 w=4.4e-07
mX_g3_MXNOE_8 csetin c X_g3_n1__8 VPW n12 l=1.3e-07 w=4.4e-07
mX_g3_MXNA1_8 X_g3_n1__8 setin VSS VPW n12 l=1.3e-07 w=4.4e-07
mX_g3_MXNA1_9 X_g3_n1__9 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_9 csetin c X_g3_n1__9 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA1_3 ECK csetin VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_4 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_5 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g5_MXPA1_2 cn c VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g8_MXPA2_2 X_g8_p1__2 SE VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1_2 nmsetin E X_g8_p1__2 VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=8.1e-07
mX_g7_MXPA1_2 setin nmsetin VDD VNW p12 l=1.3e-07 w=8.1e-07
mX_g7_MXPA1_3 setin nmsetin VDD VNW p12 l=1.3e-07 w=8e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=8e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=8e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_4 csetin cn X_g3_p1__4 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_4 X_g3_p1__4 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_5 X_g3_p1__5 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_5 csetin cn X_g3_p1__5 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_6 csetin cn X_g3_p1__6 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_6 X_g3_p1__6 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_7 X_g3_p1__7 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_7 csetin cn X_g3_p1__7 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_8 csetin cn X_g3_p1__8 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_8 X_g3_p1__8 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_9 X_g3_p1__9 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_9 csetin cn X_g3_p1__9 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK csetin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK csetin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK csetin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_7 XI1_p1__7 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 ECK csetin XI1_p1__7 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 ECK csetin XI1_p1__8 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_8 XI1_p1__8 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_9 XI1_p1__9 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_9 ECK csetin XI1_p1__9 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX2MTR ECK VDD VNW VPW VSS CK E SE
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=3e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=3e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX3MTR ECK VDD VNW VPW VSS CK E SE
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=3e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=3e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX4MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=3e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=3e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=3.2e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX6MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=3e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=4.4e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=4.6e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.3e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.9e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=8.8e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX8MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g7_MXNA1_2 setin nmsetin VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_4 X_g3_n1__4 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_4 csetin c X_g3_n1__4 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=5.9e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g7_MXPA1_2 setin nmsetin VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPA1_4 X_g3_p1__4 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN_4 csetin cn X_g3_p1__4 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=9e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=9e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI1_MXPA1_4 ECK csetin XI1_p1__4 VNW p12 l=1.3e-07 w=8.8e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNX1MTR Q QN VDD VNW VPW VSS D GN
mX_g5_MXNA1 cn GN VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 D VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI1_MXNOE pm cn XI1_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI21_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1 cn GN VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI1_MXPOEN pm c XI1_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI21_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TLATNX2MTR Q QN VDD VNW VPW VSS D GN
mX_g5_MXNA1 cn GN VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI1_MXNA1 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNOE pm cn XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI22_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 cn GN VDD VNW p12 l=1.3e-07 w=3.8e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI1_MXPA1 XI1_p1 D VDD VNW p12 l=1.3e-07 w=7e-07
mXI1_MXPOEN pm c XI1_p1 VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI22_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNX4MTR Q QN VDD VNW VPW VSS D GN
mX_g5_MXNA1 cn GN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI1_MXNA1 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNOE pm cn XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI24_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_2 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 cn GN VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 D VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI1_MXPOEN pm c XI1_p1 VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI24_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_2 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATSRX1MTR Q QN VDD VNW VPW VSS D G RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=3.1e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN1 net84 D VSS VPW n12 l=1.3e-07 w=3.9e-07
MXN0 net80 RN net84 VPW n12 l=1.3e-07 w=3.9e-07
MX_t13 pm c net80 VPW n12 l=1.3e-07 w=3.9e-07
MX_t2 pm cn net100 VPW n12 l=1.3e-07 w=2.6e-07
MXN2 net100 RN net105 VPW n12 l=1.3e-07 w=2.6e-07
MXN3 VSS m net105 VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3e-07
mX_g0_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP1 pm cn net47 VNW p12 l=1.3e-07 w=5.2e-07
MXP0 net47 nms net55 VNW p12 l=1.3e-07 w=5.2e-07
MX_t9 net55 D VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t14 net63 RN VDD VNW p12 l=1.3e-07 w=4.7e-07
MXP2 pm nms net63 VNW p12 l=1.3e-07 w=4.7e-07
MXP4 pm c net71 VNW p12 l=1.3e-07 w=3.2e-07
MXP3 net71 nms net67 VNW p12 l=1.3e-07 w=3.2e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3.2e-07
mX_g5_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g0_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TLATSRX2MTR Q QN VDD VNW VPW VSS D G RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=4.5e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=4e-07
MXN5 net84 D VSS VPW n12 l=1.3e-07 w=4.1e-07
MXN4 net80 RN net84 VPW n12 l=1.3e-07 w=4.1e-07
MX_t13 pm c net80 VPW n12 l=1.3e-07 w=4.1e-07
MX_t2 pm cn net100 VPW n12 l=1.3e-07 w=2.6e-07
MXN2 net100 RN net105 VPW n12 l=1.3e-07 w=2.6e-07
MXN3 VSS m net105 VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=2e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3e-07
mXI46_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP1 pm cn net47 VNW p12 l=1.3e-07 w=5.7e-07
MXP5 net47 nms net55 VNW p12 l=1.3e-07 w=8.6e-07
MX_t9 net55 D VDD VNW p12 l=1.3e-07 w=8.6e-07
MX_t14 net63 RN VDD VNW p12 l=1.3e-07 w=7.3e-07
MXP6 pm nms net63 VNW p12 l=1.3e-07 w=7.3e-07
MXP8 pm c net71 VNW p12 l=1.3e-07 w=3e-07
MXP7 net71 nms net67 VNW p12 l=1.3e-07 w=3e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI46_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATSRX4MTR Q QN VDD VNW VPW VSS D G RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=6.3e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=4e-07
MXN5 net84 D VSS VPW n12 l=1.3e-07 w=4.1e-07
MXN4 net80 RN net84 VPW n12 l=1.3e-07 w=4.1e-07
MX_t13 pm c net80 VPW n12 l=1.3e-07 w=4.1e-07
MX_t2 pm cn net100 VPW n12 l=1.3e-07 w=2.6e-07
MXN2 net100 RN net105 VPW n12 l=1.3e-07 w=2.6e-07
MXN3 VSS m net105 VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI46_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI46_MXNA1_2 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP1 pm cn net47 VNW p12 l=1.3e-07 w=5.7e-07
MXP5 net47 nms net55 VNW p12 l=1.3e-07 w=8.6e-07
MX_t9 net55 D VDD VNW p12 l=1.3e-07 w=8.6e-07
MX_t14 net63 RN VDD VNW p12 l=1.3e-07 w=7.3e-07
MXP6 pm nms net63 VNW p12 l=1.3e-07 w=7.3e-07
MXP8 pm c net71 VNW p12 l=1.3e-07 w=3e-07
MXP7 net71 nms net67 VNW p12 l=1.3e-07 w=3e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=4.2e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI46_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI46_MXPA1_2 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATX1MTR Q QN VDD VNW VPW VSS D G
mX_g6_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g5_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g3_MXNOE net52 c X_g3_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI5_MXNOE net52 cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m net52 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI25_MXNA1 Q net52 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g5_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g3_MXPOEN net52 cn X_g3_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI5_MXPOEN net52 c XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m net52 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI25_MXPA1 Q net52 VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TLATX2MTR Q QN VDD VNW VPW VSS D G
mX_g6_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=6.5e-07
mX_g3_MXNOE net52 c X_g3_n1 VPW n12 l=1.3e-07 w=6.5e-07
mXI5_MXNOE net52 cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m net52 VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI25_MXNA1 Q net52 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=8e-07
mX_g3_MXPOEN net52 cn X_g3_p1 VNW p12 l=1.3e-07 w=8e-07
mXI5_MXPOEN net52 c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 m net52 VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI25_MXPA1 Q net52 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATX4MTR Q QN VDD VNW VPW VSS D G
mX_g6_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g5_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNOE net52 c X_g3_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI5_MXNOE net52 cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m net52 VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI26_MXNA1 Q net52 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI26_MXNA1_2 Q net52 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g3_MXPOEN net52 cn X_g3_p1 VNW p12 l=1.3e-07 w=6.9e-07
mXI5_MXPOEN net52 c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 m net52 VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI26_MXPA1 Q net52 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI26_MXPA1_2 Q net52 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XNOR2X1MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=3e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=3e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=3.8e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=3.8e-07
.ends


.SUBCKT XNOR2X2MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=5.7e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=7.2e-07
.ends


.SUBCKT XNOR2X4MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_2 Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_2 Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN_2 Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=7.6e-07
mXI2_MXPOEN_2 Y A nb VNW p12 l=1.3e-07 w=7.6e-07
.ends


.SUBCKT XNOR2X8MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_3 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_4 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_2 Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_3 Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_4 Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_2 Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_3 Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_4 Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_3 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_4 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN_2 Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN_3 Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN_4 Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=7.6e-07
mXI2_MXPOEN_2 Y A nb VNW p12 l=1.3e-07 w=7.6e-07
mXI2_MXPOEN_3 Y A nb VNW p12 l=1.3e-07 w=7.6e-07
mXI2_MXPOEN_4 Y A nb VNW p12 l=1.3e-07 w=7.6e-07
.ends


.SUBCKT XNOR2XLMTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT XNOR3X1MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI52_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=3.7e-07
mXI53_MXNOE ny na bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI52_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=4.6e-07
mXI53_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT XNOR3X2MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=6e-07
mXI48_MXNOE ny na bnc VPW n12 l=1.3e-07 w=5.5e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI4_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI8_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=7.2e-07
mXI48_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=7.2e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XNOR3X4MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_2 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny na bnc VPW n12 l=1.3e-07 w=5.5e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.6e-07
mXI7_MXPA1_2 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI8_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=7.2e-07
mXI4_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=7.2e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XNOR3X8MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_2 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_3 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_4 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny na bnc VPW n12 l=1.3e-07 w=5.5e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.6e-07
mXI7_MXPA1_2 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.6e-07
mXI7_MXPA1_3 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI7_MXPA1_4 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI8_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=7.2e-07
mXI4_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=7.2e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XNOR3XLMTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=4.8e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=2e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=3e-07
mXI4_MXNOE ny na bnc VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=5.8e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=5.8e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=4.8e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI8_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=5.8e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT XOR2X1MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=3e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=3e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=3.8e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=3.8e-07
.ends


.SUBCKT XOR2X2MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=5.7e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=7.2e-07
.ends


.SUBCKT XOR2X3MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=4.5e-07
mXI2_MXNOE_2 Y A nb VPW n12 l=1.3e-07 w=4.5e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI4_MXNOE_2 Y na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=4.7e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=5.7e-07
mXI2_MXPOEN_2 Y na nb VNW p12 l=1.3e-07 w=5.7e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=5.7e-07
mXI4_MXPOEN_2 Y A bb VNW p12 l=1.3e-07 w=5.7e-07
.ends


.SUBCKT XOR2X4MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_2 Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_2 Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN_2 Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=7.6e-07
mXI4_MXPOEN_2 Y A bb VNW p12 l=1.3e-07 w=7.6e-07
.ends


.SUBCKT XOR2X8MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_3 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_4 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_2 Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_3 Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_4 Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_2 Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_3 Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_4 Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_3 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_4 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN_2 Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN_3 Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN_4 Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=7.6e-07
mXI4_MXPOEN_2 Y A bb VNW p12 l=1.3e-07 w=7.6e-07
mXI4_MXPOEN_3 Y A bb VNW p12 l=1.3e-07 w=7.6e-07
mXI4_MXPOEN_4 Y A bb VNW p12 l=1.3e-07 w=7.6e-07
.ends


.SUBCKT XOR2XLMTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT XOR3X1MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=3.7e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=4.6e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT XOR3X2MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=7.4e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XOR3X4MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_2 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI7_MXPA1_2 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=7.4e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XOR3X8MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_2 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_3 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_4 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI7_MXPA1_2 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI7_MXPA1_3 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI7_MXPA1_4 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=7.4e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XOR3XLMTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=4.8e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=3.7e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=2.1e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=5.8e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=5.8e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=4.8e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=2.5e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends

