* Hierarchy Level 0

* Top of hierarchy  cell=labhb1
.subckt labhb1 VDD QN Q GND RN D SN G
M1 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M4 N_22 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_22 RN N_21 GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_5 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 N_24 RN N_23 GND mn5  l=0.5u w=0.5u m=1
M10 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M11 Q N_7 GND GND mn5  l=0.5u w=0.58u m=1
M12 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_23 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_6 N_14 VDD mp5  l=0.42u w=0.52u m=1
M15 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_4 N_13 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_7 N_6 N_16 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 Q N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends labhb1
* SPICE INPUT		Wed Jul 10 13:40:34 2019	labhb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=labhb2
.subckt labhb2 VDD QN Q GND RN D SN G
M1 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M4 N_22 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_22 RN N_21 GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_5 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 N_24 RN N_23 GND mn5  l=0.5u w=0.5u m=1
M10 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M11 Q N_7 GND GND mn5  l=0.5u w=0.72u m=1
M12 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_23 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_6 N_14 VDD mp5  l=0.42u w=0.52u m=1
M15 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_4 N_13 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_7 N_6 N_16 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 Q N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends labhb2
* SPICE INPUT		Wed Jul 10 13:40:41 2019	lablb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb1
.subckt lablb1 VDD QN Q GND RN D SN GN
M1 N_6 SN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_22 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_22 RN N_21 GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_4 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 N_24 RN N_23 GND mn5  l=0.5u w=0.5u m=1
M10 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M11 Q N_7 GND GND mn5  l=0.5u w=0.58u m=1
M12 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_6 N_14 VDD mp5  l=0.42u w=0.52u m=1
M15 N_6 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_5 N_13 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_7 N_6 N_16 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 Q N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lablb1
* SPICE INPUT		Wed Jul 10 13:40:48 2019	lablb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb2
.subckt lablb2 VDD QN Q GND RN D SN GN
M1 N_6 SN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_22 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_22 RN N_21 GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_4 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 N_24 RN N_23 GND mn5  l=0.5u w=0.5u m=1
M10 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M11 Q N_7 GND GND mn5  l=0.5u w=0.72u m=1
M12 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_6 N_14 VDD mp5  l=0.42u w=0.52u m=1
M15 N_6 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_5 N_13 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_7 N_6 N_16 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 Q N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lablb2
* SPICE INPUT		Wed Jul 10 13:40:55 2019	lachb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb1
.subckt lachb1 RN D G GND QN Q VDD
M1 N_5 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_3 GND mn5  l=0.5u w=0.5u m=1
M6 N_21 RN N_20 GND mn5  l=0.5u w=0.5u m=1
M7 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_3 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_20 N_7 N_3 GND mn5  l=0.5u w=0.5u m=1
M11 N_21 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_7 G VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_3 N_7 N_31 VDD mp5  l=0.42u w=0.52u m=1
M16 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_32 N_5 N_3 VDD mp5  l=0.42u w=0.52u m=1
M18 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M19 Q N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_32 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lachb1
* SPICE INPUT		Wed Jul 10 13:41:02 2019	lachb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb2
.subckt lachb2 RN D G GND QN Q VDD
M1 N_5 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_3 GND mn5  l=0.5u w=0.5u m=1
M6 N_21 RN N_20 GND mn5  l=0.5u w=0.5u m=1
M7 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_3 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_20 N_7 N_3 GND mn5  l=0.5u w=0.5u m=1
M11 N_21 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_7 G VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_3 N_7 N_31 VDD mp5  l=0.42u w=0.52u m=1
M16 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_32 N_5 N_3 VDD mp5  l=0.42u w=0.52u m=1
M18 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 Q N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_32 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lachb2
* SPICE INPUT		Wed Jul 10 13:41:10 2019	lachq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachq1
.subckt lachq1 RN D G VDD GND Q
M1 N_3 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_6 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_16 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_17 RN N_16 GND mn5  l=0.5u w=0.5u m=1
M5 N_2 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_4 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_17 N_3 N_4 GND mn5  l=0.5u w=0.5u m=1
M8 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M9 N_18 N_6 N_4 GND mn5  l=0.5u w=0.5u m=1
M10 N_19 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_3 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 G VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 D VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_4 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M15 N_4 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M16 Q N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_29 N_3 N_4 VDD mp5  l=0.42u w=0.52u m=1
M19 N_29 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lachq1
* SPICE INPUT		Wed Jul 10 13:41:17 2019	lachq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachq2
.subckt lachq2 RN D G VDD GND Q
M1 N_3 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_6 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_16 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_17 RN N_16 GND mn5  l=0.5u w=0.5u m=1
M5 N_2 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_4 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_17 N_3 N_4 GND mn5  l=0.5u w=0.5u m=1
M8 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M9 N_18 N_6 N_4 GND mn5  l=0.5u w=0.5u m=1
M10 N_19 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_3 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 G VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 D VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_4 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M15 N_4 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M16 Q N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M17 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_29 N_3 N_4 VDD mp5  l=0.42u w=0.52u m=1
M19 N_29 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lachq2
* SPICE INPUT		Wed Jul 10 13:41:24 2019	laclb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb1
.subckt laclb1 RN D GN GND QN Q VDD
M1 N_7 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_3 GND mn5  l=0.5u w=0.5u m=1
M6 N_21 RN N_20 GND mn5  l=0.5u w=0.5u m=1
M7 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_3 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_20 N_7 N_3 GND mn5  l=0.5u w=0.5u m=1
M11 N_21 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_5 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_3 N_7 N_31 VDD mp5  l=0.42u w=0.52u m=1
M16 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_32 N_5 N_3 VDD mp5  l=0.42u w=0.52u m=1
M18 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M19 Q N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_32 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends laclb1
* SPICE INPUT		Wed Jul 10 13:41:31 2019	laclb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb2
.subckt laclb2 RN D GN GND QN Q VDD
M1 N_7 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_3 GND mn5  l=0.5u w=0.5u m=1
M6 N_21 RN N_20 GND mn5  l=0.5u w=0.5u m=1
M7 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_3 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_20 N_7 N_3 GND mn5  l=0.5u w=0.5u m=1
M11 N_21 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_5 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_3 N_7 N_31 VDD mp5  l=0.42u w=0.52u m=1
M16 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_32 N_5 N_3 VDD mp5  l=0.42u w=0.52u m=1
M18 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 Q N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_32 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends laclb2
* SPICE INPUT		Wed Jul 10 13:41:39 2019	laclq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclq1
.subckt laclq1 GN D RN VDD Q GND
M1 N_6 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_16 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 RN N_16 GND mn5  l=0.5u w=0.5u m=1
M7 N_19 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_2 GN GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_2 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_8 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M13 N_6 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_28 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_29 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_2 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_3 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_8 N_3 N_28 VDD mp5  l=0.42u w=0.52u m=1
M19 N_29 N_2 N_8 VDD mp5  l=0.42u w=0.52u m=1
.ends laclq1
* SPICE INPUT		Wed Jul 10 13:41:46 2019	laclq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclq2
.subckt laclq2 GN D RN VDD Q GND
M1 N_6 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_16 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 RN N_16 GND mn5  l=0.5u w=0.5u m=1
M7 N_19 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_2 GN GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_2 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_8 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 N_6 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_28 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_29 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_2 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_3 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_8 N_3 N_28 VDD mp5  l=0.42u w=0.52u m=1
M19 N_29 N_2 N_8 VDD mp5  l=0.42u w=0.52u m=1
.ends laclq2
* SPICE INPUT		Wed Jul 10 13:41:53 2019	lanhb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb1
.subckt lanhb1 D G GND QN Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_5 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_16 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_25 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_5 N_4 N_25 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 Q N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M18 N_26 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhb1
* SPICE INPUT		Wed Jul 10 13:42:00 2019	lanhb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb2
.subckt lanhb2 D G GND QN Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_5 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_16 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_25 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_5 N_4 N_25 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 Q N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M18 N_26 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhb2
* SPICE INPUT		Wed Jul 10 13:42:07 2019	lanhn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhn1
.subckt lanhn1 D G GND QN VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhn1
* SPICE INPUT		Wed Jul 10 13:42:14 2019	lanhn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhn2
.subckt lanhn2 D G GND QN VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhn2
* SPICE INPUT		Wed Jul 10 13:42:21 2019	lanhq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhq1
.subckt lanhq1 D G GND Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhq1
* SPICE INPUT		Wed Jul 10 13:42:29 2019	lanhq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhq2
.subckt lanhq2 D G GND Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhq2
* SPICE INPUT		Wed Jul 10 13:42:36 2019	lanht1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanht1
.subckt lanht1 GND Q VDD OE D G
M1 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 N_6 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_12 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_11 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q OE N_8 GND mn5  l=0.5u w=0.58u m=1
M10 N_3 OE GND GND mn5  l=0.5u w=0.5u m=1
M11 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_25 D VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 N_4 N_25 VDD mp5  l=0.42u w=0.52u m=1
M15 N_8 N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_26 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Q N_3 N_8 VDD mp5  l=0.42u w=0.76u m=1
M20 N_3 OE VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanht1
* SPICE INPUT		Wed Jul 10 13:42:43 2019	lanht2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanht2
.subckt lanht2 GND Q VDD OE D G
M1 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 N_6 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_12 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_11 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q OE N_8 GND mn5  l=0.5u w=0.72u m=1
M10 N_3 OE GND GND mn5  l=0.5u w=0.5u m=1
M11 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_25 D VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 N_4 N_25 VDD mp5  l=0.42u w=0.52u m=1
M15 N_8 N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_26 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Q N_3 N_8 VDD mp5  l=0.42u w=0.96u m=1
M20 N_3 OE VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanht2
* SPICE INPUT		Wed Jul 10 13:42:50 2019	lanlb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb1
.subckt lanlb1 GND QN Q VDD D GN
M1 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_7 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_6 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_11 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_10 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_6 N_5 N_22 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 Q N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_23 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_23 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlb1
* SPICE INPUT		Wed Jul 10 13:42:57 2019	lanlb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb2
.subckt lanlb2 GND QN Q VDD D GN
M1 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_7 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_6 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_11 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_10 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_6 N_5 N_22 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 Q N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_23 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_23 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlb2
* SPICE INPUT		Wed Jul 10 13:43:04 2019	lanln1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanln1
.subckt lanln1 D GN GND QN VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanln1
* SPICE INPUT		Wed Jul 10 13:43:11 2019	lanln2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanln2
.subckt lanln2 D GN GND QN VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanln2
* SPICE INPUT		Wed Jul 10 13:43:19 2019	lanlq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlq1
.subckt lanlq1 D GN GND Q VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlq1
* SPICE INPUT		Wed Jul 10 13:43:26 2019	lanlq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlq2
.subckt lanlq2 D GN GND Q VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlq2
* SPICE INPUT		Wed Jul 10 13:43:33 2019	laphb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb1
.subckt laphb1 GND QN Q VDD D SN G
M1 N_7 N_5 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M9 Q N_7 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 D VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_7 N_4 N_27 VDD mp5  l=0.42u w=0.52u m=1
M19 N_27 N_6 N_26 VDD mp5  l=0.42u w=0.52u m=1
M20 N_29 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends laphb1
* SPICE INPUT		Wed Jul 10 13:43:40 2019	laphb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb2
.subckt laphb2 GND QN Q VDD D SN G
M1 N_7 N_5 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M9 Q N_7 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 D VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_7 N_4 N_27 VDD mp5  l=0.42u w=0.52u m=1
M19 N_27 N_6 N_26 VDD mp5  l=0.42u w=0.52u m=1
M20 N_29 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M22 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends laphb2
* SPICE INPUT		Wed Jul 10 13:43:47 2019	laplb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb1
.subckt laplb1 GND QN Q VDD D SN GN
M1 N_7 N_4 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M9 Q N_7 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 D VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_7 N_5 N_27 VDD mp5  l=0.42u w=0.52u m=1
M19 N_27 N_6 N_26 VDD mp5  l=0.42u w=0.52u m=1
M20 N_29 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends laplb1
* SPICE INPUT		Wed Jul 10 13:43:55 2019	laplb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb2
.subckt laplb2 GND QN Q VDD D SN GN
M1 N_7 N_4 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M9 Q N_7 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 D VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_7 N_5 N_27 VDD mp5  l=0.42u w=0.52u m=1
M19 N_27 N_6 N_26 VDD mp5  l=0.42u w=0.52u m=1
M20 N_29 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M22 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends laplb2
* SPICE INPUT		Wed Jul 10 13:44:02 2019	mi02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR



* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad1
.subckt tlatncad1 VDD ECK GND CK E
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_21 E GND GND mn5  l=0.5u w=0.5u m=1
M3 N_21 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_22 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_22 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 ECK N_5 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_6 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_3 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_9 E VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_10 N_3 N_5 VDD mp5  l=0.42u w=0.5u m=1
M13 N_9 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M14 N_10 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M15 N_11 N_5 ECK VDD mp5  l=0.42u w=0.76u m=1
M16 N_6 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_11 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends tlatncad1
* SPICE INPUT		Wed Jul 10 14:04:29 2019	tlatncad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad2
.subckt tlatncad2 VDD ECK GND CK E
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_21 E GND GND mn5  l=0.5u w=0.5u m=1
M3 N_21 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_22 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_22 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 ECK N_5 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_6 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M8 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M9 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M10 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_9 E VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_10 N_3 N_5 VDD mp5  l=0.42u w=0.5u m=1
M13 N_9 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M14 N_10 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M15 N_11 N_5 ECK VDD mp5  l=0.42u w=0.96u m=1
M16 N_6 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_11 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends tlatncad2
* SPICE INPUT		Wed Jul 10 14:04:36 2019	tlatncad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad4
.subckt tlatncad4 GND ECK VDD E CK
M1 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 ECK N_5 GND GND mn5  l=0.5u w=0.72u m=1
M5 ECK N_5 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_10 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M10 N_10 E GND GND mn5  l=0.5u w=0.5u m=1
M11 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_6 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_28 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_27 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M18 N_28 N_3 N_5 VDD mp5  l=0.42u w=0.5u m=1
M19 N_27 E VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_15 N_5 ECK VDD mp5  l=0.42u w=0.96u m=1
M22 ECK N_5 N_15 VDD mp5  l=0.42u w=0.96u m=1
.ends tlatncad4
* SPICE INPUT		Wed Jul 10 14:04:43 2019	tlatntscad1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad1
.subckt tlatntscad1 VDD ECK GND CK SE E
M1 N_4 E GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 SE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_27 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M7 N_28 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_28 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_7 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_8 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 ECK N_3 GND GND mn5  l=0.5u w=0.58u m=1
M12 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M13 N_11 E N_4 VDD mp5  l=0.42u w=0.52u m=1
M14 N_11 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_6 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_12 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_13 N_3 N_7 VDD mp5  l=0.42u w=0.5u m=1
M19 N_12 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_7 ECK VDD mp5  l=0.42u w=0.76u m=1
M22 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M24 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends tlatntscad1
* SPICE INPUT		Wed Jul 10 14:04:51 2019	tlatntscad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad2
.subckt tlatntscad2 VDD ECK GND CK SE E
M1 N_4 E GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 SE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_28 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_29 N_6 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_8 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M11 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M12 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M13 N_12 E N_4 VDD mp5  l=0.42u w=0.52u m=1
M14 N_12 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 VDD N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M17 N_13 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_14 N_3 N_8 VDD mp5  l=0.42u w=0.5u m=1
M19 N_13 N_6 N_8 VDD mp5  l=0.42u w=0.52u m=1
M20 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_15 N_8 ECK VDD mp5  l=0.42u w=0.96u m=1
M22 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M24 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends tlatntscad2
* SPICE INPUT		Wed Jul 10 14:04:58 2019	tlatntscad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad4
.subckt tlatntscad4 GND ECK VDD CK SE E
M1 N_4 E GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 SE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_12 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_7 GND GND mn5  l=0.5u w=0.72u m=1
M10 ECK N_7 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_8 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M13 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M14 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M15 ECK N_7 N_15 VDD mp5  l=0.42u w=0.96u m=1
M16 ECK N_7 N_15 VDD mp5  l=0.42u w=0.96u m=1
M17 N_33 E N_4 VDD mp5  l=0.42u w=0.52u m=1
M18 N_33 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 VDD N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M21 N_34 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_35 N_3 N_7 VDD mp5  l=0.42u w=0.5u m=1
M23 N_34 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M24 N_35 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends tlatntscad4
* SPICE INPUT		Wed Jul 10 14:05:05 2019	xn02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR



***********************************************************

* SPICE INPUT		Wed Jul 10 13:34:20 2019	dfbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb1
.subckt dfbfb1 VDD QN Q GND RN SN CKN D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_26 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_6 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CKN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_6 N_28 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M18 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_6 N_5 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_4 N_5 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_4 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_6 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M38 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfbfb1
* SPICE INPUT		Wed Jul 10 13:34:27 2019	dfbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb2
.subckt dfbfb2 VDD QN Q GND RN SN CKN D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_26 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_6 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CKN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_6 N_28 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M20 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_6 N_5 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_4 N_5 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_4 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_6 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M40 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfbfb2
* SPICE INPUT		Wed Jul 10 13:34:34 2019	dfbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb1
.subckt dfbrb1 VDD QN Q GND RN SN CK D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_6 N_26 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CK GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_6 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_8 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M13 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M14 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M17 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_6 N_5 VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_6 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M34 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M37 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfbrb1
* SPICE INPUT		Wed Jul 10 13:34:42 2019	dfbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb2
.subckt dfbrb2 VDD QN Q GND RN SN CK D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_6 N_26 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CK GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_6 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_8 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M20 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_6 N_5 VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_6 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M40 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfbrb2
* SPICE INPUT		Wed Jul 10 13:34:49 2019	dfbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq1
.subckt dfbrq1 VDD Q GND RN D SN CK
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 SN GND GND mn5  l=0.5u w=0.58u m=1
M3 N_26 N_3 Q GND mn5  l=0.5u w=0.58u m=1
M4 N_26 N_8 Q GND mn5  l=0.5u w=0.58u m=1
M5 N_25 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_3 N_25 GND mn5  l=0.5u w=0.5u m=1
M7 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_5 N_30 GND mn5  l=0.5u w=0.5u m=1
M10 N_31 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M13 N_21 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_21 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_29 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M17 N_6 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M18 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M21 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M23 Q N_3 N_18 VDD mp5  l=0.42u w=0.76u m=1
M24 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_18 N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.5u m=1
M27 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M31 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M34 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M36 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M37 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M38 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfbrq1
* SPICE INPUT		Wed Jul 10 13:34:56 2019	dfbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq2
.subckt dfbrq2 VDD Q GND SN D RN CK
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_24 SN GND GND mn5  l=0.5u w=0.72u m=1
M6 N_24 N_3 Q GND mn5  l=0.5u w=0.72u m=1
M7 Q N_8 N_24 GND mn5  l=0.5u w=0.72u m=1
M8 N_23 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_3 N_23 GND mn5  l=0.5u w=0.5u m=1
M10 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M11 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_8 N_5 N_30 GND mn5  l=0.5u w=0.5u m=1
M13 N_31 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M14 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_19 SN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_19 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_19 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M18 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_29 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M20 N_6 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M21 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M26 Q N_3 N_18 VDD mp5  l=0.42u w=0.96u m=1
M27 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_18 N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.5u m=1
M30 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M34 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M40 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
.ends dfbrq2
* SPICE INPUT		Wed Jul 10 13:35:03 2019	dfcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb1
.subckt dfcfb1 GND QN Q VDD RN D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_14 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_15 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_8 N_4 N_16 GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M18 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M19 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_22 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M23 N_21 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M24 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M29 N_25 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M33 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M36 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfcfb1
* SPICE INPUT		Wed Jul 10 13:35:11 2019	dfcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb2
.subckt dfcfb2 GND QN Q VDD RN D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_14 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_15 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_8 N_4 N_16 GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M18 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M19 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_22 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M23 N_21 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M24 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M29 N_25 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M33 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M36 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfcfb2
* SPICE INPUT		Wed Jul 10 13:35:18 2019	dfcfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfq1
.subckt dfcfq1 GND Q VDD CKN D RN
M1 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_16 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_16 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_15 GND mn5  l=0.5u w=0.5u m=1
M9 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_14 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_13 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_25 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_24 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 N_24 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_25 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_23 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_22 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_22 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_21 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_20 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_20 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcfq1
* SPICE INPUT		Wed Jul 10 13:35:25 2019	dfcfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfq2
.subckt dfcfq2 GND Q VDD CKN D RN
M1 N_16 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_16 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 N_4 N_15 GND mn5  l=0.5u w=0.5u m=1
M5 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M7 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_14 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_13 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_35 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_35 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_34 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M21 N_36 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M22 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M24 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M25 N_34 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_33 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_33 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_32 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_31 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M30 N_32 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M31 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_36 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfcfq2
* SPICE INPUT		Wed Jul 10 13:35:32 2019	dfcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb1
.subckt dfcrb1 VDD QN Q GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_26 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_26 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M10 N_25 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_24 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_24 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_23 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_23 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M27 N_17 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_14 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M33 N_15 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M34 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrb1
* SPICE INPUT		Wed Jul 10 13:35:39 2019	dfcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb2
.subckt dfcrb2 GND QN Q VDD CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_17 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_5 N_16 GND mn5  l=0.5u w=0.5u m=1
M10 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_25 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M27 N_24 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_21 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M33 N_22 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M34 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrb2
* SPICE INPUT		Wed Jul 10 13:35:47 2019	dfcrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrn1
.subckt dfcrn1 VDD QN GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_34 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_34 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_33 GND mn5  l=0.5u w=0.5u m=1
M8 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_17 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrn1
* SPICE INPUT		Wed Jul 10 13:35:54 2019	dfcrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrn2
.subckt dfcrn2 VDD QN GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_23 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_22 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_22 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_21 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_21 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_17 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrn2
* SPICE INPUT		Wed Jul 10 13:36:01 2019	dfcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq1
.subckt dfcrq1 VDD Q GND CK D RN
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 Q N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_9 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_18 N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.52u m=1
M21 N_18 N_3 Q VDD mp5  l=0.42u w=0.76u m=1
M22 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrq1
* SPICE INPUT		Wed Jul 10 13:36:08 2019	dfcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq2
.subckt dfcrq2 VDD Q GND RN D CK
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_18 N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_18 N_3 Q VDD mp5  l=0.42u w=0.96u m=1
M21 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrq2
* SPICE INPUT		Wed Jul 10 13:36:15 2019	dfnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb1
.subckt dfnfb1 VDD QN Q GND D CKN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_5 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnfb1
* SPICE INPUT		Wed Jul 10 13:36:22 2019	dfnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb2
.subckt dfnfb2 VDD QN Q GND CKN D
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_5 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M15 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M18 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfnfb2
* SPICE INPUT		Wed Jul 10 13:36:30 2019	dfnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb1
.subckt dfnrb1 VDD QN Q GND CK D
M1 QN N_10 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_10 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_32 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_31 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_30 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M11 N_6 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_10 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_10 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 VDD N_10 N_16 VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M20 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M21 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M25 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M26 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfnrb1
* SPICE INPUT		Wed Jul 10 13:36:37 2019	dfnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb2
.subckt dfnrb2 VDD QN Q GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M17 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfnrb2
* SPICE INPUT		Wed Jul 10 13:36:44 2019	dfnrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrn1
.subckt dfnrn1 VDD QN GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrn1
* SPICE INPUT		Wed Jul 10 13:36:51 2019	dfnrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrn2
.subckt dfnrn2 VDD QN GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrn2
* SPICE INPUT		Wed Jul 10 13:36:58 2019	dfnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq1
.subckt dfnrq1 VDD Q GND CK D
M1 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrq1
* SPICE INPUT		Wed Jul 10 13:37:05 2019	dfnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq2
.subckt dfnrq2 VDD Q GND CK D
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrq2
* SPICE INPUT		Wed Jul 10 13:37:13 2019	dfpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb1
.subckt dfpfb1 VDD Q QN GND CKN D SN
M1 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_36 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_36 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_33 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_33 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfpfb1
* SPICE INPUT		Wed Jul 10 13:37:20 2019	dfpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb2
.subckt dfpfb2 VDD Q QN GND CKN D SN
M1 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_36 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_36 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M10 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_33 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M32 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M33 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfpfb2
* SPICE INPUT		Wed Jul 10 13:37:27 2019	dfprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb1
.subckt dfprb1 VDD Q QN GND SN D CK
M1 N_4 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_33 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_33 N_12 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_34 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_34 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_10 GND GND mn5  l=0.5u w=0.58u m=1
M7 QN N_8 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_10 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_35 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_35 SN N_6 GND mn5  l=0.5u w=0.5u m=1
M11 N_38 N_7 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_36 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_4 N_36 GND mn5  l=0.5u w=0.5u m=1
M14 N_37 N_12 N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_37 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_38 SN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_12 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_4 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_15 N_12 N_5 VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 Q N_10 VDD VDD mp5  l=0.42u w=0.76u m=1
M24 QN N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M25 N_10 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_6 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_6 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_12 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_17 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M32 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_8 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_12 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprb1
* SPICE INPUT		Wed Jul 10 13:37:34 2019	dfprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb2
.subckt dfprb2 VDD Q QN GND SN D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_34 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_34 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M10 N_35 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_4 N_35 GND mn5  l=0.5u w=0.5u m=1
M12 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M13 N_36 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M14 N_36 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_37 SN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_37 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_4 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_7 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_7 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M30 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M32 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfprb2
* SPICE INPUT		Wed Jul 10 13:37:41 2019	dfprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq1
.subckt dfprq1 VDD Q GND CK D SN
M1 Q N_8 N_27 GND mn5  l=0.5u w=0.58u m=1
M2 N_27 SN GND GND mn5  l=0.5u w=0.58u m=1
M3 N_33 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 N_33 GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_32 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_31 GND mn5  l=0.5u w=0.5u m=1
M8 N_31 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_30 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_30 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M19 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_9 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_14 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_7 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_7 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_11 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprq1
* SPICE INPUT		Wed Jul 10 13:37:48 2019	dfprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq2
.subckt dfprq2 VDD Q GND CK D SN
M1 Q N_10 N_29 GND mn5  l=0.5u w=0.72u m=1
M2 N_29 SN GND GND mn5  l=0.5u w=0.72u m=1
M3 N_35 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_34 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 N_10 N_35 GND mn5  l=0.5u w=0.5u m=1
M6 N_34 N_5 N_10 GND mn5  l=0.5u w=0.5u m=1
M7 N_10 N_4 N_33 GND mn5  l=0.5u w=0.5u m=1
M8 N_33 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_32 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_32 N_7 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M13 N_30 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_30 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_11 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_16 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_11 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_15 N_5 N_10 VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_9 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_13 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_5 N_7 VDD mp5  l=0.42u w=0.5u m=1
M29 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_4 N_10 VDD mp5  l=0.42u w=0.5u m=1
M31 VDD N_5 N_4 VDD mp5  l=0.42u w=0.5u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprq2


***********************************************************

* SPICE INPUT		Wed Jul 10 14:00:28 2019	sdbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb1
.subckt sdbfb1 VDD Q QN GND RN SN SI SE D CKN
M1 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M9 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M10 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M11 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_9 N_5 N_29 GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_4 N_55 GND mn5  l=0.5u w=0.5u m=1
M14 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M16 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M17 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_4 N_56 GND mn5  l=0.5u w=0.5u m=1
M20 N_57 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M21 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M23 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M24 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M25 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M26 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M28 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_4 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M34 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M44 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M45 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M46 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M47 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M48 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdbfb1
* SPICE INPUT		Wed Jul 10 14:00:35 2019	sdbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb2
.subckt sdbfb2 VDD Q QN GND RN SN SI SE D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_5 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_4 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_4 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M20 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M21 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M22 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M23 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M24 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M25 N_4 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.52u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M42 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M44 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M45 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M46 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M47 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M48 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdbfb2
* SPICE INPUT		Wed Jul 10 14:00:42 2019	sdbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb1
.subckt sdbrb1 VDD Q QN GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M18 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M19 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M20 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M21 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M22 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M23 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M24 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M42 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M44 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M45 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M46 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M47 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M48 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdbrb1
* SPICE INPUT		Wed Jul 10 14:00:50 2019	sdbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb2
.subckt sdbrb2 VDD Q QN GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M18 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M20 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M21 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M22 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M23 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M24 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M43 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M44 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M45 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M46 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M47 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M48 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
.ends sdbrb2
* SPICE INPUT		Wed Jul 10 14:00:57 2019	sdbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq1
.subckt sdbrq1 VDD Q GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_35 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_35 N_6 N_30 GND mn5  l=0.5u w=0.5u m=1
M6 N_36 SI N_30 GND mn5  l=0.5u w=0.5u m=1
M7 N_36 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_30 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_37 GND mn5  l=0.5u w=0.5u m=1
M10 N_37 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_28 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_28 N_3 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_38 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_38 GND mn5  l=0.5u w=0.5u m=1
M16 Q N_11 N_24 GND mn5  l=0.5u w=0.58u m=1
M17 N_24 N_3 Q GND mn5  l=0.5u w=0.58u m=1
M18 N_24 SN GND GND mn5  l=0.5u w=0.58u m=1
M19 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M20 N_39 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M21 N_39 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_12 N_3 N_26 GND mn5  l=0.5u w=0.5u m=1
M23 N_26 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M24 N_26 SN GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_22 N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M42 Q N_3 N_22 VDD mp5  l=0.42u w=0.76u m=1
M43 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M44 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M45 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M46 N_21 N_3 N_12 VDD mp5  l=0.42u w=0.5u m=1
M47 N_21 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M48 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdbrq1
* SPICE INPUT		Wed Jul 10 14:01:05 2019	sdbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq2
.subckt sdbrq2 VDD Q GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_35 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_35 N_6 N_30 GND mn5  l=0.5u w=0.5u m=1
M6 N_36 SI N_30 GND mn5  l=0.5u w=0.5u m=1
M7 N_36 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_30 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_37 GND mn5  l=0.5u w=0.5u m=1
M10 N_37 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_28 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_28 N_3 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_38 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_12 N_3 N_26 GND mn5  l=0.5u w=0.5u m=1
M16 N_26 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M17 N_26 SN GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 N_24 GND mn5  l=0.5u w=0.72u m=1
M19 N_24 N_3 Q GND mn5  l=0.5u w=0.72u m=1
M20 N_24 SN GND GND mn5  l=0.5u w=0.72u m=1
M21 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M22 N_11 N_5 N_38 GND mn5  l=0.5u w=0.5u m=1
M23 N_39 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M24 N_39 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_21 N_3 N_12 VDD mp5  l=0.42u w=0.5u m=1
M41 N_21 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M42 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M43 N_22 N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M44 Q N_3 N_22 VDD mp5  l=0.42u w=0.96u m=1
M45 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M46 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M47 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M48 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdbrq2
* SPICE INPUT		Wed Jul 10 14:01:12 2019	sdcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb1
.subckt sdcfb1 VDD Q QN GND RN SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_26 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M6 N_47 SI N_26 GND mn5  l=0.5u w=0.5u m=1
M7 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M9 N_48 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_11 N_5 N_49 GND mn5  l=0.5u w=0.5u m=1
M15 N_50 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M16 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M20 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M28 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M32 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M35 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M37 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M38 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M41 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M42 N_14 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M43 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M44 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends sdcfb1
* SPICE INPUT		Wed Jul 10 14:01:19 2019	sdcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb2
.subckt sdcfb2 VDD Q QN GND CKN D SE SI RN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M5 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M10 N_11 N_5 N_49 GND mn5  l=0.5u w=0.5u m=1
M11 N_50 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M12 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_28 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M14 N_47 SI N_28 GND mn5  l=0.5u w=0.5u m=1
M15 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M17 N_48 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 N_14 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M31 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M33 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M35 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M39 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M44 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdcfb2
* SPICE INPUT		Wed Jul 10 14:01:27 2019	sdcfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfq1
.subckt sdcfq1 VDD Q GND CKN D SE SI RN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_5 N_47 GND mn5  l=0.5u w=0.5u m=1
M4 N_48 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M6 N_48 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_44 D GND GND mn5  l=0.5u w=0.5u m=1
M10 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M11 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M13 N_27 N_6 N_44 GND mn5  l=0.5u w=0.5u m=1
M14 N_45 SI N_27 GND mn5  l=0.5u w=0.5u m=1
M15 N_45 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_4 N_27 GND mn5  l=0.5u w=0.5u m=1
M17 N_46 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_47 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M25 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_21 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_12 N_13 N_22 VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M33 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M38 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_10 N_13 N_19 VDD mp5  l=0.42u w=0.52u m=1
M41 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcfq1
* SPICE INPUT		Wed Jul 10 14:01:34 2019	sdcfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfq2
.subckt sdcfq2 VDD Q GND RN SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_48 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_48 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_44 D GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M12 N_25 N_6 N_44 GND mn5  l=0.5u w=0.5u m=1
M13 N_45 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M14 N_45 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M16 N_46 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_47 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_11 N_5 N_47 GND mn5  l=0.5u w=0.5u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_21 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_12 N_13 N_22 VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M30 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M37 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M38 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_10 N_13 N_19 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
.ends sdcfq2
* SPICE INPUT		Wed Jul 10 14:01:41 2019	sdcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb1
.subckt sdcrb1 VDD Q QN GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M5 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_50 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M13 N_11 N_4 N_49 GND mn5  l=0.5u w=0.5u m=1
M14 N_26 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M15 N_47 SI N_26 GND mn5  l=0.5u w=0.5u m=1
M16 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_5 N_26 GND mn5  l=0.5u w=0.5u m=1
M18 N_48 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M19 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M31 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M35 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M40 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M41 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M44 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrb1
* SPICE INPUT		Wed Jul 10 14:01:49 2019	sdcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb2
.subckt sdcrb2 VDD Q QN GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M5 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_50 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M13 N_11 N_4 N_49 GND mn5  l=0.5u w=0.5u m=1
M14 N_26 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M15 N_47 SI N_26 GND mn5  l=0.5u w=0.5u m=1
M16 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_5 N_26 GND mn5  l=0.5u w=0.5u m=1
M18 N_48 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M19 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M31 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M35 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M40 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M41 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M44 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrb2
* SPICE INPUT		Wed Jul 10 14:01:56 2019	sdcrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrn1
.subckt sdcrn1 VDD QN GND RN SI SE D CK
M1 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_42 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M9 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_24 N_6 N_42 GND mn5  l=0.5u w=0.5u m=1
M13 N_43 SI N_24 GND mn5  l=0.5u w=0.5u m=1
M14 N_43 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_5 N_24 GND mn5  l=0.5u w=0.5u m=1
M16 N_44 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_44 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M21 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M28 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_21 VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_10 N_13 N_18 VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrn1
* SPICE INPUT		Wed Jul 10 14:02:03 2019	sdcrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrn2
.subckt sdcrn2 VDD QN GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_42 D GND GND mn5  l=0.5u w=0.5u m=1
M5 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_24 N_6 N_42 GND mn5  l=0.5u w=0.5u m=1
M9 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M12 N_43 SI N_24 GND mn5  l=0.5u w=0.5u m=1
M13 N_43 SE GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_5 N_24 GND mn5  l=0.5u w=0.5u m=1
M15 N_44 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M16 N_44 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M26 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_12 N_13 N_21 VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_21 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M36 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 N_13 N_18 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
.ends sdcrn2
* SPICE INPUT		Wed Jul 10 14:02:11 2019	sdcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq1
.subckt sdcrq1 VDD Q GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_12 GND GND mn5  l=0.5u w=0.58u m=1
M4 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_13 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 RN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_47 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_43 D GND GND mn5  l=0.5u w=0.5u m=1
M10 N_47 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M11 N_11 N_4 N_46 GND mn5  l=0.5u w=0.5u m=1
M12 N_25 N_6 N_43 GND mn5  l=0.5u w=0.5u m=1
M13 N_44 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M14 N_44 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M16 N_45 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M24 Q N_12 N_15 VDD mp5  l=0.42u w=0.76u m=1
M25 N_15 N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_12 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_21 N_13 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M32 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M33 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M38 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_10 N_12 N_19 VDD mp5  l=0.42u w=0.52u m=1
M41 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_22 N_12 N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrq1
* SPICE INPUT		Wed Jul 10 14:02:18 2019	sdcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq2
.subckt sdcrq2 VDD Q GND RN SI SE D CK
M1 N_12 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M4 Q N_12 GND GND mn5  l=0.5u w=0.72u m=1
M5 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_13 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_47 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_43 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_47 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M12 N_11 N_4 N_46 GND mn5  l=0.5u w=0.5u m=1
M13 N_25 N_6 N_43 GND mn5  l=0.5u w=0.5u m=1
M14 N_44 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M15 N_44 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_45 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_12 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q N_12 N_15 VDD mp5  l=0.42u w=0.96u m=1
M26 N_15 N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_22 N_12 N_13 VDD mp5  l=0.42u w=0.52u m=1
M30 N_21 N_13 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M33 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M34 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M38 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M39 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 N_12 N_19 VDD mp5  l=0.42u w=0.52u m=1
M42 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrq2
* SPICE INPUT		Wed Jul 10 14:02:25 2019	sdnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb1
.subckt sdnfb1 GND QN Q VDD SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M6 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M7 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_17 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_11 N_5 N_18 GND mn5  l=0.5u w=0.5u m=1
M14 N_19 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M15 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M18 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M19 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M24 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M25 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_9 N_5 N_21 VDD mp5  l=0.42u w=0.52u m=1
M27 N_40 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M28 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_41 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M32 N_42 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M33 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M36 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends sdnfb1
* SPICE INPUT		Wed Jul 10 14:02:33 2019	sdnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb2
.subckt sdnfb2 GND QN Q VDD SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_19 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_5 N_18 GND mn5  l=0.5u w=0.5u m=1
M10 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M14 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_17 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M22 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M24 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_42 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_41 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M29 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M32 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M33 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_9 N_5 N_21 VDD mp5  l=0.42u w=0.52u m=1
M35 N_40 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M36 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdnfb2
* SPICE INPUT		Wed Jul 10 14:02:40 2019	sdnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb1
.subckt sdnrb1 GND QN Q VDD SI SE D CK
M1 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M3 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 N_4 N_18 GND mn5  l=0.5u w=0.5u m=1
M8 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M10 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M13 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M14 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M16 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M18 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M19 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_42 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M25 N_41 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M26 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M33 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M34 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_9 N_4 N_21 VDD mp5  l=0.42u w=0.52u m=1
M36 N_40 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
.ends sdnrb1
* SPICE INPUT		Wed Jul 10 14:02:47 2019	sdnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb2
.subckt sdnrb2 GND QN Q VDD SI SE D CK
M1 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_19 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 N_4 N_18 GND mn5  l=0.5u w=0.5u m=1
M6 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M8 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M14 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M19 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_42 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M23 N_41 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M24 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M31 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M32 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_9 N_4 N_21 VDD mp5  l=0.42u w=0.52u m=1
M34 N_40 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdnrb2
* SPICE INPUT		Wed Jul 10 14:02:54 2019	sdnrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrn1
.subckt sdnrn1 GND QN VDD SI SE D CK
M1 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M7 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M9 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M12 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M13 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M14 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M15 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M16 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M18 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M23 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M24 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_20 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_37 N_6 N_20 VDD mp5  l=0.42u w=0.52u m=1
M32 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_9 N_4 N_20 VDD mp5  l=0.42u w=0.52u m=1
M34 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
.ends sdnrn1
* SPICE INPUT		Wed Jul 10 14:03:02 2019	sdnrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrn2
.subckt sdnrn2 GND QN VDD CK D SE SI
M1 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M14 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M21 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M22 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M27 N_9 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M28 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_37 N_6 N_22 VDD mp5  l=0.42u w=0.52u m=1
M30 N_22 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdnrn2
* SPICE INPUT		Wed Jul 10 14:03:09 2019	sdnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq1
.subckt sdnrq1 GND Q VDD CK D SE SI
M1 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M2 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M10 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M12 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M13 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M14 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M19 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M20 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M24 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_9 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M26 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M29 N_37 N_6 N_22 VDD mp5  l=0.42u w=0.52u m=1
M30 N_22 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdnrq1
* SPICE INPUT		Wed Jul 10 14:03:16 2019	sdnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq2
.subckt sdnrq2 GND Q VDD CK D SE SI
M1 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M5 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M14 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M21 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M23 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M27 N_9 N_4 N_19 VDD mp5  l=0.42u w=0.52u m=1
M28 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_37 N_6 N_19 VDD mp5  l=0.42u w=0.52u m=1
M30 N_19 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdnrq2
* SPICE INPUT		Wed Jul 10 14:03:23 2019	sdpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb1
.subckt sdpfb1 VDD Q QN GND CKN D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.58u m=1
M2 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M5 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_46 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_5 N_45 GND mn5  l=0.5u w=0.5u m=1
M9 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M11 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_43 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M15 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M18 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.76u m=1
M23 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M25 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M29 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M30 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M38 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M39 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdpfb1
* SPICE INPUT		Wed Jul 10 14:03:31 2019	sdpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb2
.subckt sdpfb2 VDD Q QN GND CKN D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_46 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M5 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_5 N_45 GND mn5  l=0.5u w=0.5u m=1
M7 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M9 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M10 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_43 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M15 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M18 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.96u m=1
M23 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M28 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M32 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M38 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M39 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdpfb2
* SPICE INPUT		Wed Jul 10 14:03:38 2019	sdprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb1
.subckt sdprb1 VDD Q QN GND CK D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M5 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M10 N_43 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M12 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M13 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M15 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M18 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.76u m=1
M23 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M28 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M32 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M33 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M35 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M38 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M39 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprb1
* SPICE INPUT		Wed Jul 10 14:03:45 2019	sdprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb2
.subckt sdprb2 VDD Q QN GND CK D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M7 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M9 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_43 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M12 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M13 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M14 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M15 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M18 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.96u m=1
M23 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M28 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M32 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M33 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M35 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M36 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M38 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M39 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M41 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprb2
* SPICE INPUT		Wed Jul 10 14:03:53 2019	sdprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq1
.subckt sdprq1 VDD Q GND CK D SN SE SI
M1 N_43 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M2 N_43 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_42 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_44 SN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_41 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_4 N_42 GND mn5  l=0.5u w=0.5u m=1
M7 N_41 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_11 N_44 GND mn5  l=0.5u w=0.5u m=1
M9 Q N_11 N_37 GND mn5  l=0.5u w=0.58u m=1
M10 N_40 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_40 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M12 N_9 N_5 N_24 GND mn5  l=0.5u w=0.5u m=1
M13 N_37 SN GND GND mn5  l=0.5u w=0.58u m=1
M14 N_39 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_39 SI N_24 GND mn5  l=0.5u w=0.5u m=1
M16 N_24 N_6 N_38 GND mn5  l=0.5u w=0.5u m=1
M17 N_38 D GND GND mn5  l=0.5u w=0.5u m=1
M18 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M19 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M20 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_18 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_17 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M23 N_17 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_18 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M29 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_16 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_16 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M32 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M33 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M34 N_15 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_15 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_7 SE N_14 VDD mp5  l=0.42u w=0.5u m=1
M37 N_14 D VDD VDD mp5  l=0.42u w=0.5u m=1
M38 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprq1
* SPICE INPUT		Wed Jul 10 14:04:00 2019	sdprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq2
.subckt sdprq2 GND Q VDD CK D SE SI SN
M1 N_20 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_20 N_4 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 N_3 N_19 GND mn5  l=0.5u w=0.5u m=1
M4 N_19 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_18 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_18 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 Q N_10 N_14 GND mn5  l=0.5u w=0.72u m=1
M10 N_17 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M12 N_14 SN GND GND mn5  l=0.5u w=0.72u m=1
M13 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M14 N_16 SI N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_6 N_5 N_15 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 SE GND GND mn5  l=0.5u w=0.5u m=1
M19 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M20 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_44 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_44 N_3 N_10 VDD mp5  l=0.42u w=0.5u m=1
M23 N_43 N_4 N_10 VDD mp5  l=0.42u w=0.52u m=1
M24 N_43 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_9 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_42 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 Q N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_11 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_42 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M31 N_8 N_3 N_25 VDD mp5  l=0.42u w=0.5u m=1
M32 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M33 N_41 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_41 N_5 N_25 VDD mp5  l=0.42u w=0.5u m=1
M35 N_11 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M36 N_25 SE N_40 VDD mp5  l=0.42u w=0.5u m=1
M37 N_40 D VDD VDD mp5  l=0.42u w=0.5u m=1
M38 N_5 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprq2


