* SPICE INPUT		Tue Jan 14 09:25:35 2020	buftld4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld4
.subckt buftld4 OE A GND Y VDD
M1 GND N_5 Y GND mn5  l=0.5u w=0.72u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_5 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M7 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M8 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 N_2 N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld4
* SPICE INPUT		Tue Jan 14 09:25:40 2020	buftld6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld6
.subckt buftld6 A OE VDD GND Y
M1 N_4 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M8 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M11 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_6 N_4 N_3 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld6
* SPICE INPUT		Tue Jan 14 09:25:45 2020	buftld8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld8
.subckt buftld8 OE A Y VDD GND
M1 GND N_5 Y GND mn5  l=0.5u w=0.72u m=1
M2 GND N_5 Y GND mn5  l=0.5u w=0.72u m=1
M3 GND N_5 Y GND mn5  l=0.5u w=0.72u m=1
M4 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M6 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_5 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_5 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M10 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M11 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M12 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_6 N_2 N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld8
* SPICE INPUT		Wed Jul 10 13:23:44 2019	ad01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d0
.subckt ad01d0 GND S CO VDD B CI A
M1 N_4 N_15 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_3 CI N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_10 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_14 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_15 CI GND GND mn5  l=0.5u w=0.5u m=1
M11 CO N_14 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_10 N_9 N_3 GND mn5  l=0.5u w=0.5u m=1
M13 S N_2 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_10 N_3 GND mn5  l=0.5u w=0.5u m=1
M15 N_3 N_15 N_2 VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 CI N_2 VDD mp5  l=0.42u w=0.52u m=1
M17 N_10 A VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_3 N_7 N_10 VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_7 N_10 N_3 VDD mp5  l=0.42u w=0.52u m=1
M21 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_4 N_14 VDD mp5  l=0.42u w=0.52u m=1
M23 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 CI VDD VDD mp5  l=0.42u w=0.52u m=1
M25 CO N_14 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_4 N_9 N_10 VDD mp5  l=0.42u w=0.52u m=1
M27 S N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
.ends ad01d0
* SPICE INPUT		Wed Jul 10 13:23:52 2019	ad01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d1
.subckt ad01d1 VDD S CO GND A B CI
M1 N_4 N_15 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_3 CI N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_9 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_14 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_15 CI GND GND mn5  l=0.5u w=0.5u m=1
M11 CO N_14 GND GND mn5  l=0.5u w=0.58u m=1
M12 N_9 N_8 N_3 GND mn5  l=0.5u w=0.5u m=1
M13 S N_2 GND GND mn5  l=0.5u w=0.58u m=1
M14 N_8 N_9 N_3 GND mn5  l=0.5u w=0.5u m=1
M15 N_3 N_15 N_2 VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 CI N_2 VDD mp5  l=0.42u w=0.52u m=1
M17 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_3 N_7 N_9 VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_7 N_9 N_3 VDD mp5  l=0.42u w=0.52u m=1
M21 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_4 N_14 VDD mp5  l=0.42u w=0.52u m=1
M23 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 CI VDD VDD mp5  l=0.42u w=0.52u m=1
M25 CO N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 N_4 N_8 N_9 VDD mp5  l=0.42u w=0.52u m=1
M27 S N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M28 N_4 N_9 N_8 VDD mp5  l=0.42u w=0.52u m=1
.ends ad01d1
* SPICE INPUT		Wed Jul 10 13:23:59 2019	ad01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d2
.subckt ad01d2 VDD S CO GND A B CI
M1 N_4 N_15 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_3 CI N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_9 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_14 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_15 CI GND GND mn5  l=0.5u w=0.5u m=1
M11 CO N_14 GND GND mn5  l=0.5u w=0.72u m=1
M12 N_9 N_8 N_3 GND mn5  l=0.5u w=0.5u m=1
M13 S N_2 GND GND mn5  l=0.5u w=0.72u m=1
M14 N_8 N_9 N_3 GND mn5  l=0.5u w=0.5u m=1
M15 N_3 N_15 N_2 VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 CI N_2 VDD mp5  l=0.42u w=0.52u m=1
M17 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_3 N_7 N_9 VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_7 N_9 N_3 VDD mp5  l=0.42u w=0.52u m=1
M21 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_4 N_14 VDD mp5  l=0.42u w=0.52u m=1
M23 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 CI VDD VDD mp5  l=0.42u w=0.52u m=1
M25 CO N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 N_4 N_8 N_9 VDD mp5  l=0.42u w=0.52u m=1
M27 S N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_4 N_9 N_8 VDD mp5  l=0.42u w=0.52u m=1
.ends ad01d2
* SPICE INPUT		Wed Jul 10 13:24:06 2019	ah01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d0
.subckt ah01d0 VDD CO S GND B A
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 S N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M3 GND A N_6 GND mn5  l=0.5u w=0.5u m=1
M4 CO N_8 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_21 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M7 S B N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_21 A N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 N_7 S VDD mp5  l=0.42u w=0.52u m=1
M11 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M12 CO N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M14 S B N_4 VDD mp5  l=0.42u w=0.52u m=1
M15 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_8 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ah01d0
* SPICE INPUT		Wed Jul 10 13:24:13 2019	ah01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d1
.subckt ah01d1 VDD CO S GND A B
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 S N_7 N_4 GND mn5  l=0.5u w=0.58u m=1
M3 GND A N_5 GND mn5  l=0.5u w=0.5u m=1
M4 S B N_5 GND mn5  l=0.5u w=0.58u m=1
M5 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_21 A N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_21 B GND GND mn5  l=0.5u w=0.5u m=1
M8 CO N_8 GND GND mn5  l=0.5u w=0.58u m=1
M9 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 S N_7 N_5 VDD mp5  l=0.42u w=0.76u m=1
M11 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M12 S B N_4 VDD mp5  l=0.42u w=0.76u m=1
M13 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_8 A VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M16 CO N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends ah01d1
* SPICE INPUT		Wed Jul 10 13:24:20 2019	ah01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d2
.subckt ah01d2 VDD CO S GND B A
M1 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M2 S N_4 N_5 GND mn5  l=0.5u w=0.72u m=1
M3 N_6 B S GND mn5  l=0.5u w=0.72u m=1
M4 N_6 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 A N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_12 B GND GND mn5  l=0.5u w=0.5u m=1
M7 CO N_8 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_5 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 S N_4 N_6 VDD mp5  l=0.42u w=0.96u m=1
M11 N_8 A VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M14 CO N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_5 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 S B N_5 VDD mp5  l=0.42u w=0.96u m=1
.ends ah01d2
* SPICE INPUT		Wed Jul 10 13:24:28 2019	an02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d0
.subckt an02d0 B A VDD Y GND
M1 N_8 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an02d0
* SPICE INPUT		Wed Jul 10 13:24:35 2019	an02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d1
.subckt an02d1 B A VDD Y GND
M1 N_8 A N_2 GND mn5  l=0.5u w=0.58u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.58u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an02d1
* SPICE INPUT		Wed Jul 10 13:24:42 2019	an02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d2
.subckt an02d2 B A VDD Y GND
M1 N_8 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends an02d2
* SPICE INPUT		Wed Jul 10 13:24:49 2019	an03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d0
.subckt an03d0 C B A GND Y VDD
M1 N_9 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 C VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an03d0
* SPICE INPUT		Wed Jul 10 13:24:56 2019	an03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d1
.subckt an03d1 C B A Y GND VDD
M1 N_9 A N_2 GND mn5  l=0.5u w=0.58u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.58u m=1
M3 N_10 C GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 C VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an03d1
* SPICE INPUT		Wed Jul 10 13:25:04 2019	an03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d2
.subckt an03d2 C B A Y GND VDD
M1 N_9 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 C VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends an03d2
* SPICE INPUT		Wed Jul 10 13:25:11 2019	an04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d0
.subckt an04d0 GND Y VDD D C B A
M1 N_6 A N_4 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.58u m=1
M3 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 D GND GND mn5  l=0.5u w=0.58u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 C VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 D VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an04d0
* SPICE INPUT		Wed Jul 10 13:25:18 2019	an04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d1
.subckt an04d1 GND Y VDD D C B A
M1 N_6 A N_4 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.58u m=1
M3 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 D GND GND mn5  l=0.5u w=0.58u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 C VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 D VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an04d1
* SPICE INPUT		Wed Jul 10 13:25:25 2019	an04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d2
.subckt an04d2 GND Y VDD A B C D
M1 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.58u m=1
M3 N_6 A N_4 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 D GND GND mn5  l=0.5u w=0.58u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 C VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 D VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends an04d2
* SPICE INPUT		Wed Jul 10 13:25:33 2019	an12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an12d0
.subckt an12d0 B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_14 N_4 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_14 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an12d0
* SPICE INPUT		Wed Jul 10 13:25:40 2019	an12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an12d1
.subckt an12d1 B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_14 N_4 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_14 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an12d1
* SPICE INPUT		Wed Jul 10 13:25:47 2019	an12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an12d2
.subckt an12d2 B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 N_4 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends an12d2
* SPICE INPUT		Wed Jul 10 13:25:54 2019	an13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an13d0
.subckt an13d0 C B AN GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an13d0
* SPICE INPUT		Wed Jul 10 13:26:01 2019	an13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an13d1
.subckt an13d1 C B AN VDD GND Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an13d1
* SPICE INPUT		Wed Jul 10 13:26:08 2019	an13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an13d2
.subckt an13d2 C B AN VDD GND Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an13d2
* SPICE INPUT		Wed Jul 10 13:26:15 2019	an23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an23d0
.subckt an23d0 C BN AN VDD Y GND
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_3 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_12 C GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_5 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an23d0
* SPICE INPUT		Wed Jul 10 13:26:23 2019	an23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an23d1
.subckt an23d1 C BN AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_5 N_2 GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_2 C VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an23d1
* SPICE INPUT		Wed Jul 10 13:26:30 2019	an23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an23d2
.subckt an23d2 C BN AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_3 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_12 C GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_6 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an23d2


* Top of hierarchy  cell=aoi211d0
.subckt aoi211d0 A0 A1 B0 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 Y A1 N_15 GND mn5  l=0.5u w=0.5u m=1
M4 N_15 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M6 N_6 B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M7 N_6 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi211d0
* SPICE INPUT		Wed Jul 10 13:26:51 2019	aoi211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d1
.subckt aoi211d1 A0 A1 B0 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.58u m=1
M2 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M3 Y A1 N_10 GND mn5  l=0.5u w=0.58u m=1
M4 N_10 A0 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y C0 N_16 VDD mp5  l=0.42u w=0.76u m=1
M6 N_6 B0 N_16 VDD mp5  l=0.42u w=0.76u m=1
M7 N_6 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_6 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aoi211d1
* SPICE INPUT		Wed Jul 10 13:26:58 2019	aoi211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d2
.subckt aoi211d2 A0 A1 B0 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A1 N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_10 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y C0 N_16 VDD mp5  l=0.42u w=0.96u m=1
M6 N_6 B0 N_16 VDD mp5  l=0.42u w=0.96u m=1
M7 N_6 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_6 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi211d2
* SPICE INPUT		Wed Jul 10 13:27:05 2019	aoi21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d0
.subckt aoi21d0 A0 A1 B0 GND Y VDD
M1 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_12 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y B0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M5 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi21d0
* SPICE INPUT		Wed Jul 10 13:27:13 2019	aoi21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d1
.subckt aoi21d1 A0 A1 B0 GND Y VDD
M1 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 A1 Y GND mn5  l=0.5u w=0.58u m=1
M3 N_9 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y B0 N_7 VDD mp5  l=0.42u w=0.76u m=1
M5 N_7 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 N_7 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aoi21d1
* SPICE INPUT		Wed Jul 10 13:27:20 2019	aoi21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d2
.subckt aoi21d2 A0 A1 B0 GND Y VDD
M1 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 A1 Y GND mn5  l=0.5u w=0.72u m=1
M3 N_9 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 N_7 VDD mp5  l=0.42u w=0.96u m=1
M5 N_7 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_7 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi21d2
* SPICE INPUT		Wed Jul 10 13:27:27 2019	aoi221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d0
.subckt aoi221d0 C0 A0 A1 B1 B0 VDD GND Y
M1 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B1 N_12 GND mn5  l=0.5u w=0.5u m=1
M3 N_13 A1 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_13 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y C0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_11 A1 N_7 VDD mp5  l=0.42u w=0.52u m=1
M10 N_11 A0 N_7 VDD mp5  l=0.42u w=0.52u m=1
.ends aoi221d0
* SPICE INPUT		Wed Jul 10 13:27:34 2019	aoi221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d1
.subckt aoi221d1 B0 A0 A1 B1 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.58u m=1
M2 Y B1 N_12 GND mn5  l=0.5u w=0.58u m=1
M3 N_13 A1 Y GND mn5  l=0.5u w=0.58u m=1
M4 N_13 A0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.58u m=1
M6 Y C0 N_8 VDD mp5  l=0.42u w=0.76u m=1
M7 N_7 B1 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_7 A1 N_8 VDD mp5  l=0.42u w=0.76u m=1
M9 N_7 A0 N_8 VDD mp5  l=0.42u w=0.76u m=1
M10 N_7 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aoi221d1
* SPICE INPUT		Wed Jul 10 13:27:41 2019	aoi221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d2
.subckt aoi221d2 B0 A0 A1 B1 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y B1 N_12 GND mn5  l=0.5u w=0.72u m=1
M3 N_13 A1 Y GND mn5  l=0.5u w=0.72u m=1
M4 N_13 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y C0 N_8 VDD mp5  l=0.42u w=0.96u m=1
M7 N_7 B1 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_7 A1 N_8 VDD mp5  l=0.42u w=0.96u m=1
M9 N_7 A0 N_8 VDD mp5  l=0.42u w=0.96u m=1
M10 N_7 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi221d2
* SPICE INPUT		Wed Jul 10 13:27:49 2019	aoi22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d0
.subckt aoi22d0 B0 B1 A1 A0 GND VDD Y
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 Y B1 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_8 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_8 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 B0 Y VDD mp5  l=0.42u w=0.52u m=1
.ends aoi22d0
* SPICE INPUT		Wed Jul 10 13:27:56 2019	aoi22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d1
.subckt aoi22d1 B0 B1 A1 A0 Y VDD GND
M1 N_11 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 Y A1 N_11 GND mn5  l=0.5u w=0.58u m=1
M3 Y B1 N_10 GND mn5  l=0.5u w=0.58u m=1
M4 N_10 B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_6 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 N_6 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_6 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M8 N_6 B0 Y VDD mp5  l=0.42u w=0.76u m=1
.ends aoi22d1
* SPICE INPUT		Wed Jul 10 13:28:03 2019	aoi22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d2
.subckt aoi22d2 A0 A1 B0 B1 GND Y VDD
M1 Y B1 N_10 GND mn5  l=0.5u w=0.72u m=1
M2 N_10 B0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A1 N_11 GND mn5  l=0.5u w=0.72u m=1
M4 N_11 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_8 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M6 N_8 B0 Y VDD mp5  l=0.42u w=0.96u m=1
M7 N_8 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_8 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi22d2
* SPICE INPUT		Wed Jul 10 13:28:11 2019	aoi31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d0
.subckt aoi31d0 A0 A1 A2 B0 VDD Y GND
M1 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A2 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_11 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M6 N_7 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi31d0
* SPICE INPUT		Wed Jul 10 13:28:18 2019	aoi31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d1
.subckt aoi31d1 B0 A2 A1 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_11 A1 N_10 GND mn5  l=0.5u w=0.58u m=1
M3 N_11 A2 Y GND mn5  l=0.5u w=0.58u m=1
M4 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_9 A2 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y B0 N_9 VDD mp5  l=0.42u w=0.76u m=1
.ends aoi31d1
* SPICE INPUT		Wed Jul 10 13:28:25 2019	aoi31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d2
.subckt aoi31d2 B0 A2 A1 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_11 A1 N_10 GND mn5  l=0.5u w=0.72u m=1
M3 N_11 A2 Y GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_9 A2 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y B0 N_9 VDD mp5  l=0.42u w=0.96u m=1
.ends aoi31d2
* SPICE INPUT		Wed Jul 10 13:28:32 2019	aoi32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d0
.subckt aoi32d0 GND Y VDD A1 A0 A2 B1 B0
M1 N_5 B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B1 N_5 GND mn5  l=0.5u w=0.5u m=1
M3 Y A2 N_7 GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A1 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_6 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_12 B0 Y VDD mp5  l=0.42u w=0.52u m=1
M7 N_12 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_12 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi32d0
* SPICE INPUT		Wed Jul 10 13:28:40 2019	aoi32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d1
.subckt aoi32d1 GND Y VDD B0 B1 A2 A1 A0
M1 N_6 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_7 A1 N_6 GND mn5  l=0.5u w=0.58u m=1
M3 Y A2 N_7 GND mn5  l=0.5u w=0.58u m=1
M4 Y B1 N_5 GND mn5  l=0.5u w=0.58u m=1
M5 N_5 B0 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_9 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_9 A2 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_9 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M10 N_9 B0 Y VDD mp5  l=0.42u w=0.76u m=1
.ends aoi32d1
* SPICE INPUT		Wed Jul 10 13:28:47 2019	aoi32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d2
.subckt aoi32d2 GND Y VDD A0 A1 A2 B1 B0
M1 N_5 B0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_6 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B1 N_5 GND mn5  l=0.5u w=0.72u m=1
M4 Y A2 N_7 GND mn5  l=0.5u w=0.72u m=1
M5 N_7 A1 N_6 GND mn5  l=0.5u w=0.72u m=1
M6 N_12 B0 Y VDD mp5  l=0.42u w=0.96u m=1
M7 N_12 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_12 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M9 N_12 A2 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_12 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi32d2
* SPICE INPUT		Wed Jul 10 13:28:54 2019	aoi33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d0
.subckt aoi33d0 GND Y VDD B0 B1 B2 A2 A1 A0
M1 N_6 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A1 N_6 GND mn5  l=0.5u w=0.5u m=1
M3 Y A2 N_7 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 B2 Y GND mn5  l=0.5u w=0.5u m=1
M5 N_8 B1 N_5 GND mn5  l=0.5u w=0.5u m=1
M6 N_5 B0 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y B2 N_10 VDD mp5  l=0.42u w=0.52u m=1
M11 Y B1 N_10 VDD mp5  l=0.42u w=0.52u m=1
M12 Y B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends aoi33d0
* SPICE INPUT		Wed Jul 10 13:29:01 2019	aoi33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d1
.subckt aoi33d1 GND Y VDD B0 B1 B2 A2 A1 A0
M1 N_6 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_7 A1 N_6 GND mn5  l=0.5u w=0.58u m=1
M3 Y A2 N_7 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 B2 Y GND mn5  l=0.5u w=0.58u m=1
M5 N_8 B1 N_5 GND mn5  l=0.5u w=0.58u m=1
M6 N_5 B0 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_11 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_11 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_11 A2 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y B2 N_11 VDD mp5  l=0.42u w=0.76u m=1
M11 Y B1 N_11 VDD mp5  l=0.42u w=0.76u m=1
M12 Y B0 N_11 VDD mp5  l=0.42u w=0.76u m=1
.ends aoi33d1
* SPICE INPUT		Wed Jul 10 13:29:08 2019	aoi33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d2
.subckt aoi33d2 GND Y VDD A0 A1 B1 A2 B2 B0
M1 N_8 B1 N_5 GND mn5  l=0.5u w=0.72u m=1
M2 N_6 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_8 B2 Y GND mn5  l=0.5u w=0.72u m=1
M4 Y A2 N_7 GND mn5  l=0.5u w=0.72u m=1
M5 N_5 B0 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_7 A1 N_6 GND mn5  l=0.5u w=0.72u m=1
M7 Y B1 N_14 VDD mp5  l=0.42u w=0.96u m=1
M8 N_14 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y B2 N_14 VDD mp5  l=0.42u w=0.96u m=1
M10 N_14 A2 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 Y B0 N_14 VDD mp5  l=0.42u w=0.96u m=1
M12 N_14 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi33d2
* SPICE INPUT		Wed Jul 10 13:29:15 2019	aoim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d0
.subckt aoim21d0 A1N A0N B0 GND VDD Y
M1 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 A0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1N GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 N_13 VDD mp5  l=0.42u w=0.52u m=1
M6 N_13 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_14 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A1N N_14 VDD mp5  l=0.42u w=0.52u m=1
.ends aoim21d0
* SPICE INPUT		Wed Jul 10 13:29:22 2019	aoim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d1
.subckt aoim21d1 B0 A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_14 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_13 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y B0 N_13 VDD mp5  l=0.42u w=0.76u m=1
.ends aoim21d1
* SPICE INPUT		Wed Jul 10 13:29:30 2019	aoim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d2
.subckt aoim21d2 B0 A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_14 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_13 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y B0 N_13 VDD mp5  l=0.42u w=0.96u m=1
.ends aoim21d2
* SPICE INPUT		Wed Jul 10 13:29:37 2019	aoim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d0
.subckt aoim22d0 B1 B0 A1N A0N GND VDD Y
M1 N_2 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_16 B0 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_16 B1 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 A1N N_11 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_10 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends aoim22d0
* SPICE INPUT		Wed Jul 10 13:29:45 2019	aoim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d1
.subckt aoim22d1 B0 B1 A1N A0N VDD Y GND
M1 N_2 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B1 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_11 B0 Y GND mn5  l=0.5u w=0.58u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_18 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 A1N N_18 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B1 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_10 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y N_2 N_10 VDD mp5  l=0.42u w=0.76u m=1
.ends aoim22d1
* SPICE INPUT		Wed Jul 10 13:29:52 2019	aoim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d2
.subckt aoim22d2 B0 B1 A1N A0N GND Y VDD
M1 N_2 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B1 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_11 B0 Y GND mn5  l=0.5u w=0.72u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_18 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 A1N N_18 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B1 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_10 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y N_2 N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends aoim22d2
* SPICE INPUT		Wed Jul 10 13:29:59 2019	aoim31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim31d0
.subckt aoim31d0 B0 A2N A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_12 A1N N_11 VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 A2N N_12 VDD mp5  l=0.42u w=0.52u m=1
M9 N_10 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends aoim31d0
* SPICE INPUT		Wed Jul 10 13:30:07 2019	aoim31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim31d1
.subckt aoim31d1 B0 A2N A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_15 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_16 A1N N_15 VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 A2N N_16 VDD mp5  l=0.42u w=0.52u m=1
M9 N_14 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y B0 N_14 VDD mp5  l=0.42u w=0.76u m=1
.ends aoim31d1
* SPICE INPUT		Wed Jul 10 13:30:14 2019	aoim31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim31d2
.subckt aoim31d2 B0 A2N A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_15 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_16 A1N N_15 VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 A2N N_16 VDD mp5  l=0.42u w=0.52u m=1
M9 N_14 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y B0 N_14 VDD mp5  l=0.42u w=0.96u m=1
.ends aoim31d2
* SPICE INPUT		Wed Jul 10 13:30:21 2019	aor211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d0
.subckt aor211d0 C0 B0 A0 A1 GND Y VDD
M1 N_11 A1 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 C0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 C0 N_18 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor211d0
* SPICE INPUT		Wed Jul 10 13:30:29 2019	aor211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d1
.subckt aor211d1 C0 B0 A0 A1 VDD Y GND
M1 N_11 A1 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 C0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 C0 N_18 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aor211d1
* SPICE INPUT		Wed Jul 10 13:30:36 2019	aor211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d2
.subckt aor211d2 A1 A0 B0 C0 GND Y VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_6 C0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 A1 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_6 C0 N_18 VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 B0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor211d2
* SPICE INPUT		Wed Jul 10 13:30:43 2019	aor21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d0
.subckt aor21d0 B0 A1 A0 VDD Y GND
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor21d0
* SPICE INPUT		Wed Jul 10 13:30:50 2019	aor21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d1
.subckt aor21d1 B0 A1 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_3 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_3 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
.ends aor21d1
* SPICE INPUT		Wed Jul 10 13:30:58 2019	aor21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d2
.subckt aor21d2 B0 A1 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_3 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_3 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
.ends aor21d2
* SPICE INPUT		Wed Jul 10 13:31:05 2019	aor221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d0
.subckt aor221d0 GND Y VDD C0 A0 A1 B1 B0
M1 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B1 N_4 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_14 A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A0 N_14 VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_14 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_14 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor221d0
* SPICE INPUT		Wed Jul 10 13:31:12 2019	aor221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d1
.subckt aor221d1 GND Y VDD C0 A0 A1 B1 B0
M1 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_8 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B1 N_4 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_14 A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A0 N_14 VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M11 N_14 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_14 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor221d1
* SPICE INPUT		Wed Jul 10 13:31:19 2019	aor221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d2
.subckt aor221d2 GND Y VDD C0 A0 A1 B1 B0
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_8 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B1 N_4 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_14 A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A0 N_14 VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 N_14 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_14 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor221d2
* SPICE INPUT		Wed Jul 10 13:31:26 2019	aor22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d0
.subckt aor22d0 B0 B1 A1 A0 Y GND VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_12 B1 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B1 N_9 VDD mp5  l=0.42u w=0.52u m=1
M10 N_9 B0 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends aor22d0
* SPICE INPUT		Wed Jul 10 13:31:34 2019	aor22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d1
.subckt aor22d1 A0 A1 B1 B0 GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 B1 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_8 B0 N_6 VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B1 N_8 VDD mp5  l=0.42u w=0.52u m=1
M9 N_8 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_8 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor22d1
* SPICE INPUT		Wed Jul 10 13:31:41 2019	aor22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d2
.subckt aor22d2 A0 A1 B1 B0 Y VDD GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 B1 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_7 B0 N_6 VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B1 N_7 VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor22d2
* SPICE INPUT		Wed Jul 10 13:31:48 2019	aor311d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor311d0
.subckt aor311d0 GND Y VDD A2 A0 A1 B0 C0
M1 N_7 A1 N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A0 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_15 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor311d0
* SPICE INPUT		Wed Jul 10 13:31:55 2019	aor311d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor311d1
.subckt aor311d1 GND Y VDD A2 A0 A1 B0 C0
M1 N_7 A1 N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A0 N_7 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_15 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aor311d1
* SPICE INPUT		Wed Jul 10 13:32:02 2019	aor311d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor311d2
.subckt aor311d2 GND Y VDD A2 A0 A1 B0 C0
M1 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A1 N_4 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A0 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_15 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aor311d2
* SPICE INPUT		Wed Jul 10 13:32:10 2019	aor31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d0
.subckt aor31d0 B0 A2 A1 A0 Y VDD GND
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A2 N_12 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_9 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor31d0
* SPICE INPUT		Wed Jul 10 13:32:17 2019	aor31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d1
.subckt aor31d1 B0 A2 A1 A0 GND Y VDD
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A2 N_12 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aor31d1
* SPICE INPUT		Wed Jul 10 13:32:24 2019	aor31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d2
.subckt aor31d2 B0 A2 A1 A0 GND Y VDD
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A2 N_12 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aor31d2
* SPICE INPUT		Wed Jul 10 13:32:31 2019	buffd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd0
.subckt buffd0 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends buffd0
* SPICE INPUT		Wed Jul 10 13:32:39 2019	buffd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd1
.subckt buffd1 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends buffd1
* SPICE INPUT		Wed Jul 10 13:32:46 2019	buffd10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd10
.subckt buffd10 GND Y VDD A
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M7 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 N_4 A VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_4 A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buffd10
* SPICE INPUT		Wed Jul 10 13:32:53 2019	buffd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd2
.subckt buffd2 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.58u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends buffd2
* SPICE INPUT		Wed Jul 10 13:33:00 2019	buffd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd3
.subckt buffd3 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.74u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.34u m=1
M3 N_4 A GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.72u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.72u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends buffd3
* SPICE INPUT		Wed Jul 10 13:33:08 2019	buffd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd4
.subckt buffd4 GND Y VDD A
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buffd4
* SPICE INPUT		Wed Jul 10 13:33:15 2019	buffd5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd5
.subckt buffd5 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.613u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.613u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.574u m=1
M4 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y N_4 VDD VDD mp5  l=0.42u w=0.48u m=1
M8 VDD A N_4 VDD mp5  l=0.42u w=0.96u m=1
.ends buffd5
* SPICE INPUT		Wed Jul 10 13:33:22 2019	buffd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd6
.subckt buffd6 GND Y VDD A
M1 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buffd6
* SPICE INPUT		Wed Jul 10 13:33:30 2019	buffd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd8
.subckt buffd8 GND Y VDD A
M1 N_4 A GND GND mn5  l=0.5u w=0.54u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.54u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_4 A VDD VDD mp5  l=0.42u w=0.72u m=1
M8 N_4 A VDD VDD mp5  l=0.42u w=0.72u m=1
M9 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buffd8
* SPICE INPUT		Wed Jul 10 13:33:37 2019	buftd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd0
.subckt buftd0 OE A GND Y VDD
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_3 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 OE GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_3 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 OE N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftd0
* SPICE INPUT		Wed Jul 10 13:33:44 2019	buftd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd1
.subckt buftd1 OE A GND Y VDD
M1 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_3 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 OE GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_3 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 OE N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftd1
* SPICE INPUT		Wed Jul 10 13:33:51 2019	buftd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd2
.subckt buftd2 A OE Y GND VDD
M1 N_4 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_6 OE N_2 VDD mp5  l=0.42u w=0.52u m=1
.ends buftd2
* SPICE INPUT		Wed Jul 10 13:33:59 2019	buftld0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld0
.subckt buftld0 A OE GND VDD Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 N_2 N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld0
* SPICE INPUT		Wed Jul 10 13:34:06 2019	buftld1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld1
.subckt buftld1 A OE GND VDD Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 N_2 N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld1
* SPICE INPUT		Wed Jul 10 13:34:13 2019	buftld2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld2
.subckt buftld2 A OE VDD Y GND
M1 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_5 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_6 N_5 N_2 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld2



* SPICE INPUT		Wed Jul 10 13:37:55 2019	dl01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d0
.subckt dl01d0 A GND VDD Y
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dl01d0
* SPICE INPUT		Wed Jul 10 13:38:03 2019	dl01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d1
.subckt dl01d1 A GND VDD Y
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dl01d1
* SPICE INPUT		Wed Jul 10 13:38:10 2019	dl01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d2
.subckt dl01d2 A GND VDD Y
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dl01d2
* SPICE INPUT		Wed Jul 10 13:38:17 2019	dl02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d0
.subckt dl02d0 A Y VDD GND
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=1u w=0.5u m=1
M3 N_4 N_3 GND GND mn5  l=1u w=0.5u m=1
M4 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_5 N_4 VDD VDD mp5  l=0.84u w=0.52u m=1
M7 N_4 N_3 VDD VDD mp5  l=0.84u w=0.52u m=1
M8 N_3 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dl02d0
* SPICE INPUT		Wed Jul 10 13:38:24 2019	dl02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d1
.subckt dl02d1 A VDD Y GND
M1 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_4 GND GND mn5  l=1u w=0.5u m=1
M3 N_4 N_3 GND GND mn5  l=1u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_3 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.84u w=0.52u m=1
M7 N_4 N_3 VDD VDD mp5  l=0.84u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dl02d1
* SPICE INPUT		Wed Jul 10 13:38:32 2019	dl02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d2
.subckt dl02d2 A VDD Y GND
M1 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_4 GND GND mn5  l=1u w=0.5u m=1
M3 N_4 N_3 GND GND mn5  l=1u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_3 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.84u w=0.52u m=1
M7 N_4 N_3 VDD VDD mp5  l=0.84u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dl02d2


* SPICE INPUT		Wed Jul 10 13:38:39 2019	inv0d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d0
.subckt inv0d0 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.5u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends inv0d0
* SPICE INPUT		Wed Jul 10 13:38:46 2019	inv0d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d1
.subckt inv0d1 VDD Y GND A
M1 Y A GND GND mn5  l=0.5u w=0.58u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends inv0d1
* SPICE INPUT		Wed Jul 10 13:38:53 2019	inv0d10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d10
.subckt inv0d10 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A GND GND mn5  l=0.5u w=0.72u m=1
M5 Y A GND GND mn5  l=0.5u w=0.72u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d10
* SPICE INPUT		Wed Jul 10 13:39:00 2019	inv0d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d2
.subckt inv0d2 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d2
* SPICE INPUT		Wed Jul 10 13:39:08 2019	inv0d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d3
.subckt inv0d3 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.54u m=1
M2 Y A GND GND mn5  l=0.5u w=0.54u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.72u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.72u m=1
.ends inv0d3
* SPICE INPUT		Wed Jul 10 13:39:15 2019	inv0d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d4
.subckt inv0d4 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d4
* SPICE INPUT		Wed Jul 10 13:39:22 2019	inv0d5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d5
.subckt inv0d5 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.6u m=1
M2 Y A GND GND mn5  l=0.5u w=0.6u m=1
M3 Y A GND GND mn5  l=0.5u w=0.6u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.8u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.8u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.8u m=1
.ends inv0d5
* SPICE INPUT		Wed Jul 10 13:39:29 2019	inv0d6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d6
.subckt inv0d6 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d6
* SPICE INPUT		Wed Jul 10 13:39:36 2019	inv0d8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d8
.subckt inv0d8 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A GND GND mn5  l=0.5u w=0.72u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d8
* SPICE INPUT		Wed Jul 10 13:39:43 2019	invtd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtd0
.subckt invtd0 GND Y VDD OE A
M1 N_4 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_6 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y OE N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends invtd0
* SPICE INPUT		Wed Jul 10 13:39:51 2019	invtd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtd1
.subckt invtd1 A OE VDD GND Y
M1 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A GND GND mn5  l=0.5u w=0.58u m=1
M3 Y N_2 N_9 GND mn5  l=0.5u w=0.58u m=1
M4 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_14 A VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y OE N_14 VDD mp5  l=0.42u w=0.76u m=1
.ends invtd1
* SPICE INPUT		Wed Jul 10 13:39:58 2019	invtd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtd2
.subckt invtd2 A OE VDD GND Y
M1 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y N_2 N_9 GND mn5  l=0.5u w=0.72u m=1
M4 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_14 A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y OE N_14 VDD mp5  l=0.42u w=0.96u m=1
.ends invtd2
* SPICE INPUT		Wed Jul 10 13:40:05 2019	invtld0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld0
.subckt invtld0 GND Y VDD OE A
M1 N_4 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 Y OE N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_6 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 Y N_4 N_13 VDD mp5  l=0.42u w=0.52u m=1
M6 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends invtld0
* SPICE INPUT		Wed Jul 10 13:40:12 2019	invtld1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld1
.subckt invtld1 OE A GND VDD Y
M1 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A GND GND mn5  l=0.5u w=0.58u m=1
M3 Y OE N_9 GND mn5  l=0.5u w=0.58u m=1
M4 N_5 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_14 A VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y N_5 N_14 VDD mp5  l=0.42u w=0.76u m=1
.ends invtld1
* SPICE INPUT		Wed Jul 10 13:40:19 2019	invtld2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld2
.subckt invtld2 OE A GND VDD Y
M1 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y OE N_9 GND mn5  l=0.5u w=0.72u m=1
M4 N_5 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_14 A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y N_5 N_14 VDD mp5  l=0.42u w=0.96u m=1
.ends invtld2

* SPICE INPUT		Wed Jul 10 13:44:02 2019	mi02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d0
.subckt mi02d0 VDD Y GND S0 B A
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 N_3 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_5 S0 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y S0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mi02d0
* SPICE INPUT		Wed Jul 10 13:44:09 2019	mi02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d1
.subckt mi02d1 GND Y VDD A B S0
M1 N_5 B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 N_4 GND mn5  l=0.5u w=0.58u m=1
M3 Y S0 N_5 GND mn5  l=0.5u w=0.58u m=1
M4 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_3 N_5 VDD mp5  l=0.42u w=0.76u m=1
M7 N_5 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y S0 N_4 VDD mp5  l=0.42u w=0.76u m=1
M9 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mi02d1
* SPICE INPUT		Wed Jul 10 13:44:16 2019	mi02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d2
.subckt mi02d2 GND Y VDD S0 B A
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 N_4 GND mn5  l=0.5u w=0.72u m=1
M3 Y S0 N_5 GND mn5  l=0.5u w=0.72u m=1
M4 N_5 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y S0 N_4 VDD mp5  l=0.42u w=0.96u m=1
M8 Y N_3 N_5 VDD mp5  l=0.42u w=0.96u m=1
M9 N_5 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mi02d2
* SPICE INPUT		Wed Jul 10 13:44:23 2019	mi04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi04d0
.subckt mi04d0 VDD Y GND D C S0 B A S1
M1 N_11 N_13 N_15 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_7 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_10 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_7 S0 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_15 S1 N_12 GND mn5  l=0.5u w=0.5u m=1
M10 N_13 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M12 N_6 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 N_7 N_5 GND mn5  l=0.5u w=0.5u m=1
M14 N_5 C GND GND mn5  l=0.5u w=0.5u m=1
M15 Y N_15 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_15 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M17 N_12 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_11 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 S0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 S0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M23 N_10 N_7 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 S1 N_11 VDD mp5  l=0.42u w=0.52u m=1
M25 N_13 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 D VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 N_7 N_4 VDD mp5  l=0.42u w=0.52u m=1
M29 N_5 C VDD VDD mp5  l=0.42u w=0.52u m=1
M30 Y N_15 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mi04d0
* SPICE INPUT		Wed Jul 10 13:44:30 2019	mi04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi04d1
.subckt mi04d1 VDD Y GND C D S0 B A S1
M1 N_11 N_15 N_14 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_7 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_10 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_7 S0 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_14 S1 N_12 GND mn5  l=0.5u w=0.5u m=1
M10 N_15 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M12 N_6 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 N_7 N_5 GND mn5  l=0.5u w=0.5u m=1
M14 N_5 C GND GND mn5  l=0.5u w=0.5u m=1
M15 Y N_14 GND GND mn5  l=0.5u w=0.58u m=1
M16 N_14 N_15 N_12 VDD mp5  l=0.42u w=0.52u m=1
M17 N_12 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_11 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 S0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 S0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M23 N_10 N_7 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 S1 N_11 VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 D VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 N_7 N_4 VDD mp5  l=0.42u w=0.52u m=1
M29 N_5 C VDD VDD mp5  l=0.42u w=0.52u m=1
M30 Y N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends mi04d1
* SPICE INPUT		Wed Jul 10 13:44:37 2019	mi04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi04d2
.subckt mi04d2 GND Y VDD C D S0 B A S1
M1 N_11 N_13 N_14 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_10 N_7 N_9 GND mn5  l=0.5u w=0.5u m=1
M6 N_6 S0 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_9 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_7 S0 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_14 S1 N_12 GND mn5  l=0.5u w=0.5u m=1
M10 N_13 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_6 N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M14 N_4 C GND GND mn5  l=0.5u w=0.5u m=1
M15 Y N_14 GND GND mn5  l=0.5u w=0.72u m=1
M16 N_14 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M17 N_12 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_10 A VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_4 S0 N_6 VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 S0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M23 N_9 N_7 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 S1 N_11 VDD mp5  l=0.42u w=0.52u m=1
M25 N_13 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 D VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_5 N_7 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_4 C VDD VDD mp5  l=0.42u w=0.52u m=1
M30 Y N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends mi04d2
* SPICE INPUT		Wed Jul 10 13:44:45 2019	mx02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d0
.subckt mx02d0 VDD Y GND S0 B A
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 S0 N_5 VDD mp5  l=0.42u w=0.52u m=1
M11 N_7 N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mx02d0
* SPICE INPUT		Wed Jul 10 13:44:52 2019	mx02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d1
.subckt mx02d1 GND Y VDD S0 B A
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 S0 N_5 VDD mp5  l=0.42u w=0.52u m=1
M11 N_7 N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mx02d1
* SPICE INPUT		Wed Jul 10 13:44:59 2019	mx02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d2
.subckt mx02d2 GND Y VDD S0 B A
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 S0 N_5 VDD mp5  l=0.42u w=0.52u m=1
M11 N_7 N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mx02d2
* SPICE INPUT		Wed Jul 10 13:45:06 2019	mx04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d0
.subckt mx04d0 GND Y VDD S1 A B S0 D C
M1 N_3 N_14 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 S1 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_8 D GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 B GND GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_10 N_3 GND mn5  l=0.5u w=0.5u m=1
M9 N_13 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_14 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_4 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_10 S0 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_3 S0 N_11 GND mn5  l=0.5u w=0.5u m=1
M14 N_4 N_14 N_2 VDD mp5  l=0.42u w=0.5u m=1
M15 N_2 S1 N_3 VDD mp5  l=0.42u w=0.5u m=1
M16 N_7 C VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_8 N_10 N_4 VDD mp5  l=0.42u w=0.5u m=1
M18 N_8 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_11 B VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_3 N_10 N_11 VDD mp5  l=0.42u w=0.5u m=1
M22 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_4 S0 N_7 VDD mp5  l=0.42u w=0.5u m=1
M25 N_10 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_3 S0 N_13 VDD mp5  l=0.42u w=0.5u m=1
.ends mx04d0
* SPICE INPUT		Wed Jul 10 13:45:13 2019	mx04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d1
.subckt mx04d1 GND Y VDD S1 A B S0 D C
M1 N_3 N_14 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 S1 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_8 D GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 B GND GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_10 N_3 GND mn5  l=0.5u w=0.5u m=1
M9 N_13 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_14 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_4 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_10 S0 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_3 S0 N_11 GND mn5  l=0.5u w=0.5u m=1
M14 N_4 N_14 N_2 VDD mp5  l=0.42u w=0.5u m=1
M15 N_2 S1 N_3 VDD mp5  l=0.42u w=0.5u m=1
M16 N_7 C VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_8 N_10 N_4 VDD mp5  l=0.42u w=0.5u m=1
M18 N_8 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_11 B VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_3 N_10 N_11 VDD mp5  l=0.42u w=0.5u m=1
M22 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_4 S0 N_7 VDD mp5  l=0.42u w=0.5u m=1
M25 N_10 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_3 S0 N_13 VDD mp5  l=0.42u w=0.5u m=1
.ends mx04d1
* SPICE INPUT		Wed Jul 10 13:45:20 2019	mx04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d2
.subckt mx04d2 GND Y VDD S1 A B S0 D C
M1 N_3 N_14 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 S1 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_8 D GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 B GND GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_10 N_3 GND mn5  l=0.5u w=0.5u m=1
M9 N_13 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_14 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_4 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_10 S0 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_3 S0 N_11 GND mn5  l=0.5u w=0.5u m=1
M14 N_4 N_14 N_2 VDD mp5  l=0.42u w=0.5u m=1
M15 N_2 S1 N_3 VDD mp5  l=0.42u w=0.5u m=1
M16 N_7 C VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_8 N_10 N_4 VDD mp5  l=0.42u w=0.5u m=1
M18 N_8 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_11 B VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_3 N_10 N_11 VDD mp5  l=0.42u w=0.5u m=1
M22 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_4 S0 N_7 VDD mp5  l=0.42u w=0.5u m=1
M25 N_10 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_3 S0 N_13 VDD mp5  l=0.42u w=0.5u m=1
.ends mx04d2
* SPICE INPUT		Wed Jul 10 13:45:27 2019	nd02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d0
.subckt nd02d0 VDD Y GND B A
M1 Y A N_8 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd02d0
* SPICE INPUT		Wed Jul 10 13:45:35 2019	nd02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d1
.subckt nd02d1 VDD Y GND B A
M1 Y A N_8 GND mn5  l=0.5u w=0.58u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.58u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.76u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd02d1
* SPICE INPUT		Wed Jul 10 13:45:42 2019	nd02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d2
.subckt nd02d2 GND Y VDD B A
M1 Y A N_5 GND mn5  l=0.5u w=0.72u m=1
M2 N_5 B GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd02d2
* SPICE INPUT		Wed Jul 10 13:45:49 2019	nd03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d0
.subckt nd03d0 C B A Y VDD GND
M1 Y A N_8 GND mn5  l=0.5u w=0.5u m=1
M2 N_9 B N_8 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 C GND GND mn5  l=0.5u w=0.5u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd03d0
* SPICE INPUT		Wed Jul 10 13:45:56 2019	nd03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d1
.subckt nd03d1 A B C VDD GND Y
M1 N_9 C GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 B N_8 GND mn5  l=0.5u w=0.58u m=1
M3 Y A N_8 GND mn5  l=0.5u w=0.58u m=1
M4 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M5 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd03d1
* SPICE INPUT		Wed Jul 10 13:46:03 2019	nd03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d2
.subckt nd03d2 C B A Y VDD GND
M1 Y A N_8 GND mn5  l=0.5u w=0.72u m=1
M2 N_9 B N_8 GND mn5  l=0.5u w=0.72u m=1
M3 N_9 C GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M5 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd03d2
* SPICE INPUT		Wed Jul 10 13:46:10 2019	nd04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d0
.subckt nd04d0 C B D A GND VDD Y
M1 Y A N_9 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B N_9 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 C N_10 GND mn5  l=0.5u w=0.5u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y D VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd04d0
* SPICE INPUT		Wed Jul 10 13:46:17 2019	nd04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d1
.subckt nd04d1 GND Y VDD A B C D
M1 N_6 D GND GND mn5  l=0.5u w=0.58u m=1
M2 N_7 C N_6 GND mn5  l=0.5u w=0.58u m=1
M3 N_7 B N_5 GND mn5  l=0.5u w=0.58u m=1
M4 Y A N_5 GND mn5  l=0.5u w=0.58u m=1
M5 Y D VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M7 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd04d1
* SPICE INPUT		Wed Jul 10 13:46:24 2019	nd04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d2
.subckt nd04d2 D C B A Y VDD GND
M1 Y A N_9 GND mn5  l=0.5u w=0.72u m=1
M2 N_11 B N_9 GND mn5  l=0.5u w=0.72u m=1
M3 N_11 C N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_10 D GND GND mn5  l=0.5u w=0.72u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y D VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd04d2
* SPICE INPUT		Wed Jul 10 13:46:32 2019	nd12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d0
.subckt nd12d0 B AN Y VDD GND
M1 Y N_4 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd12d0
* SPICE INPUT		Wed Jul 10 13:46:39 2019	nd12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d1
.subckt nd12d1 B AN Y VDD GND
M1 Y N_4 N_12 GND mn5  l=0.5u w=0.58u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 B GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd12d1
* SPICE INPUT		Wed Jul 10 13:46:46 2019	nd12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d2
.subckt nd12d2 B AN Y VDD GND
M1 Y N_4 N_8 GND mn5  l=0.5u w=0.72u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd12d2
* SPICE INPUT		Wed Jul 10 13:46:53 2019	nd13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d0
.subckt nd13d0 GND Y VDD B C AN
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 C GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd13d0
* SPICE INPUT		Wed Jul 10 13:47:00 2019	nd13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d1
.subckt nd13d1 C AN B Y VDD GND
M1 Y N_5 N_9 GND mn5  l=0.5u w=0.58u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.58u m=1
M3 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.58u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd13d1
* SPICE INPUT		Wed Jul 10 13:47:07 2019	nd13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d2
.subckt nd13d2 C AN B Y VDD GND
M1 Y N_5 N_9 GND mn5  l=0.5u w=0.72u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.72u m=1
M3 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd13d2
* SPICE INPUT		Wed Jul 10 13:47:15 2019	nd14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d0
.subckt nd14d0 GND Y VDD B C D AN
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 C N_7 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 B N_6 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y D VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd14d0
* SPICE INPUT		Wed Jul 10 13:47:22 2019	nd14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d1
.subckt nd14d1 GND Y VDD B C D AN
M1 N_8 B N_6 GND mn5  l=0.5u w=0.58u m=1
M2 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M3 N_7 D GND GND mn5  l=0.5u w=0.58u m=1
M4 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 N_6 GND mn5  l=0.5u w=0.58u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
M7 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y D VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd14d1
* SPICE INPUT		Wed Jul 10 13:47:29 2019	nd14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d2
.subckt nd14d2 GND Y VDD B C D AN
M1 N_8 B N_6 GND mn5  l=0.5u w=0.72u m=1
M2 N_8 C N_7 GND mn5  l=0.5u w=0.72u m=1
M3 N_7 D GND GND mn5  l=0.5u w=0.72u m=1
M4 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 N_6 GND mn5  l=0.5u w=0.72u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y D VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd14d2
* SPICE INPUT		Wed Jul 10 13:47:36 2019	nd23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd23d0
.subckt nd23d0 AN C BN GND Y VDD
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd23d0
* SPICE INPUT		Wed Jul 10 13:47:44 2019	nd23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd23d1
.subckt nd23d1 AN C BN GND Y VDD
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 N_11 GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_4 N_10 GND mn5  l=0.5u w=0.58u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.58u m=1
M5 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M10 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd23d1
* SPICE INPUT		Wed Jul 10 13:47:51 2019	nd23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd23d2
.subckt nd23d2 AN C BN GND Y VDD
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 N_11 GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_4 N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.72u m=1
M5 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd23d2
* SPICE INPUT		Wed Jul 10 13:47:58 2019	nd24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d0
.subckt nd24d0 GND Y VDD D AN C BN
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 C N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
M11 Y D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd24d0
* SPICE INPUT		Wed Jul 10 13:48:05 2019	nd24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d1
.subckt nd24d1 GND Y VDD D AN C BN
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 N_9 GND mn5  l=0.5u w=0.58u m=1
M3 N_9 N_3 N_8 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M5 N_7 D GND GND mn5  l=0.5u w=0.58u m=1
M6 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M11 Y D VDD VDD mp5  l=0.42u w=0.76u m=1
M12 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd24d1
* SPICE INPUT		Wed Jul 10 13:48:12 2019	nd24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d2
.subckt nd24d2 GND Y VDD D AN C BN
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 N_9 GND mn5  l=0.5u w=0.72u m=1
M3 N_9 N_3 N_8 GND mn5  l=0.5u w=0.72u m=1
M4 N_8 C N_7 GND mn5  l=0.5u w=0.72u m=1
M5 N_7 D GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M11 Y D VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd24d2
* SPICE INPUT		Wed Jul 10 13:48:19 2019	nr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d0
.subckt nr02d0 GND Y VDD B A
M1 Y A GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A VDD VDD mp5  l=0.42u w=0.52u m=1
M4 Y B N_7 VDD mp5  l=0.42u w=0.52u m=1
.ends nr02d0
* SPICE INPUT		Wed Jul 10 13:48:26 2019	nr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d1
.subckt nr02d1 GND Y VDD B A
M1 Y A GND GND mn5  l=0.5u w=0.58u m=1
M2 Y B GND GND mn5  l=0.5u w=0.58u m=1
M3 N_7 A VDD VDD mp5  l=0.42u w=0.76u m=1
M4 Y B N_7 VDD mp5  l=0.42u w=0.76u m=1
.ends nr02d1
* SPICE INPUT		Wed Jul 10 13:48:34 2019	nr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d2
.subckt nr02d2 GND Y VDD B A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y B GND GND mn5  l=0.5u w=0.72u m=1
M3 N_7 A VDD VDD mp5  l=0.42u w=0.96u m=1
M4 Y B N_7 VDD mp5  l=0.42u w=0.96u m=1
.ends nr02d2
* SPICE INPUT		Wed Jul 10 13:48:41 2019	nr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d0
.subckt nr03d0 A B C Y VDD GND
M1 Y C GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y A GND GND mn5  l=0.5u w=0.5u m=1
M4 Y C N_8 VDD mp5  l=0.42u w=0.52u m=1
M5 N_9 B N_8 VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr03d0
* SPICE INPUT		Wed Jul 10 13:48:48 2019	nr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d1
.subckt nr03d1 A B C GND VDD Y
M1 Y C GND GND mn5  l=0.5u w=0.58u m=1
M2 Y B GND GND mn5  l=0.5u w=0.58u m=1
M3 Y A GND GND mn5  l=0.5u w=0.58u m=1
M4 Y C N_11 VDD mp5  l=0.42u w=0.76u m=1
M5 N_12 B N_11 VDD mp5  l=0.42u w=0.76u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nr03d1
* SPICE INPUT		Wed Jul 10 13:48:55 2019	nr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d2
.subckt nr03d2 A B C GND VDD Y
M1 Y C GND GND mn5  l=0.5u w=0.72u m=1
M2 Y B GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C N_11 VDD mp5  l=0.42u w=0.96u m=1
M5 N_12 B N_11 VDD mp5  l=0.42u w=0.96u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nr03d2
* SPICE INPUT		Wed Jul 10 13:49:02 2019	nr04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d0
.subckt nr04d0 A B C D Y VDD GND
M1 Y D GND GND mn5  l=0.5u w=0.5u m=1
M2 Y C GND GND mn5  l=0.5u w=0.5u m=1
M3 Y B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y D N_9 VDD mp5  l=0.42u w=0.52u m=1
M6 N_11 C N_9 VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 B N_10 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr04d0
* SPICE INPUT		Wed Jul 10 13:49:10 2019	nr04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d1
.subckt nr04d1 A B C D GND VDD Y
M1 Y D GND GND mn5  l=0.5u w=0.58u m=1
M2 Y C GND GND mn5  l=0.5u w=0.58u m=1
M3 Y B GND GND mn5  l=0.5u w=0.58u m=1
M4 Y A GND GND mn5  l=0.5u w=0.58u m=1
M5 Y D N_12 VDD mp5  l=0.42u w=0.76u m=1
M6 N_14 C N_12 VDD mp5  l=0.42u w=0.76u m=1
M7 N_14 B N_13 VDD mp5  l=0.42u w=0.76u m=1
M8 N_13 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nr04d1
* SPICE INPUT		Wed Jul 10 13:49:17 2019	nr04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d2
.subckt nr04d2 A B C D GND VDD Y
M1 Y D GND GND mn5  l=0.5u w=0.72u m=1
M2 Y C GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A GND GND mn5  l=0.5u w=0.72u m=1
M5 Y D N_12 VDD mp5  l=0.42u w=0.96u m=1
M6 N_14 C N_12 VDD mp5  l=0.42u w=0.96u m=1
M7 N_14 B N_13 VDD mp5  l=0.42u w=0.96u m=1
M8 N_13 A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nr04d2
* SPICE INPUT		Wed Jul 10 13:49:24 2019	nr12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d0
.subckt nr12d0 AN B Y VDD GND
M1 Y B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 Y B N_8 VDD mp5  l=0.42u w=0.52u m=1
M5 N_8 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr12d0
* SPICE INPUT		Wed Jul 10 13:49:31 2019	nr12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d1
.subckt nr12d1 B AN GND VDD Y
M1 N_2 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.58u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_2 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M5 Y B N_12 VDD mp5  l=0.42u w=0.76u m=1
M6 N_12 N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nr12d1
* SPICE INPUT		Wed Jul 10 13:49:38 2019	nr12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d2
.subckt nr12d2 B AN GND VDD Y
M1 N_2 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.72u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_2 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M5 Y B N_12 VDD mp5  l=0.42u w=0.96u m=1
M6 N_12 N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nr12d2
* SPICE INPUT		Wed Jul 10 13:49:45 2019	nr13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d0
.subckt nr13d0 AN B C Y VDD GND
M1 Y C GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_3 AN GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C N_9 VDD mp5  l=0.42u w=0.52u m=1
M6 N_10 B N_9 VDD mp5  l=0.42u w=0.52u m=1
M7 N_10 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr13d0
* SPICE INPUT		Wed Jul 10 13:49:53 2019	nr13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d1
.subckt nr13d1 C B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M3 Y B GND GND mn5  l=0.5u w=0.58u m=1
M4 Y C GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_10 N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_10 B N_9 VDD mp5  l=0.42u w=0.76u m=1
M8 Y C N_9 VDD mp5  l=0.42u w=0.76u m=1
.ends nr13d1
* SPICE INPUT		Wed Jul 10 13:50:00 2019	nr13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d2
.subckt nr13d2 C B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_14 B N_13 VDD mp5  l=0.42u w=0.96u m=1
M8 Y C N_13 VDD mp5  l=0.42u w=0.96u m=1
.ends nr13d2
* SPICE INPUT		Wed Jul 10 13:50:07 2019	nr14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d0
.subckt nr14d0 D C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 Y B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y C GND GND mn5  l=0.5u w=0.5u m=1
M5 Y D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_16 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M10 Y D N_14 VDD mp5  l=0.42u w=0.52u m=1
.ends nr14d0
* SPICE INPUT		Wed Jul 10 13:50:14 2019	nr14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d1
.subckt nr14d1 D C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M3 Y B GND GND mn5  l=0.5u w=0.58u m=1
M4 Y C GND GND mn5  l=0.5u w=0.58u m=1
M5 Y D GND GND mn5  l=0.5u w=0.58u m=1
M6 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_12 B N_11 VDD mp5  l=0.42u w=0.76u m=1
M9 N_12 C N_10 VDD mp5  l=0.42u w=0.76u m=1
M10 Y D N_10 VDD mp5  l=0.42u w=0.76u m=1
.ends nr14d1
* SPICE INPUT		Wed Jul 10 13:50:21 2019	nr14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d2
.subckt nr14d2 D C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C GND GND mn5  l=0.5u w=0.72u m=1
M5 Y D GND GND mn5  l=0.5u w=0.72u m=1
M6 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_12 B N_11 VDD mp5  l=0.42u w=0.96u m=1
M9 N_12 C N_10 VDD mp5  l=0.42u w=0.96u m=1
M10 Y D N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends nr14d2
* SPICE INPUT		Wed Jul 10 13:50:29 2019	nr23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr23d0
.subckt nr23d0 C AN BN GND VDD Y
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C GND GND mn5  l=0.5u w=0.5u m=1
M6 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_11 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M10 Y C N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends nr23d0
* SPICE INPUT		Wed Jul 10 13:50:36 2019	nr23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr23d1
.subckt nr23d1 C AN BN GND VDD Y
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y C GND GND mn5  l=0.5u w=0.58u m=1
M6 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_11 N_3 N_10 VDD mp5  l=0.42u w=0.76u m=1
M10 Y C N_10 VDD mp5  l=0.42u w=0.76u m=1
.ends nr23d1
* SPICE INPUT		Wed Jul 10 13:50:43 2019	nr23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr23d2
.subckt nr23d2 C AN BN GND VDD Y
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y C GND GND mn5  l=0.5u w=0.72u m=1
M6 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_11 N_3 N_10 VDD mp5  l=0.42u w=0.96u m=1
M10 Y C N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends nr23d2
* SPICE INPUT		Wed Jul 10 13:50:50 2019	nr24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d0
.subckt nr24d0 D C AN BN Y VDD GND
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y D GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_13 N_4 N_12 VDD mp5  l=0.42u w=0.52u m=1
M11 N_13 C N_11 VDD mp5  l=0.42u w=0.52u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends nr24d0
* SPICE INPUT		Wed Jul 10 13:50:57 2019	nr24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d1
.subckt nr24d1 D C AN BN Y VDD GND
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y C GND GND mn5  l=0.5u w=0.58u m=1
M6 Y D GND GND mn5  l=0.5u w=0.58u m=1
M7 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 N_13 N_4 N_12 VDD mp5  l=0.42u w=0.76u m=1
M11 N_13 C N_11 VDD mp5  l=0.42u w=0.76u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=0.76u m=1
.ends nr24d1
* SPICE INPUT		Wed Jul 10 13:51:04 2019	nr24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d2
.subckt nr24d2 D C AN BN Y VDD GND
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y C GND GND mn5  l=0.5u w=0.72u m=1
M6 Y D GND GND mn5  l=0.5u w=0.72u m=1
M7 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_13 N_4 N_12 VDD mp5  l=0.42u w=0.96u m=1
M11 N_13 C N_11 VDD mp5  l=0.42u w=0.96u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=0.96u m=1
.ends nr24d2
* SPICE INPUT		Wed Jul 10 13:51:12 2019	oai211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d0
.subckt oai211d0 C0 B0 A1 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 B0 N_16 GND mn5  l=0.5u w=0.5u m=1
M4 Y C0 N_16 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y A1 N_10 VDD mp5  l=0.42u w=0.52u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai211d0
* SPICE INPUT		Wed Jul 10 13:51:19 2019	oai211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d1
.subckt oai211d1 C0 B0 A1 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 B0 N_16 GND mn5  l=0.5u w=0.58u m=1
M4 Y C0 N_16 GND mn5  l=0.5u w=0.58u m=1
M5 N_10 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y A1 N_10 VDD mp5  l=0.42u w=0.76u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oai211d1
* SPICE INPUT		Wed Jul 10 13:51:26 2019	oai211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d2
.subckt oai211d2 A0 C0 A1 B0 Y VDD GND
M1 N_9 B0 N_10 GND mn5  l=0.5u w=0.72u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y C0 N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_9 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y A1 N_16 VDD mp5  l=0.42u w=0.96u m=1
M7 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_16 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oai211d2
* SPICE INPUT		Wed Jul 10 13:51:33 2019	oai21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d0
.subckt oai21d0 A0 B0 A1 VDD Y GND
M1 N_5 A1 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B0 N_5 GND mn5  l=0.5u w=0.5u m=1
M3 N_5 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 A1 Y VDD mp5  l=0.42u w=0.52u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_12 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai21d0
* SPICE INPUT		Wed Jul 10 13:51:41 2019	oai21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d1
.subckt oai21d1 A0 A1 B0 Y VDD GND
M1 N_5 B0 Y GND mn5  l=0.5u w=0.58u m=1
M2 N_5 A1 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_5 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M5 N_9 A1 Y VDD mp5  l=0.42u w=0.76u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oai21d1
* SPICE INPUT		Wed Jul 10 13:51:48 2019	oai21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d2
.subckt oai21d2 A0 A1 B0 Y VDD GND
M1 N_5 B0 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_5 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_5 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M5 N_9 A1 Y VDD mp5  l=0.42u w=0.96u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oai21d2
* SPICE INPUT		Wed Jul 10 13:51:55 2019	oai221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d0
.subckt oai221d0 C0 B1 A1 A0 B0 Y VDD GND
M1 N_7 B0 N_8 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 B1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_7 GND mn5  l=0.5u w=0.5u m=1
M6 N_13 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_12 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M10 N_13 B1 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oai221d0
* SPICE INPUT		Wed Jul 10 13:52:02 2019	oai221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d1
.subckt oai221d1 C0 B1 A1 A0 B0 Y VDD GND
M1 N_7 B0 N_8 GND mn5  l=0.5u w=0.58u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_8 B1 N_7 GND mn5  l=0.5u w=0.58u m=1
M5 Y C0 N_7 GND mn5  l=0.5u w=0.58u m=1
M6 N_13 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_12 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y A1 N_12 VDD mp5  l=0.42u w=0.76u m=1
M10 N_13 B1 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai221d1
* SPICE INPUT		Wed Jul 10 13:52:10 2019	oai221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d2
.subckt oai221d2 C0 B1 B0 A1 A0 Y VDD GND
M1 N_7 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_7 B0 N_8 GND mn5  l=0.5u w=0.72u m=1
M4 N_7 B1 N_8 GND mn5  l=0.5u w=0.72u m=1
M5 Y C0 N_8 GND mn5  l=0.5u w=0.72u m=1
M6 N_12 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y A1 N_12 VDD mp5  l=0.42u w=0.96u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_13 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_13 B1 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai221d2
* SPICE INPUT		Wed Jul 10 13:52:17 2019	oai222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d0
.subckt oai222d0 B0 A0 A1 B1 C0 C1 Y VDD GND
M1 N_11 C1 Y GND mn5  l=0.5u w=0.5u m=1
M2 N_11 C0 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B1 N_8 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_8 B0 N_11 GND mn5  l=0.5u w=0.5u m=1
M7 N_20 C1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C0 N_20 VDD mp5  l=0.42u w=0.52u m=1
M9 Y B1 N_9 VDD mp5  l=0.42u w=0.52u m=1
M10 Y A1 N_21 VDD mp5  l=0.42u w=0.52u m=1
M11 N_21 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_9 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai222d0
* SPICE INPUT		Wed Jul 10 13:52:24 2019	oai222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d1
.subckt oai222d1 C1 C0 B1 A1 A0 B0 GND VDD Y
M1 N_13 B0 N_10 GND mn5  l=0.5u w=0.58u m=1
M2 N_13 A0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_13 A1 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_10 B1 N_13 GND mn5  l=0.5u w=0.58u m=1
M5 N_10 C0 Y GND mn5  l=0.5u w=0.58u m=1
M6 Y C1 N_10 GND mn5  l=0.5u w=0.58u m=1
M7 N_12 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_21 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y A1 N_21 VDD mp5  l=0.42u w=0.76u m=1
M10 Y B1 N_12 VDD mp5  l=0.42u w=0.76u m=1
M11 Y C0 N_20 VDD mp5  l=0.42u w=0.76u m=1
M12 N_20 C1 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oai222d1
* SPICE INPUT		Wed Jul 10 13:52:31 2019	oai222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d2
.subckt oai222d2 GND Y VDD B0 A0 C1 B1 C0 A1
M1 N_4 C0 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_6 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_6 B0 N_4 GND mn5  l=0.5u w=0.72u m=1
M4 N_6 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 B1 N_6 GND mn5  l=0.5u w=0.72u m=1
M6 N_4 C1 Y GND mn5  l=0.5u w=0.72u m=1
M7 Y A1 N_24 VDD mp5  l=0.42u w=0.96u m=1
M8 N_13 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_24 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y C0 N_25 VDD mp5  l=0.42u w=0.96u m=1
M11 Y B1 N_13 VDD mp5  l=0.42u w=0.96u m=1
M12 VDD C1 N_25 VDD mp5  l=0.42u w=0.96u m=1
.ends oai222d2
* SPICE INPUT		Wed Jul 10 13:52:39 2019	oai22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d0
.subckt oai22d0 A0 A1 B1 B0 GND VDD Y
M1 Y B0 N_7 GND mn5  l=0.5u w=0.5u m=1
M2 Y B1 N_7 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_11 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M7 Y A1 N_10 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai22d0
* SPICE INPUT		Wed Jul 10 13:52:46 2019	oai22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d1
.subckt oai22d1 A1 A0 B0 B1 VDD Y GND
M1 Y B1 N_7 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B0 Y GND mn5  l=0.5u w=0.58u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_7 A1 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_11 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M6 N_11 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_10 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y A1 N_10 VDD mp5  l=0.42u w=0.76u m=1
.ends oai22d1
* SPICE INPUT		Wed Jul 10 13:52:53 2019	oai22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d2
.subckt oai22d2 A1 A0 B0 B1 VDD Y GND
M1 Y B1 N_7 GND mn5  l=0.5u w=0.72u m=1
M2 N_7 B0 Y GND mn5  l=0.5u w=0.72u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_7 A1 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_11 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M6 N_11 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_10 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y A1 N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends oai22d2
* SPICE INPUT		Wed Jul 10 13:53:00 2019	oai311d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai311d0
.subckt oai311d0 VDD Y GND C0 B0 A0 A1 A2
M1 N_11 A2 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_20 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_20 GND mn5  l=0.5u w=0.5u m=1
M6 N_7 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M7 N_8 A1 N_7 VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 VDD C0 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oai311d0
* SPICE INPUT		Wed Jul 10 13:53:07 2019	oai311d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai311d1
.subckt oai311d1 C0 A2 A1 A0 B0 VDD Y GND
M1 N_9 B0 N_18 GND mn5  l=0.5u w=0.58u m=1
M2 N_9 A0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 A1 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_9 A2 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y C0 N_18 GND mn5  l=0.5u w=0.58u m=1
M6 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_12 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_12 A1 N_11 VDD mp5  l=0.42u w=0.76u m=1
M9 N_11 A2 Y VDD mp5  l=0.42u w=0.76u m=1
M10 VDD C0 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai311d1
* SPICE INPUT		Wed Jul 10 13:53:14 2019	oai311d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai311d2
.subckt oai311d2 A0 B0 C0 A1 A2 Y VDD GND
M1 N_10 A2 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_10 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y C0 N_11 GND mn5  l=0.5u w=0.72u m=1
M4 N_10 B0 N_11 GND mn5  l=0.5u w=0.72u m=1
M5 N_10 A0 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_17 A2 Y VDD mp5  l=0.42u w=0.96u m=1
M7 N_18 A1 N_17 VDD mp5  l=0.42u w=0.96u m=1
M8 VDD C0 Y VDD mp5  l=0.42u w=0.96u m=1
M9 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_18 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oai311d2
* SPICE INPUT		Wed Jul 10 13:53:21 2019	oai31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d0
.subckt oai31d0 A2 A0 A1 B0 Y VDD GND
M1 Y B0 N_7 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_11 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 A0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A2 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oai31d0
* SPICE INPUT		Wed Jul 10 13:53:29 2019	oai31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d1
.subckt oai31d1 A2 A0 A1 B0 Y VDD GND
M1 Y B0 N_7 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_7 A2 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 N_11 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_11 A0 N_10 VDD mp5  l=0.42u w=0.76u m=1
M8 N_10 A2 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai31d1
* SPICE INPUT		Wed Jul 10 13:53:36 2019	oai31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d2
.subckt oai31d2 A2 B0 A0 A1 GND VDD Y
M1 N_8 A1 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B0 N_8 GND mn5  l=0.5u w=0.72u m=1
M4 N_8 A2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_15 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_15 A0 N_14 VDD mp5  l=0.42u w=0.96u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_14 A2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai31d2
* SPICE INPUT		Wed Jul 10 13:53:43 2019	oai321d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai321d0
.subckt oai321d0 B1 B0 A0 A1 A2 C0 VDD Y GND
M1 Y C0 N_10 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A2 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_10 B1 N_11 GND mn5  l=0.5u w=0.5u m=1
M7 N_17 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_19 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_19 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M12 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai321d0
* SPICE INPUT		Wed Jul 10 13:53:50 2019	oai321d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai321d1
.subckt oai321d1 A2 A1 A0 B0 B1 C0 GND Y VDD
M1 Y C0 N_11 GND mn5  l=0.5u w=0.58u m=1
M2 N_11 B1 N_10 GND mn5  l=0.5u w=0.58u m=1
M3 N_10 B0 N_11 GND mn5  l=0.5u w=0.58u m=1
M4 N_10 A0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_10 A1 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_10 A2 GND GND mn5  l=0.5u w=0.58u m=1
M7 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_15 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M9 N_15 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 N_14 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M11 N_14 A1 N_13 VDD mp5  l=0.42u w=0.76u m=1
M12 N_13 A2 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai321d1
* SPICE INPUT		Wed Jul 10 13:53:57 2019	oai321d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai321d2
.subckt oai321d2 A2 B0 B1 A1 A0 C0 GND Y VDD
M1 Y C0 N_9 GND mn5  l=0.5u w=0.72u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_8 B1 N_9 GND mn5  l=0.5u w=0.72u m=1
M5 N_8 B0 N_9 GND mn5  l=0.5u w=0.72u m=1
M6 N_8 A2 GND GND mn5  l=0.5u w=0.72u m=1
M7 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_14 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_14 A1 N_13 VDD mp5  l=0.42u w=0.96u m=1
M10 N_15 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M11 N_15 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_13 A2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai321d2
* SPICE INPUT		Wed Jul 10 13:54:05 2019	oai322d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai322d0
.subckt oai322d0 VDD Y GND B0 A0 A1 A2 B1 C0 C1
M1 N_11 B0 N_13 GND mn5  l=0.5u w=0.5u m=1
M2 Y C1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 C0 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_13 B1 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_13 A2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_13 A1 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 A0 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_8 C1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y C0 N_8 VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M11 Y A2 N_9 VDD mp5  l=0.42u w=0.52u m=1
M12 N_10 A1 N_9 VDD mp5  l=0.42u w=0.52u m=1
M13 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_3 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai322d0
* SPICE INPUT		Wed Jul 10 13:54:13 2019	oai322d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai322d1
.subckt oai322d1 Y VDD GND B0 A0 A1 A2 B1 C0 C1
M1 N_14 B0 N_12 GND mn5  l=0.5u w=0.58u m=1
M2 Y C1 N_12 GND mn5  l=0.5u w=0.58u m=1
M3 N_12 C0 Y GND mn5  l=0.5u w=0.58u m=1
M4 N_14 B1 N_12 GND mn5  l=0.5u w=0.58u m=1
M5 N_14 A2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_14 A1 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_14 A0 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_9 C1 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_9 C0 Y VDD mp5  l=0.42u w=0.76u m=1
M10 N_3 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M11 N_10 A2 Y VDD mp5  l=0.42u w=0.76u m=1
M12 N_11 A1 N_10 VDD mp5  l=0.42u w=0.76u m=1
M13 N_11 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M14 N_3 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oai322d1
* SPICE INPUT		Wed Jul 10 13:54:20 2019	oai322d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai322d2
.subckt oai322d2 GND Y VDD A1 C1 A0 A2 B0 B1 C0
M1 N_3 B0 N_2 GND mn5  l=0.5u w=0.72u m=1
M2 N_2 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y C1 N_3 GND mn5  l=0.5u w=0.72u m=1
M4 N_2 B1 N_3 GND mn5  l=0.5u w=0.72u m=1
M5 N_2 A2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_3 C0 Y GND mn5  l=0.5u w=0.72u m=1
M7 N_2 A1 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_26 C1 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_12 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M10 N_26 C0 Y VDD mp5  l=0.42u w=0.96u m=1
M11 N_12 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_28 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 N_27 A2 Y VDD mp5  l=0.42u w=0.96u m=1
M14 N_28 A1 N_27 VDD mp5  l=0.42u w=0.96u m=1
.ends oai322d2
* SPICE INPUT		Wed Jul 10 13:54:27 2019	oai32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d0
.subckt oai32d0 A0 B1 A1 A2 B0 Y VDD GND
M1 N_7 B0 Y GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A2 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 B1 Y GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_16 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_17 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y B1 N_15 VDD mp5  l=0.42u w=0.52u m=1
M10 N_17 A0 N_16 VDD mp5  l=0.42u w=0.52u m=1
.ends oai32d0
* SPICE INPUT		Wed Jul 10 13:54:34 2019	oai32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d1
.subckt oai32d1 A2 B1 B0 A0 A1 GND VDD Y
M1 N_9 A1 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 A0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 B0 Y GND mn5  l=0.5u w=0.58u m=1
M4 N_9 B1 Y GND mn5  l=0.5u w=0.58u m=1
M5 N_9 A2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_13 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_13 A0 N_12 VDD mp5  l=0.42u w=0.76u m=1
M8 N_11 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y B1 N_11 VDD mp5  l=0.42u w=0.76u m=1
M10 N_12 A2 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai32d1
* SPICE INPUT		Wed Jul 10 13:54:41 2019	oai32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d2
.subckt oai32d2 A2 B1 B0 A0 A1 GND VDD Y
M1 N_9 A1 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 B0 Y GND mn5  l=0.5u w=0.72u m=1
M4 N_9 B1 Y GND mn5  l=0.5u w=0.72u m=1
M5 N_9 A2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_13 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_13 A0 N_12 VDD mp5  l=0.42u w=0.96u m=1
M8 N_11 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y B1 N_11 VDD mp5  l=0.42u w=0.96u m=1
M10 N_12 A2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai32d2
* SPICE INPUT		Wed Jul 10 13:54:49 2019	oai33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d0
.subckt oai33d0 VDD Y GND B2 B1 B0 A1 A0 A2
M1 Y B0 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B2 N_12 GND mn5  l=0.5u w=0.5u m=1
M6 Y B1 N_12 GND mn5  l=0.5u w=0.5u m=1
M7 N_9 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_8 A0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M10 N_7 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M11 Y B2 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_9 B1 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends oai33d0
* SPICE INPUT		Wed Jul 10 13:54:56 2019	oai33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d1
.subckt oai33d1 VDD Y GND B2 B1 B0 A1 A0 A2
M1 Y B0 N_12 GND mn5  l=0.5u w=0.58u m=1
M2 N_12 A1 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_12 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_12 A2 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y B2 N_12 GND mn5  l=0.5u w=0.58u m=1
M6 Y B1 N_12 GND mn5  l=0.5u w=0.58u m=1
M7 N_9 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_8 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_8 A0 N_7 VDD mp5  l=0.42u w=0.76u m=1
M10 N_7 A2 Y VDD mp5  l=0.42u w=0.76u m=1
M11 Y B2 N_6 VDD mp5  l=0.42u w=0.76u m=1
M12 N_9 B1 N_6 VDD mp5  l=0.42u w=0.76u m=1
.ends oai33d1
* SPICE INPUT		Wed Jul 10 13:55:03 2019	oai33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d2
.subckt oai33d2 VDD Y GND B2 B1 B0 A1 A0 A2
M1 N_14 A2 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_14 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B1 N_14 GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 N_14 GND mn5  l=0.5u w=0.72u m=1
M5 N_14 A1 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y B2 N_14 GND mn5  l=0.5u w=0.72u m=1
M7 N_7 A2 Y VDD mp5  l=0.42u w=0.96u m=1
M8 N_8 A0 N_7 VDD mp5  l=0.42u w=0.96u m=1
M9 N_9 B1 N_6 VDD mp5  l=0.42u w=0.96u m=1
M10 N_9 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 N_8 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 Y B2 N_6 VDD mp5  l=0.42u w=0.96u m=1
.ends oai33d2
* SPICE INPUT		Wed Jul 10 13:55:10 2019	oaim211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim211d0
.subckt oaim211d0 B0 C0 A0N A1N GND VDD Y
M1 N_11 A1N N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y C0 N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim211d0
* SPICE INPUT		Wed Jul 10 13:55:17 2019	oaim211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim211d1
.subckt oaim211d1 GND Y VDD C0 B0 A0N A1N
M1 N_7 A1N N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A0N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 N_4 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_8 B0 N_6 GND mn5  l=0.5u w=0.58u m=1
M5 Y C0 N_6 GND mn5  l=0.5u w=0.58u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oaim211d1
* SPICE INPUT		Wed Jul 10 13:55:25 2019	oaim211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim211d2
.subckt oaim211d2 GND Y VDD B0 C0 A0N A1N
M1 N_7 A1N N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A0N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C0 N_6 GND mn5  l=0.5u w=0.72u m=1
M5 N_8 B0 N_6 GND mn5  l=0.5u w=0.72u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oaim211d2
* SPICE INPUT		Wed Jul 10 13:55:32 2019	oaim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d0
.subckt oaim21d0 B0 A1N A0N VDD GND Y
M1 N_10 A0N N_3 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 N_9 GND mn5  l=0.5u w=0.5u m=1
M4 N_9 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim21d0
* SPICE INPUT		Wed Jul 10 13:55:39 2019	oaim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d1
.subckt oaim21d1 B0 A1N A0N VDD GND Y
M1 N_10 A0N N_3 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 N_9 GND mn5  l=0.5u w=0.58u m=1
M4 N_9 B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_3 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oaim21d1
* SPICE INPUT		Wed Jul 10 13:55:46 2019	oaim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d2
.subckt oaim21d2 B0 A1N A0N VDD GND Y
M1 N_10 A0N N_3 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 N_9 GND mn5  l=0.5u w=0.72u m=1
M4 N_9 B0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_3 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oaim21d2
* SPICE INPUT		Wed Jul 10 13:55:53 2019	oaim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d0
.subckt oaim22d0 B1 B0 A0N A1N Y VDD GND
M1 N_11 A1N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A0N N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 N_4 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_7 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_7 B1 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_18 B1 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oaim22d0
* SPICE INPUT		Wed Jul 10 13:56:00 2019	oaim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d1
.subckt oaim22d1 B1 B0 A0N A1N Y VDD GND
M1 N_11 A1N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A0N N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 N_4 Y GND mn5  l=0.5u w=0.58u m=1
M4 N_7 B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_7 B1 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_18 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 N_18 B1 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oaim22d1
* SPICE INPUT		Wed Jul 10 13:56:08 2019	oaim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d2
.subckt oaim22d2 B1 B0 A0N A1N Y VDD GND
M1 N_11 A1N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A0N N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 N_4 Y GND mn5  l=0.5u w=0.72u m=1
M4 N_7 B0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_7 B1 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_18 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_18 B1 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oaim22d2
* SPICE INPUT		Wed Jul 10 13:56:15 2019	oaim2m11d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim2m11d0
.subckt oaim2m11d0 C0 A0N B0N A1N VDD GND Y
M1 N_11 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_12 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A0N N_12 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_11 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_7 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B0N N_7 VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim2m11d0
* SPICE INPUT		Wed Jul 10 13:56:22 2019	oaim2m11d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim2m11d1
.subckt oaim2m11d1 C0 A0N B0N A1N VDD GND Y
M1 N_11 N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_12 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A0N N_12 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_11 GND mn5  l=0.5u w=0.58u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_7 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B0N N_7 VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oaim2m11d1
* SPICE INPUT		Wed Jul 10 13:56:30 2019	oaim2m11d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim2m11d2
.subckt oaim2m11d2 C0 B0N A1N A0N VDD Y GND
M1 N_3 A0N N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 B0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y C0 N_11 GND mn5  l=0.5u w=0.72u m=1
M6 N_9 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 B0N N_9 VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oaim2m11d2
* SPICE INPUT		Wed Jul 10 13:56:37 2019	oaim31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim31d0
.subckt oaim31d0 GND Y VDD A1N A2N B0 A0N
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1N N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0N N_4 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A2N VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim31d0
* SPICE INPUT		Wed Jul 10 13:56:44 2019	oaim31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim31d1
.subckt oaim31d1 GND Y VDD A1N A2N A0N B0
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.58u m=1
M2 N_6 B0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_8 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1N N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0N N_4 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_4 A2N VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim31d1
* SPICE INPUT		Wed Jul 10 13:56:51 2019	oaim31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim31d2
.subckt oaim31d2 GND Y VDD A1N A2N B0 A0N
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.72u m=1
M2 N_6 B0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_8 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1N N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0N N_4 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_4 A2N VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim31d2
* SPICE INPUT		Wed Jul 10 13:56:58 2019	or02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d0
.subckt or02d0 A B VDD GND Y
M1 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 B N_3 VDD mp5  l=0.42u w=0.52u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or02d0
* SPICE INPUT		Wed Jul 10 13:57:05 2019	or02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d1
.subckt or02d1 A B VDD GND Y
M1 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_12 B N_2 VDD mp5  l=0.42u w=0.52u m=1
M5 N_12 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends or02d1
* SPICE INPUT		Wed Jul 10 13:57:12 2019	or02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d2
.subckt or02d2 A B GND VDD Y
M1 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 B N_3 VDD mp5  l=0.42u w=0.52u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or02d2
* SPICE INPUT		Wed Jul 10 13:57:20 2019	or03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d0
.subckt or03d0 B A C GND VDD Y
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_13 C N_3 VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_14 B N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends or03d0
* SPICE INPUT		Wed Jul 10 13:57:27 2019	or03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d1
.subckt or03d1 B A C GND VDD Y
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_13 C N_3 VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_14 B N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends or03d1
* SPICE INPUT		Wed Jul 10 13:57:34 2019	or03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d2
.subckt or03d2 B A C GND VDD Y
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_13 C N_3 VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_14 B N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends or03d2
* SPICE INPUT		Wed Jul 10 13:57:41 2019	or04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d0
.subckt or04d0 A B D C VDD Y GND
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_14 D N_3 VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_16 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or04d0
* SPICE INPUT		Wed Jul 10 13:57:48 2019	or04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d1
.subckt or04d1 D A C B VDD Y GND
M1 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 D GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_14 D N_2 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends or04d1
* SPICE INPUT		Wed Jul 10 13:57:55 2019	or04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d2
.subckt or04d2 D A B C VDD Y GND
M1 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 D GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_15 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_14 D N_2 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends or04d2
* SPICE INPUT		Wed Jul 10 13:58:03 2019	or12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or12d0
.subckt or12d0 B AN VDD GND Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_14 B N_2 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or12d0
* SPICE INPUT		Wed Jul 10 13:58:10 2019	or12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or12d1
.subckt or12d1 AN B Y VDD GND
M1 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_2 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_14 B N_4 VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_2 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_14 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or12d1
* SPICE INPUT		Wed Jul 10 13:58:17 2019	or12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or12d2
.subckt or12d2 AN B Y VDD GND
M1 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_14 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 B N_2 VDD mp5  l=0.42u w=0.52u m=1
M7 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends or12d2
* SPICE INPUT		Wed Jul 10 13:58:24 2019	or13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or13d0
.subckt or13d0 C B AN Y VDD GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_15 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C N_16 VDD mp5  l=0.42u w=0.52u m=1
.ends or13d0
* SPICE INPUT		Wed Jul 10 13:58:32 2019	or13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or13d1
.subckt or13d1 AN C B GND VDD Y
M1 N_5 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_5 B GND GND mn5  l=0.5u w=0.5u m=1
M4 N_5 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 C N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or13d1
* SPICE INPUT		Wed Jul 10 13:58:39 2019	or13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or13d2
.subckt or13d2 C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 C N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends or13d2
* SPICE INPUT		Wed Jul 10 13:58:46 2019	or23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or23d0
.subckt or23d0 AN C BN Y VDD GND
M1 N_6 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 BN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_3 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_18 N_7 N_17 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C N_18 VDD mp5  l=0.42u w=0.52u m=1
M11 N_17 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_3 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or23d0
* SPICE INPUT		Wed Jul 10 13:58:53 2019	or23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or23d1
.subckt or23d1 AN C BN Y VDD GND
M1 N_5 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_5 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_2 C N_18 VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 N_5 N_17 VDD mp5  l=0.42u w=0.52u m=1
M10 N_17 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends or23d1
* SPICE INPUT		Wed Jul 10 13:59:00 2019	or23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or23d2
.subckt or23d2 BN C AN Y VDD GND
M1 N_6 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 BN GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_6 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_17 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 N_5 N_17 VDD mp5  l=0.42u w=0.52u m=1
M10 N_2 C N_18 VDD mp5  l=0.42u w=0.52u m=1
M11 N_5 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends or23d2
* SPICE INPUT		Wed Jul 10 13:59:08 2019	ora211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d0
.subckt ora211d0 C0 B0 A1 A0 GND Y VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_6 C0 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_17 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora211d0
* SPICE INPUT		Wed Jul 10 13:59:15 2019	ora211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d1
.subckt ora211d1 A1 B0 C0 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_5 C0 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A1 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_5 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
.ends ora211d1
* SPICE INPUT		Wed Jul 10 13:59:22 2019	ora211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d2
.subckt ora211d2 A1 B0 C0 A0 VDD Y GND
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_5 C0 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A1 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_5 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
.ends ora211d2
* SPICE INPUT		Wed Jul 10 13:59:30 2019	ora21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d0
.subckt ora21d0 B0 A1 A0 Y VDD GND
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_6 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B0 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_5 A1 N_14 VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora21d0
* SPICE INPUT		Wed Jul 10 13:59:37 2019	ora21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d1
.subckt ora21d1 B0 A1 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 N_9 GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_14 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 A1 N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends ora21d1
* SPICE INPUT		Wed Jul 10 13:59:44 2019	ora21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d2
.subckt ora21d2 A1 B0 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_4 B0 N_9 GND mn5  l=0.5u w=0.5u m=1
M4 N_9 A1 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_14 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_4 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A1 N_14 VDD mp5  l=0.42u w=0.52u m=1
.ends ora21d2
* SPICE INPUT		Wed Jul 10 13:59:51 2019	ora311d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora311d1
.subckt ora311d1 C0 B0 A2 A1 A0 Y VDD GND
M1 Y N_7 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 B0 N_12 GND mn5  l=0.5u w=0.5u m=1
M6 N_12 C0 N_7 GND mn5  l=0.5u w=0.5u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_19 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_19 A1 N_18 VDD mp5  l=0.42u w=0.52u m=1
M10 N_18 A2 N_7 VDD mp5  l=0.42u w=0.52u m=1
M11 N_7 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_7 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora311d1
* SPICE INPUT		Wed Jul 10 13:59:58 2019	ora311d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora311d2
.subckt ora311d2 A0 A1 A2 B0 C0 Y VDD GND
M1 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_12 C0 N_7 GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B0 N_12 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_7 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_18 A2 N_7 VDD mp5  l=0.42u w=0.52u m=1
M11 N_19 A1 N_18 VDD mp5  l=0.42u w=0.52u m=1
M12 N_19 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora311d2
* SPICE INPUT		Wed Jul 10 14:00:06 2019	ora31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d0
.subckt ora31d0 B0 A2 A0 A1 Y VDD GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 B0 N_7 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 A0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A2 N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora31d0
* SPICE INPUT		Wed Jul 10 14:00:13 2019	ora31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d1
.subckt ora31d1 A0 A2 B0 A1 GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_10 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_15 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A2 N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_16 A0 N_15 VDD mp5  l=0.42u w=0.52u m=1
.ends ora31d1
* SPICE INPUT		Wed Jul 10 14:00:20 2019	ora31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d2
.subckt ora31d2 A0 A2 B0 A1 GND VDD Y
M1 N_10 A1 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_5 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_5 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 A2 N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_16 A0 N_15 VDD mp5  l=0.42u w=0.52u m=1
.ends ora31d2


* Hierarchy Level 0

* Top of hierarchy  cell=xn02d0
.subckt xn02d0 VDD Y GND A B
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_8 A N_6 VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends xn02d0
* SPICE INPUT		Wed Jul 10 14:05:12 2019	xn02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d1
.subckt xn02d1 VDD Y GND A B
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_8 A N_6 VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends xn02d1
* SPICE INPUT		Wed Jul 10 14:05:19 2019	xn02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d2
.subckt xn02d2 VDD Y GND A B
M1 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A N_4 GND mn5  l=0.5u w=0.5u m=1
M6 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_7 N_5 N_4 VDD mp5  l=0.42u w=0.52u m=1
M11 N_8 A N_7 VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends xn02d2
* SPICE INPUT		Wed Jul 10 14:05:26 2019	xn03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d0
.subckt xn03d0 VDD Y GND C B A
M1 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M8 Y N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_9 C N_12 GND mn5  l=0.5u w=0.5u m=1
M11 N_12 N_11 N_6 GND mn5  l=0.5u w=0.5u m=1
M12 N_11 C VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.52u m=1
M16 N_9 B N_4 VDD mp5  l=0.42u w=0.52u m=1
M17 N_6 B N_5 VDD mp5  l=0.42u w=0.52u m=1
M18 N_10 B VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 C N_12 VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 N_11 N_12 VDD mp5  l=0.42u w=0.52u m=1
.ends xn03d0
* SPICE INPUT		Wed Jul 10 14:05:34 2019	xn03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d1
.subckt xn03d1 VDD Y GND C A B
M1 N_12 N_11 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_9 C N_12 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M6 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M8 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M10 Y N_12 GND GND mn5  l=0.5u w=0.58u m=1
M11 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M12 N_11 C VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_9 B N_4 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 B N_5 VDD mp5  l=0.42u w=0.52u m=1
M15 N_10 B VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 C N_12 VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 N_11 N_12 VDD mp5  l=0.42u w=0.52u m=1
.ends xn03d1
* SPICE INPUT		Wed Jul 10 14:05:41 2019	xn03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d2
.subckt xn03d2 VDD Y GND C A B
M1 N_12 N_11 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_9 C N_12 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M6 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M8 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M10 Y N_12 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M12 N_11 C VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_9 B N_4 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 B N_5 VDD mp5  l=0.42u w=0.52u m=1
M15 N_10 B VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 C N_12 VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 N_11 N_12 VDD mp5  l=0.42u w=0.52u m=1
.ends xn03d2
* SPICE INPUT		Wed Jul 10 14:05:48 2019	xr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d0
.subckt xr02d0 VDD Y GND B A
M1 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_6 N_5 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_4 A N_6 VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_8 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends xr02d0
* SPICE INPUT		Wed Jul 10 14:05:55 2019	xr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d1
.subckt xr02d1 VDD Y GND B A
M1 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_6 N_5 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_4 A N_6 VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M11 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_8 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends xr02d1
* SPICE INPUT		Wed Jul 10 14:06:02 2019	xr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d2
.subckt xr02d2 VDD Y GND B A
M1 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A N_7 GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_5 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_7 A N_4 VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_8 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
.ends xr02d2
* SPICE INPUT		Wed Jul 10 14:06:10 2019	xr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d0
.subckt xr03d0 VDD Y GND C B A
M1 N_9 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 C N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M9 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M10 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M11 Y N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_4 A VDD VDD mp5  l=0.42u w=0.5u m=1
M13 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M14 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.5u m=1
M15 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.5u m=1
M16 N_9 B N_4 VDD mp5  l=0.42u w=0.5u m=1
M17 N_6 B N_5 VDD mp5  l=0.42u w=0.5u m=1
M18 N_10 B VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_11 C VDD VDD mp5  l=0.42u w=0.5u m=1
M20 Y N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 N_11 N_12 VDD mp5  l=0.42u w=0.5u m=1
M22 N_9 C N_12 VDD mp5  l=0.42u w=0.5u m=1
.ends xr03d0
* SPICE INPUT		Wed Jul 10 14:06:17 2019	xr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d1
.subckt xr03d1 VDD Y GND C A B
M1 N_9 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 C N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 Y N_12 GND GND mn5  l=0.5u w=0.58u m=1
M9 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M12 N_9 B N_4 VDD mp5  l=0.42u w=0.5u m=1
M13 N_6 B N_5 VDD mp5  l=0.42u w=0.5u m=1
M14 N_10 B VDD VDD mp5  l=0.42u w=0.5u m=1
M15 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.5u m=1
M16 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.5u m=1
M17 Y N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 N_4 A VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_11 C VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_6 N_11 N_12 VDD mp5  l=0.42u w=0.5u m=1
M22 N_9 C N_12 VDD mp5  l=0.42u w=0.5u m=1
.ends xr03d1
* SPICE INPUT		Wed Jul 10 14:06:24 2019	xr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d2
.subckt xr03d2 VDD Y GND A B C
M1 N_9 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 C N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 Y N_12 GND GND mn5  l=0.5u w=0.72u m=1
M9 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M12 N_9 B N_4 VDD mp5  l=0.42u w=0.5u m=1
M13 N_6 B N_5 VDD mp5  l=0.42u w=0.5u m=1
M14 N_10 B VDD VDD mp5  l=0.42u w=0.5u m=1
M15 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.5u m=1
M16 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.5u m=1
M17 Y N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 N_4 A VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_11 C VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_6 N_11 N_12 VDD mp5  l=0.42u w=0.5u m=1
M22 N_9 C N_12 VDD mp5  l=0.42u w=0.5u m=1
.ends xr03d2
