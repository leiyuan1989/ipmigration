****Sub-Circuit for DGRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNHSV1 CK D Q QN RN VDD VSS
MM39 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM3 m c net43 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=250.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=250.00n L=60.00n
MM0 m pm VSS VPW N12LL W=340.00n L=60.00n
MM40 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM4 m cn net43 VNW P12LL W=500.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=330.00n L=60.00n
MM1 m pm VDD VNW P12LL W=500.00n L=60.00n
.ENDS DGRNHSV1
****Sub-Circuit for DGRNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNHSV2 CK D Q QN RN VDD VSS
MM39 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM3 m c net43 VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM40 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM4 m cn net43 VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=450.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS DGRNHSV2
****Sub-Circuit for DGRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNHSV4 CK D Q QN RN VDD VSS
MM39 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM3 m c net43 VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=360.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 m pm VSS VPW N12LL W=390.00n L=60.00n
MM40 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM4 m cn net43 VNW P12LL W=580.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=540.0n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=580.00n L=60.00n
.ENDS DGRNHSV4
****Sub-Circuit for DGRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNQHSV1 CK D Q RN VDD VSS
MM3 m c net43 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=250.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=250.00n L=60.00n
MM0 m pm VSS VPW N12LL W=340.00n L=60.00n
MM4 m cn net43 VNW P12LL W=500.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=330.00n L=60.00n
MM1 m pm VDD VNW P12LL W=500.00n L=60.00n
.ENDS DGRNQHSV1
****Sub-Circuit for DGRNQHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT DGRNQHSV2 CK D Q RN VDD VSS
MM3 m c net43 VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=270.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=270.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM4 m cn net43 VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=450.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=350.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS DGRNQHSV2
****Sub-Circuit for DGRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNQHSV4 CK D Q RN VDD VSS
MM3 m c net43 VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=340.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=270.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=270.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM4 m cn net43 VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.0n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=350.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS DGRNQHSV4
****Sub-Circuit for DGRSNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRSNHSV1 CK D Q QN RN SN VDD VSS
MM43 snn SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN net073 VSS VPW N12LL W=290.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=340.00n L=60.00n
MM42 net69 snn net_0162 VPW N12LL W=250.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=250.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=290.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=250.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=340.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=450.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=380.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=440.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=500.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=440.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=380.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=380.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=500.00n L=60.00n
.ENDS DGRSNHSV1
****Sub-Circuit for DGRSNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRSNHSV2 CK D Q QN RN SN VDD VSS
MM43 snn SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN net073 VSS VPW N12LL W=430.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=360.00n L=60.00n
MM42 net69 snn net_0162 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=430.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=360.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=450.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=650.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=650.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGRSNHSV2
****Sub-Circuit for DGRSNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRSNHSV4 CK D Q QN RN SN VDD VSS
MM43 snn SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN net073 VSS VPW N12LL W=860.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=360.00n L=60.00n
MM42 net69 snn net_0162 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=860.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=360.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=450.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=1.3u L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=1.3u L=60.00n
MM18 net063 net073 VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGRSNHSV4
****Sub-Circuit for DGSNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGSNHSV1 CK D Q QN SN VDD VSS
MM39 QN net073 VSS VPW N12LL W=290.00n L=60.00n
MM43 snn SN VSS VPW N12LL W=200.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=270.00n L=60.00n
MM42 net69 snn VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=290.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=250.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=270.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=440.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=440.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=300.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=440.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=440.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=400.00n L=60.00n
.ENDS DGSNHSV1
****Sub-Circuit for DGSNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGSNHSV2 CK D Q QN SN VDD VSS
MM39 QN net073 VSS VPW N12LL W=430.00n L=60.00n
MM43 snn SN VSS VPW N12LL W=200.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=350.00n L=60.00n
MM42 net69 snn VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=380.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=430.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=260.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=260.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=350.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=650.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=300.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=570.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=650.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGSNHSV2
****Sub-Circuit for DGSNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGSNHSV4 CK D Q QN SN VDD VSS
MM39 QN net073 VSS VPW N12LL W=860.00n L=60.00n
MM43 snn SN VSS VPW N12LL W=200.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=340.00n L=60.00n
MM42 net69 snn VSS VPW N12LL W=250.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=860.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=270.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=270.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=340.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=1.3u L=60.00n
MM44 snn SN VDD VNW P12LL W=300.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=1.3u L=60.00n
MM18 net063 net073 VDD VNW P12LL W=490.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGSNHSV4
****Sub-Circuit for DHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DHSV1 CK D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=290.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM43 QN s VDD VNW P12LL W=440.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DHSV1
****Sub-Circuit for DHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DHSV2 CK D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=430.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=640.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=640.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DHSV2
****Sub-Circuit for DHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DHSV4 CK D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 net43 c net_099 VPW N12LL W=300.00n L=60.00n m=2
MM40 net_099 m VSS VPW N12LL W=300.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM17 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 net43 cn net_0158 VNW P12LL W=450.00n L=60.00n m=2
MM41 net_0158 m VDD VNW P12LL W=450.00n L=60.00n m=2
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM18 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DHSV4
****Sub-Circuit for DQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DQHSV1 CK D Q VDD VSS
MM39 net43 c net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS DQHSV1
****Sub-Circuit for DQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DQHSV2 CK D Q VDD VSS
MM39 net43 c net_099 VPW N12LL W=430.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=290.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=290.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=440.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=440.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DQHSV2
****Sub-Circuit for DQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DQHSV4 CK D Q VDD VSS
MM39 net43 c net_099 VPW N12LL W=600.0n L=60.00n
MM40 net_099 m VSS VPW N12LL W=600.0n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=290.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=290.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=910.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=910.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=440.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=440.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DQHSV4
****Sub-Circuit for DRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNHSV1 CK D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DRNHSV1
****Sub-Circuit for DRNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNHSV2 CK D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNHSV2
****Sub-Circuit for DRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNHSV4 CK D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=330.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=330.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNHSV4
****Sub-Circuit for DRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNQHSV1 CK D Q RDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DRNQHSV1
****Sub-Circuit for DRNQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNQHSV2 CK D Q RDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNQHSV2
****Sub-Circuit for DRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNQHSV4 CK D Q RDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=330.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=330.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNQHSV4
****Sub-Circuit for DRSNHSV1, Mon May 30 16:01:10 CST 2011****
.SUBCKT DRSNHSV1 CK D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=290.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=220.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=220.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=360.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=440.00n L=60.00n
.ENDS DRSNHSV1
****Sub-Circuit for DRSNHSV2, Mon May 30 19:07:49 CST 2011****
.SUBCKT DRSNHSV2 CK D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=360.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=380.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=400.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=390.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=220.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=220.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=400.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=600.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=600.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=600.00n L=60.00n
.ENDS DRSNHSV2
****Sub-Circuit for DRSNHSV4, Mon May 30 19:07:49 CST 2011****
.SUBCKT DRSNHSV4 CK D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=360.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=410.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n m=2
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=320.00n L=60.00n m=2
MM40 net43 R net_0132 VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=220.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=220.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 s net43 VDD VNW P12LL W=600.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=650.00n L=60.00n m=2
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=290.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=290.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=630.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=650.00n L=60.00n
.ENDS DRSNHSV4
****Sub-Circuit for DSNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DSNHSV1 CK D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=400.00n L=60.00n
.ENDS DSNHSV1
****Sub-Circuit for DSNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DSNHSV2 CK D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=300.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=390.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS DSNHSV2
****Sub-Circuit for DSNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DSNHSV4 CK D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=780.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=780.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM38 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=570.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=910.00n L=60.00n
.ENDS DSNHSV4
****Sub-Circuit for DXHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DXHSV1 CK DA DB Q QN SA VDD VSS
MM33 m c net43 VPW N12LL W=350.00n L=60.00n
MM16 net_0144 DB VSS VPW N12LL W=350.00n L=60.00n
MM31 san SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=350.00n L=60.00n
MM19 QN s VSS VPW N12LL W=350.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=310.00n L=60.00n
MM3 net_0148 SA n43 VPW N12LL W=240.00n L=60.00n
MM7 net69 n43 VSS VPW N12LL W=310.00n L=60.00n
MM5 net_0144 san n43 VPW N12LL W=240.00n L=60.00n
MM2 net_0148 DA VSS VPW N12LL W=350.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM38 m cn net43 VNW P12LL W=440.00n L=60.00n
MM37 net_0144 DB VDD VNW P12LL W=440.00n L=60.00n
MM15 net_0148 DA VDD VNW P12LL W=440.00n L=60.00n
MM32 san SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM20 QN s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 n43 VDD VNW P12LL W=390.00n L=60.00n
MM4 net_0148 san n43 VNW P12LL W=300.00n L=60.00n
MM6 net_0144 SA n43 VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DXHSV1
****Sub-Circuit for DXHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DXHSV2 CK DA DB Q QN SA VDD VSS
MM5 net_0150 san n43 VPW N12LL W=240.00n L=60.00n
MM2 net_0138 DA VSS VPW N12LL W=350.00n L=60.00n
MM31 san SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM19 QN s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM33 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=310.00n L=60.00n
MM16 net_0150 DB VSS VPW N12LL W=350.00n L=60.00n
MM7 net69 n43 VSS VPW N12LL W=430.00n L=60.00n
MM3 net_0138 SA n43 VPW N12LL W=240.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM15 net_0138 DA VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0150 DB VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0138 san n43 VNW P12LL W=300.00n L=60.00n
MM6 net_0150 SA n43 VNW P12LL W=300.00n L=60.00n
MM32 san SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=550.00n L=60.00n
MM20 QN s VDD VNW P12LL W=550.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 m cn net43 VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 n43 VDD VNW P12LL W=550.00n L=60.00n
MM1 m pm VDD VNW P12LL W=550.00n L=60.00n
.ENDS DXHSV2
****Sub-Circuit for DXHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DXHSV4 CK DA DB Q QN SA VDD VSS
MM2 net_0156 DA VSS VPW N12LL W=350.00n L=60.00n
MM5 net_0144 san n43 VPW N12LL W=240.00n L=60.00n
MM3 net_0156 SA n43 VPW N12LL W=240.00n L=60.00n
MM16 net_0144 DB VSS VPW N12LL W=350.00n L=60.00n
MM31 san SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM19 QN s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM33 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=260.00n L=60.00n
MM7 net69 n43 VSS VPW N12LL W=260.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM6 net_0144 SA n43 VNW P12LL W=300.00n L=60.00n
MM4 net_0156 san n43 VNW P12LL W=300.00n L=60.00n
MM15 net_0156 DA VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0144 DB VDD VNW P12LL W=440.00n L=60.00n
MM32 san SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.1u L=60.00n
MM20 QN s VDD VNW P12LL W=1.1u L=60.00n
MM18 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM38 m cn net43 VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 n43 VDD VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=550.00n L=60.00n
.ENDS DXHSV4
****Sub-Circuit for EDGRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNHSV1 CK D E Q QN RN VDD VSS
MM43 QN s VSS VPW N12LL W=290.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=280.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=280.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM44 QN s VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNHSV1
****Sub-Circuit for EDGRNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNHSV2 CK D E Q QN RN VDD VSS
MM43 QN s VSS VPW N12LL W=390.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=390.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM44 QN s VDD VNW P12LL W=610.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=610.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=440.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNHSV2
****Sub-Circuit for EDGRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNHSV4 CK D E Q QN RN VDD VSS
MM43 QN s VSS VPW N12LL W=860.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=260.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=260.00n L=60.00n
MM44 QN s VDD VNW P12LL W=1.3u L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=500.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=400.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=400.00n L=60.00n
.ENDS EDGRNHSV4
****Sub-Circuit for EDGRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNQHSV1 CK D E Q RN VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=300.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=280.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=280.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=415.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNQHSV1
****Sub-Circuit for EDGRNQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNQHSV2 CK D E Q RN VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=420.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=420.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=440.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNQHSV2
****Sub-Circuit for EDGRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNQHSV4 CK D E Q RN VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=300.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.0n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=450.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=440.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNQHSV4
****Sub-Circuit for EDHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDHSV1 CK D E Q QN VDD VSS
MM43 QN s VSS VPW N12LL W=290.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=395.00n L=60.00n
MM42 QN s VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=495.00n L=60.00n
.ENDS EDHSV1
****Sub-Circuit for EDHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT EDHSV2 CK D E Q QN VDD VSS
MM43 QN s VSS VPW N12LL W=430.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=340.00n L=60.00n
MM42 QN s VDD VNW P12LL W=650.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=400.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=400.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=550.00n L=60.00n
.ENDS EDHSV2
****Sub-Circuit for EDHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDHSV4 CK D E Q QN VDD VSS
MM43 QN s VSS VPW N12LL W=860.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 QN s VDD VNW P12LL W=1.3u L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDHSV4
****Sub-Circuit for EDQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDQHSV1 CK D E Q VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=395.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=495.00n L=60.00n
.ENDS EDQHSV1
****Sub-Circuit for EDQHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT EDQHSV2 CK D E Q VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=340.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=400.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=400.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=550.00n L=60.00n
.ENDS EDQHSV2
****Sub-Circuit for EDQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDQHSV4 CK D E Q VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDQHSV4
****Sub-Circuit for EDRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNHSV1 CK D E Q QN RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM47 QN s VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM48 QN s VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=320.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=320.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNHSV1
****Sub-Circuit for EDRNHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT EDRNHSV2 CK D E Q QN RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM47 QN s VSS VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM48 QN s VDD VNW P12LL W=650.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=430.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=430.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNHSV2
****Sub-Circuit for EDRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNHSV4 CK D E Q QN RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM47 QN s VSS VPW N12LL W=860.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM48 QN s VDD VNW P12LL W=1.3u L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNHSV4
****Sub-Circuit for EDRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNQHSV1 CK D E Q RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=320.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=320.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNQHSV1
****Sub-Circuit for EDRNQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNQHSV2 CK D E Q RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=430.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=430.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNQHSV2
****Sub-Circuit for EDRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNQHSV4 CK D E Q RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNQHSV4



****Sub-Circuit for NDHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDHSV1 CKN D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=290.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM43 QN s VDD VNW P12LL W=440.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDHSV1
****Sub-Circuit for NDHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDHSV2 CKN D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=230.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=230.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=480.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDHSV2
****Sub-Circuit for NDHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDHSV4 CKN D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 net43 c net_099 VPW N12LL W=400.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=400.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM17 s net43 VSS VPW N12LL W=400.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 net43 cn net_0158 VNW P12LL W=450.00n L=60.00n m=2
MM41 net_0158 m VDD VNW P12LL W=450.00n L=60.00n m=2
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM18 s net43 VDD VNW P12LL W=600.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDHSV4
****Sub-Circuit for NDRNHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRNHSV1 CKN D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=200.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=200.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS NDRNHSV1
****Sub-Circuit for NDRNHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRNHSV2 CKN D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=200.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=300.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=200.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS NDRNHSV2
****Sub-Circuit for NDRNHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRNHSV4 CKN D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM3 net_0154 c net43 VPW N12LL W=360.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=200.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=190.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=280.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=280.00n L=60.00n m=2
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=190.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=190.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=260.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=560n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=650.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=610.00n L=60.00n
.ENDS NDRNHSV4
****Sub-Circuit for NDRSNHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRSNHSV1 CKN D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=200.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=200.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=380.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=440.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=350.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=440.00n L=60.00n
.ENDS NDRSNHSV1
****Sub-Circuit for NDRSNHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRSNHSV2 CKN D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=250.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=260.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=240.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=250.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=250.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=240.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=320.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=460.00n L=60.00n m=1
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=650.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=580.00n L=60.00n
.ENDS NDRSNHSV2
****Sub-Circuit for NDRSNHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRSNHSV4 CKN D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=260.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=240.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=420.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=240.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 s net43 VDD VNW P12LL W=470.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=460n L=60.00n
MM29 cn c VDD VNW P12LL W=640.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=650.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=430.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=620.00n L=60.00n
.ENDS NDRSNHSV4
****Sub-Circuit for NDSNHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDSNHSV1 CKN D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=290.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=270.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=290.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDSNHSV1
****Sub-Circuit for NDSNHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDSNHSV2 CKN D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=260.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=390.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=390.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=395.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=395.00n L=60.00n
.ENDS NDSNHSV2
****Sub-Circuit for NDSNHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDSNHSV4 CKN D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=390.00n L=60.00n
MM30 cn c VSS VPW N12LL W=400.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=400.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 s net43 VDD VNW P12LL W=580.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=600.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=600.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=620.00n L=60.00n
.ENDS NDSNHSV4