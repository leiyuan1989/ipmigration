//* No part of this file can be released without the consent of SMIC.
//************************************************************************************************************                                                                                                                                                   
//* SMIC 0.11um Mixed Signal 1P6M(1P5M, 1P7M, 1P8M) 1.2V/3.3V SPICE model (for SPECTRE only) //*                                                                                                                                                     
//************************************************************************************************************                                                                                                                                                   
//*                                                                                                                                                                                                                                                              
//* Release version    : 1.14                                                                                                                                                                                                                                     
//*                                                                                                                                                                                                                                                              
//* Release date       : 03/28/2016                                                                                                                                                                                                                              
//*                                                                                                                                                                                                                                                              
//* Simulation tool    : Cadence spectre V10.1.1                                                                                                                                                                                                 
//*                                                                                                                                                                                                                                                              
//*  Inductor   :                                                                                                                                                                                                                                                
//* *  *------------------------*-----------------------------------------------------------------------------------------------------*
//*    |  Turn, Radius & Width  |T=1~3 step 0.5,W=5~13.5um,R=1.7071*W+16.378~120um;T=3.5~5.0 step 0.5,W=5~8um,R=1.7071*W+16.378~120um |
//* *  *------------------------*-----------------------------------------------------------------------------------------------------*
//*    |        Model Name      |      diff_ind_rf_pgs_psub_n                       								  |            
//* *  *------------------------*-----------------------------------------------------------------------------------------------------*
simulator lang=spectre  insensitive=yes
subckt diff_ind_rf_pgs_psub_n (PLUS MINUS PSUB)
parameters r=6e-05 radius_=0.00833333*(r/1e-06-0) w=8e-06 w_=0.0666667*(w/1e-06-0) n=3  \
T0=(n==1.5) \
T1=(radius_>=0.416958) \
T2=(w_+7.291667e-01*radius_>=0.904432) \
T3=(w_>=0.6004) \
T4=(radius_>=0.416375) \
T5=(radius_>=0.708625) \
T6=(w_+7.291667e-01*radius_>=0.903207) \
T7=(w_>=0.5996) \
T8=(radius_>=0.708042) \
T9=(n==1) \
T10=(n==2.5) \
T11=(n==2) \
T12=(n==3.5) \
T13=(n==3) \
T14=(n==4.5) \
T15=(n==4) \
T16=(n==5) \
S0=T0*(1-T1)*(1-T2) \
noS0=(1-S0) \
S1=T0*(1-T3)*T4*(1-T5)*noS0 \
noS1=(1-S1)*noS0 \
S2=T0*T6*T7*(1-T5)*noS1 \
noS2=(1-S2)*noS1 \
S3=T0*(1-T3)*T8*noS2 \
noS3=(1-S3)*noS2 \
S4=T0*T8*T7*noS3 \
noS4=(1-S4)*noS3 \
S5=T9*(1-T1)*(1-T2)*noS4 \
noS5=(1-S5)*noS4 \
S6=T9*(1-T3)*T4*(1-T5)*noS5 \
noS6=(1-S6)*noS5 \
S7=T9*T6*T7*(1-T5)*noS6 \
noS7=(1-S7)*noS6 \
S8=T9*(1-T3)*T8*noS7 \
noS8=(1-S8)*noS7 \
S9=T9*T8*T7*noS8 \
noS9=(1-S9)*noS8 \
S10=T10*(1-T1)*(1-T2)*noS9 \
noS10=(1-S10)*noS9 \
S11=T10*(1-T3)*T4*(1-T5)*noS10 \
noS11=(1-S11)*noS10 \
S12=T10*T6*T7*(1-T5)*noS11 \
noS12=(1-S12)*noS11 \
S13=T10*(1-T3)*T8*noS12 \
noS13=(1-S13)*noS12 \
S14=T10*T8*T7*noS13 \
noS14=(1-S14)*noS13 \
S15=T11*(1-T1)*(1-T2)*noS14 \
noS15=(1-S15)*noS14 \
S16=T11*(1-T3)*T4*(1-T5)*noS15 \
noS16=(1-S16)*noS15 \
S17=T11*T6*T7*(1-T5)*noS16 \
noS17=(1-S17)*noS16 \
S18=T11*(1-T3)*T8*noS17 \
noS18=(1-S18)*noS17 \
S19=T11*T8*T7*noS18 \
noS19=(1-S19)*noS18 \
S20=T12*(1-T1)*noS19 \
noS20=(1-S20)*noS19 \
S21=T12*T4*(1-T5)*noS20 \
noS21=(1-S21)*noS20 \
S22=T12*T8*noS21 \
noS22=(1-S22)*noS21 \
S23=T13*(1-T1)*(1-T2)*noS22 \
noS23=(1-S23)*noS22 \
S24=T13*(1-T3)*T4*(1-T5)*noS23 \
noS24=(1-S24)*noS23 \
S25=T13*T6*T7*(1-T5)*noS24 \
noS25=(1-S25)*noS24 \
S26=T13*(1-T3)*T8*noS25 \
noS26=(1-S26)*noS25 \
S27=T13*T8*T7*noS26 \
noS27=(1-S27)*noS26 \
S28=T14*(1-T1)*noS27 \
noS28=(1-S28)*noS27 \
S29=T14*T4*(1-T5)*noS28 \
noS29=(1-S29)*noS28 \
S30=T14*T8*noS29 \
noS30=(1-S30)*noS29 \
S31=T15*(1-T1)*noS30 \
noS31=(1-S31)*noS30 \
S32=T15*T4*(1-T5)*noS31 \
noS32=(1-S32)*noS31 \
S33=T15*T8*noS32 \
noS33=(1-S33)*noS32 \
S34=T16*(1-T1)*noS33 \
noS34=(1-S34)*noS33 \
S35=T16*T4*(1-T5)*noS34 \
noS35=(1-S35)*noS34 \
S36=T16*T8*noS35 \
noS36=(1-S36)*noS35 \
V0_part1=0.000000e+00*S0+(-2.188913e+00)*S1+(-1.222321e+01)*S2+1.266025e+00*S3+(-8.910136e+00)*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V0_part2=V0_part1+2.850805e-01*S10+3.686949e+00*S11+5.663831e+00*S12+6.850846e+00*S13+(-2.980274e+01)*S14+(-4.343037e+00)*S15+(-4.894421e+00)*S16+(-2.723354e+00)*S17+(-3.417343e-01)*S18+(-2.290001e+00)*S19 \
V0_part3=V0_part2+2.577640e+00*S20+3.943746e+00*S21+(-2.586079e+00)*S22+1.638807e-01*S23+8.985351e+00*S24+0.000000e+00*S25+(-3.155055e+01)*S26+(-2.131377e+01)*S27+(-3.610296e+00)*S28+6.419885e+00*S29 \
V0=V0_part3+6.613859e+00*S30+4.907798e+00*S31+1.207101e+01*S32+(-1.543649e+01)*S33+(-4.671759e+00)*S34+1.444530e+01*S35+2.336190e+01*S36 \
V1_part1=0.000000e+00*S0+1.558597e+01*S1+2.929961e+01*S2+2.101637e+01*S3+1.952267e+01*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V1_part2=V1_part1+2.497215e+01*S10+2.300462e+01*S11+2.051031e+01*S12+2.237192e+01*S13+5.938577e+01*S14+3.223314e+01*S15+2.751532e+01*S16+2.771719e+01*S17+3.032280e+01*S18+2.337416e+01*S19 \
V1_part3=V1_part2+5.113689e+01*S20+4.788171e+01*S21+6.519320e+01*S22+6.032734e+01*S23+2.519095e+01*S24+0.000000e+00*S25+7.047157e+01*S26+4.684035e+01*S27+1.033268e+02*S28+7.632438e+01*S29 \
V1=V1_part3+7.604024e+01*S30+6.027022e+01*S31+5.376599e+01*S32+8.972297e+01*S33+1.222638e+02*S34+8.461609e+01*S35+7.985180e+01*S36 \
V2_part1=0.000000e+00*S0+(-1.934879e+00)*S1+6.221866e+00*S2+(-2.162807e+01)*S3+1.828117e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V2_part2=V2_part1+9.270080e-01*S10+(-8.996662e+00)*S11+(-9.583669e+00)*S12+(-1.874151e+01)*S13+1.457216e+01*S14+(-1.320362e+00)*S15+3.270971e-01*S16+(-3.943386e+00)*S17+(-2.762510e+01)*S18+(-2.911584e+00)*S19 \
V2_part3=V2_part2+2.686540e+00*S20+(-1.079198e+00)*S21+(-2.226540e+00)*S22+9.492091e-01*S23+(-1.809293e+01)*S24+0.000000e+00*S25+2.199950e+01*S26+1.947594e+01*S27+2.305971e+01*S28+2.291534e+00*S29 \
V2=V2_part3+(-3.729510e+00)*S30+(-1.742953e+00)*S31+(-2.173379e+01)*S32+1.805506e+00*S33+3.174499e+01*S34+(-1.871980e+01)*S35+(-3.992889e+01)*S36 \
V3_part1=3.382088e-01*S0+(-4.271846e-01)*S1+(-3.309507e-01)*S2+(-1.191771e+00)*S3+(-3.026173e-01)*S4+(-1.564318e-01)*S5+(-2.601445e-01)*S6+(-1.082656e-01)*S7+(-4.552855e-01)*S8+(-3.320446e-01)*S9 \
V3_part2=V3_part1+(-2.884163e-01)*S10+(-1.624855e+00)*S11+(-1.542167e-01)*S12+(-1.639843e+00)*S13+(-6.046250e-01)*S14+(-2.425435e-01)*S15+(-3.832261e-01)*S16+(-2.031645e-01)*S17+(-8.397946e-01)*S18+(-6.205529e-01)*S19 \
V3_part3=V3_part2+(-2.612782e-01)*S20+(-5.240519e-01)*S21+(-8.624852e+00)*S22+(-2.075498e-02)*S23+(-4.819097e-01)*S24+(-2.436149e-01)*S25+(-1.417964e+00)*S26+(-7.174262e-01)*S27+1.135721e+00*S28+(-4.561517e-01)*S29 \
V3=V3_part3+(-1.269719e+00)*S30+2.095714e-01*S31+(-4.305274e-01)*S32+(-8.070793e+00)*S33+(-2.101369e-01)*S34+(-5.985787e-01)*S35+(-1.434599e+00)*S36 \
V4_part1=1.082494e+00*S0+3.445881e+00*S1+3.498244e-01*S2+6.531851e-01*S3+7.761950e-01*S4+6.926253e-01*S5+7.132896e-01*S6+3.622430e-01*S7+8.167986e-01*S8+6.412253e-01*S9 \
V4_part2=V4_part1+(-3.657466e+00)*S10+1.527639e+00*S11+7.134715e-01*S12+(-1.884475e+00)*S13+1.408899e+00*S14+1.368132e+00*S15+1.462114e+00*S16+7.845700e-01*S17+1.492018e+00*S18+4.829800e-01*S19 \
V4_part3=V4_part2+1.976063e+00*S20+2.527356e+00*S21+1.188260e+00*S22+1.234614e+00*S23+2.207110e+00*S24+9.904278e-01*S25+(-1.246506e+00)*S26+1.849108e+00*S27+3.643818e+00*S28+3.146511e+00*S29 \
V4=V4_part3+3.948827e+00*S30+3.389348e+00*S31+2.794748e+00*S32+(-2.412462e-01)*S33+1.912805e+00*S34+3.474482e+00*S35+4.167145e+00*S36 \
V5_part1=8.515581e-02*S0+(-4.620254e-02)*S1+7.402240e-01*S2+1.609091e+00*S3+2.430989e-01*S4+5.956362e-02*S5+8.890476e-02*S6+7.903161e-02*S7+1.208175e-01*S8+1.169772e-01*S9 \
V5_part2=V5_part1+2.976188e+00*S10+1.822768e+00*S11+3.057848e-01*S12+4.855744e+00*S13+4.828337e-01*S14+1.244481e-01*S15+1.757368e-01*S16+1.924777e-01*S17+2.992184e-01*S18+1.152313e+00*S19 \
V5_part3=V5_part2+2.719205e-01*S20+2.951137e-01*S21+6.552327e+00*S22+9.794549e-01*S23+2.597345e-01*S24+3.192219e-01*S25+3.888535e+00*S26+5.476166e-01*S27+1.253428e+00*S28+3.501540e-01*S29 \
V5=V5_part3+4.928423e-01*S30+1.601172e+00*S31+3.017539e-01*S32+7.354509e+00*S33+1.854546e+00*S34+4.607935e-01*S35+6.002647e-01*S36 \
V6_part1=(-9.178359e-03)*S0+(-1.809311e-02)*S1+(-3.469446e-03)*S2+(-2.409103e-02)*S3+(-3.385986e-02)*S4+(-9.275531e-03)*S5+(-1.805718e-02)*S6+(-9.484982e-03)*S7+(-3.438445e-02)*S8+(-1.927470e-02)*S9 \
V6_part2=V6_part1+3.632143e-01*S10+(-9.597518e-03)*S11+(-3.454997e-02)*S12+3.443363e-01*S13+(-1.417962e-01)*S14+(-1.218714e-02)*S15+(-5.491354e-02)*S16+(-2.988085e-02)*S17+(-9.804144e-02)*S18+(-7.730735e-03)*S19 \
V6_part3=V6_part2+(-7.418317e-02)*S20+(-1.950086e-01)*S21+3.926309e-01*S22+(-3.502991e-02)*S23+(-1.204508e-01)*S24+(-6.806617e-02)*S25+3.257160e-01*S26+(-2.089747e-01)*S27+(-5.148758e-02)*S28+(-3.138669e-01)*S29 \
V6=V6_part3+(-5.716185e-01)*S30+(-3.768676e-02)*S31+(-2.365265e-01)*S32+3.884376e-01*S33+(-2.050724e-02)*S34+(-3.479937e-01)*S35+(-6.295238e-01)*S36 \
V7_part1=6.833163e-01*S0+7.561579e-01*S1+6.675984e-01*S2+8.339878e-01*S3+8.590395e-01*S4+3.163946e-01*S5+3.454767e-01*S6+3.068772e-01*S7+3.726964e-01*S8+3.456088e-01*S9 \
V7_part2=V7_part1+1.719641e+00*S10+1.824388e+00*S11+1.743307e+00*S12+1.831417e+00*S13+2.141787e+00*S14+9.694227e-01*S15+1.195592e+00*S16+1.060461e+00*S17+1.309719e+00*S18+1.091236e+00*S19 \
V7_part3=V7_part2+3.185151e+00*S20+3.533666e+00*S21+3.554583e+00*S22+2.106694e+00*S23+2.532385e+00*S24+2.236702e+00*S25+2.324928e+00*S26+2.741149e+00*S27+4.686802e+00*S28+5.529250e+00*S29 \
V7=V7_part3+6.193530e+00*S30+3.692982e+00*S31+4.233638e+00*S32+4.193925e+00*S33+5.381640e+00*S34+6.378476e+00*S35+7.119152e+00*S36 \
V8_part1=(-4.383708e-02)*S0+(-8.597002e-02)*S1+(-4.321802e-02)*S2+(-1.720254e-01)*S3+(-1.063938e-01)*S4+(-2.139286e-02)*S5+(-2.902345e-02)*S6+(-1.906875e-02)*S7+(-4.666726e-02)*S8+(-4.146824e-02)*S9 \
V8_part2=V8_part1+(-3.947516e-01)*S10+(-2.592933e-01)*S11+(-5.678236e-02)*S12+(-6.730331e-01)*S13+(-1.584772e-01)*S14+(-5.952370e-02)*S15+(-9.025088e-02)*S16+(-3.827326e-02)*S17+(-1.696063e-01)*S18+(-1.626632e-01)*S19 \
V8_part3=V8_part2+2.085043e-02*S20+2.096491e-02*S21+(-1.477562e+00)*S22+(-1.046401e-01)*S23+(-1.195593e-01)*S24+(-3.596326e-02)*S25+(-7.693320e-01)*S26+(-1.416558e-01)*S27+(-6.009981e-02)*S28+1.855852e-01*S29 \
V8=V8_part3+(-1.184776e-01)*S30+(-1.206864e-01)*S31+4.719416e-02*S32+(-1.524471e+00)*S33+(-8.566338e-02)*S34+2.481137e-01*S35+(-2.386518e-01)*S36 \
V9_part1=(-6.758253e-01)*S0+(-8.750606e-01)*S1+(-2.485939e-01)*S2+(-1.091367e+00)*S3+(-1.086963e+00)*S4+(-1.531793e-01)*S5+(-9.523292e-01)*S6+(-3.526650e-01)*S7+(-8.538565e-01)*S8+(-3.839888e-01)*S9 \
V9_part2=V9_part1+(-4.145268e-01)*S10+(-1.047160e+00)*S11+(-7.561890e-03)*S12+(-1.805322e+00)*S13+(-1.270891e+00)*S14+4.271534e-01*S15+(-2.659487e+00)*S16+(-1.127542e+00)*S17+(-2.332753e+00)*S18+(-1.050307e+00)*S19 \
V9_part3=V9_part2+(-1.888562e+00)*S20+(-1.349614e+01)*S21+(-2.259070e+00)*S22+(-6.137476e-01)*S23+(-4.461402e+00)*S24+(-1.177431e-01)*S25+(-2.247320e+00)*S26+(-1.552832e+00)*S27+(-7.676994e-01)*S28+(-1.610898e+01)*S29 \
V9=V9_part3+(-1.343332e+01)*S30+(-6.856369e-01)*S31+(-1.290856e+01)*S32+(-2.577915e+00)*S33+(-8.490440e-01)*S34+(-1.148649e+01)*S35+(-1.379285e+01)*S36 \
V10_part1=1.985890e+00*S0+9.545226e-01*S1+1.811707e+00*S2+1.932202e+00*S3+9.240795e-01*S4+(-1.848339e-01)*S5+3.368350e-01*S6+1.823905e-02*S7+(-4.263155e-01)*S8+3.986291e-02*S9 \
V10_part2=V10_part1+3.144473e+00*S10+3.563031e+00*S11+3.229059e+00*S12+3.091691e+00*S13+1.407929e+00*S14+(-3.169985e+00)*S15+1.849462e+00*S16+3.204414e-01*S17+2.950336e-02*S18+2.093796e+00*S19 \
V10_part3=V10_part2+9.682997e+00*S20+4.780046e+00*S21+5.164032e+00*S22+4.292168e+00*S23+3.617757e+00*S24+(-2.744105e-01)*S25+4.061435e+00*S26+1.712774e+00*S27+5.978439e+00*S28+5.490714e+00*S29 \
V10=V10_part3+3.472945e+00*S30+4.802567e+00*S31+6.584434e+00*S32+5.658433e+00*S33+7.649563e+00*S34+7.350689e+00*S35+4.648340e+00*S36 \
V11_part1=4.664570e-01*S0+8.251728e-01*S1+2.216757e-01*S2+5.138601e-01*S3+2.023354e+00*S4+6.271485e-01*S5+1.072014e+00*S6+1.161425e+00*S7+1.558678e+00*S8+1.086997e+00*S9 \
V11_part2=V11_part1+3.184116e-01*S10+5.582572e-01*S11+4.211039e+00*S12+8.056062e-01*S13+2.579952e+00*S14+2.307703e+00*S15+2.493685e+00*S16+3.200584e+00*S17+3.779531e+00*S18+6.862381e-01*S19 \
V11_part3=V11_part2+4.570256e+00*S20+9.537577e+00*S21+9.165855e-01*S22+4.357983e-01*S23+4.006873e+00*S24+6.437970e+00*S25+8.971227e-01*S26+2.599221e+00*S27+8.012144e-01*S28+1.181164e+01*S29 \
V11=V11_part3+1.042663e+01*S30+6.295279e-01*S31+8.637656e+00*S32+1.053254e+00*S33+7.814198e-01*S34+8.813074e+00*S35+1.069784e+01*S36 \
V12_part1=(-5.646991e-03)*S0+8.118506e-02*S1+(-1.227034e-02)*S2+(-1.186737e-01)*S3+(-1.625476e-02)*S4+3.335165e-03*S5+5.604596e-03*S6+1.054736e-02*S7+(-6.801009e-04)*S8+(-1.081705e-02)*S9 \
V12_part2=V12_part1+(-1.889167e-02)*S10+(-1.624207e-01)*S11+(-1.865629e-03)*S12+(-2.810779e-01)*S13+(-3.631755e-02)*S14+2.801820e-01*S15+(-2.813407e-02)*S16+7.638286e-02*S17+5.963018e-02*S18+(-1.667878e-01)*S19 \
V12_part3=V12_part2+(-7.780753e-02)*S20+3.761305e-01*S21+(-7.607695e-01)*S22+(-1.114816e-01)*S23+(-4.563381e-02)*S24+2.424058e-01*S25+(-3.771362e-01)*S26+(-8.224900e-02)*S27+(-1.762747e-01)*S28+5.253212e-01*S29 \
V12=V12_part3+5.674396e-01*S30+(-1.625236e-01)*S31+1.293946e-01*S32+(-8.188660e-01)*S33+(-2.661477e-01)*S34+1.381255e-02*S35+5.658013e-02*S36 \
V13_part1=1.545670e+00*S0+1.555944e+00*S1+1.487378e+00*S2+1.824851e+00*S3+1.515025e+00*S4+5.382520e-01*S5+5.966428e-01*S6+5.460831e-01*S7+6.299755e-01*S8+6.023586e-01*S9 \
V13_part2=V13_part1+3.231111e+00*S10+3.960172e+00*S11+3.421932e+00*S12+4.295828e+00*S13+3.616184e+00*S14+1.961994e+00*S15+2.165537e+00*S16+1.918596e+00*S17+2.289883e+00*S18+2.508926e+00*S19 \
V13_part3=V13_part2+6.342498e+00*S20+6.560658e+00*S21+7.930114e+00*S22+4.592601e+00*S23+4.657388e+00*S24+4.201294e+00*S25+5.498596e+00*S26+4.620085e+00*S27+9.991043e+00*S28+1.028386e+01*S29 \
V13=V13_part3+1.125094e+01*S30+7.670970e+00*S31+7.916265e+00*S32+9.446110e+00*S33+1.161675e+01*S34+1.192692e+01*S35+1.305156e+01*S36 \
V14_part1=(-1.164187e-01)*S0+(-2.910763e-01)*S1+(-8.472639e-02)*S2+(-2.829068e-01)*S3+(-2.184733e-01)*S4+(-4.964753e-02)*S5+(-9.542180e-02)*S6+(-4.975470e-02)*S7+(-1.298068e-01)*S8+(-8.198766e-02)*S9 \
V14_part2=V14_part1+(-1.767027e-01)*S10+(-2.482124e-01)*S11+(-1.910247e-01)*S12+(-5.515618e-01)*S13+(-4.951622e-01)*S14+(-3.312513e-01)*S15+(-3.063804e-01)*S16+(-1.938236e-01)*S17+(-5.600537e-01)*S18+(-2.124790e-01)*S19 \
V14_part3=V14_part2+(-2.483154e-01)*S20+(-1.562971e+00)*S21+(-4.299175e-01)*S22+(-8.660448e-02)*S23+(-6.541776e-01)*S24+(-3.852601e-01)*S25+(-6.346846e-01)*S26+(-5.822711e-01)*S27+3.303193e-01*S28+(-2.129807e+00)*S29 \
V14=V14_part3+(-3.613834e+00)*S30+1.089078e-01*S31+(-1.364143e+00)*S32+(-7.541026e-01)*S33+6.883644e-01*S34+(-1.361851e+00)*S35+(-3.112719e+00)*S36 \
V15_part1=3.852049e+00*S0+3.689209e+00*S1+6.274034e-01*S2+1.378736e+00*S3+1.891388e+00*S4+4.385865e-02*S5+(-8.369962e-02)*S6+2.784376e-01*S7+(-1.761560e+00)*S8+(-1.289785e+00)*S9 \
V15_part2=V15_part1+(-1.294789e-01)*S10+7.389699e-01*S11+7.322539e-01*S12+(-3.147867e-01)*S13+1.298601e+00*S14+(-1.418962e-01)*S15+5.704166e-01*S16+7.338866e-02*S17+(-1.231387e-01)*S18+9.286650e-01*S19 \
V15_part3=V15_part2+8.103033e-01*S20+(-3.145247e-01)*S21+(-4.297708e-01)*S22+9.386627e-01*S23+3.622025e-01*S24+8.090447e-02*S25+(-5.771549e-01)*S26+1.563673e+00*S27+1.187950e+00*S28+(-2.622908e-01)*S29 \
V15=V15_part3+(-3.688760e-01)*S30+7.715072e-01*S31+(-8.133342e-02)*S32+(-6.661839e-01)*S33+7.199981e-01*S34+7.097110e-01*S35+1.555650e-01*S36 \
V16_part1=(-1.407897e+00)*S0+(-7.714105e-01)*S1+1.523557e+00*S2+6.725178e-01*S3+(-1.675887e-01)*S4+2.958450e+00*S5+2.278677e+00*S6+1.257942e+00*S7+3.987252e+00*S8+3.669764e+00*S9 \
V16_part2=V16_part1+2.543869e+00*S10+1.458508e+00*S11+3.772085e-01*S12+1.317286e+00*S13+3.543203e-01*S14+3.852867e+00*S15+1.797758e+00*S16+1.567939e+00*S17+1.970192e+00*S18+6.621261e-01*S19 \
V16_part3=V16_part2+7.729232e-01*S20+2.017569e+00*S21+1.659762e+00*S22+1.482272e+00*S23+1.647716e+00*S24+1.106200e+00*S25+1.749144e+00*S26+2.089900e-01*S27+1.520128e+00*S28+1.939707e+00*S29 \
V16=V16_part3+2.059199e+00*S30+1.160851e+00*S31+1.985786e+00*S32+2.097422e+00*S33+2.072520e+00*S34+1.779016e+00*S35+2.323083e+00*S36 \
V17_part1=(-1.996081e+00)*S0+(-1.882683e+00)*S1+2.037182e+00*S2+(-1.427535e-01)*S3+7.656564e-01*S4+1.110008e+00*S5+1.089440e+00*S6+6.792394e-01*S7+1.713784e+00*S8+1.513722e+00*S9 \
V17_part2=V17_part1+1.271494e+00*S10+(-2.267441e-01)*S11+(-1.328657e-01)*S12+1.387605e-01*S13+(-1.483100e-02)*S14+1.280523e+00*S15+7.383108e-01*S16+2.452597e-01*S17+5.250735e-02*S18+3.906910e-02*S19 \
V17_part3=V17_part2+(-5.579494e-01)*S20+9.270595e-01*S21+6.294347e-01*S22+(-2.249989e-02)*S23+8.473955e-01*S24+1.044139e-01*S25+4.626887e-01*S26+(-6.805874e-02)*S27+(-8.566468e-01)*S28+1.168070e+00*S29 \
V17=V17_part3+7.288186e-01*S30+(-4.293945e-01)*S31+1.338553e+00*S32+8.763015e-01*S33+2.617258e-03*S34+4.043942e-02*S35+2.593425e-02*S36 \
V18_part1=(-1.406908e+00)*S0+(-8.234607e-01)*S1+(-9.568327e-02)*S2+(-1.412503e+00)*S3+(-8.281259e-01)*S4+(-1.198460e-02)*S5+1.491933e+00*S6+(-2.128034e+01)*S7+1.802392e+00*S8+1.683354e+00*S9 \
V18_part2=V18_part1+(-1.534031e+00)*S10+(-2.961085e+00)*S11+(-4.521273e+00)*S12+(-4.346002e+00)*S13+1.769887e+00*S14+1.052313e-01*S15+(-4.130523e-01)*S16+(-1.940281e+00)*S17+(-1.477554e+00)*S18+(-2.275629e+00)*S19 \
V18_part3=V18_part2+(-2.480659e+00)*S20+(-3.942189e+00)*S21+(-2.808569e+00)*S22+(-1.094926e+00)*S23+(-3.458240e+00)*S24+(-1.900145e+00)*S25+3.367659e+00*S26+2.163170e-01*S27+(-9.500672e-01)*S28+(-4.850446e+00)*S29 \
V18=V18_part3+(-6.959113e+00)*S30+(-2.685733e+00)*S31+(-4.467860e+00)*S32+(-1.851746e-02)*S33+(-9.812939e-01)*S34+(-5.745217e+00)*S35+(-8.253955e+00)*S36 \
V19_part1=8.237290e+00*S0+4.837152e+00*S1+3.347280e+00*S2+2.479039e+00*S3+4.085802e+00*S4+3.873746e+00*S5+(-3.156997e-01)*S6+3.751004e+01*S7+(-2.221536e-01)*S8+4.459656e-01*S9 \
V19_part2=V19_part1+8.638049e+00*S10+9.008084e+00*S11+1.231766e+01*S12+9.146378e+00*S13+3.277702e+00*S14+2.514278e+00*S15+3.046456e+00*S16+4.257060e+00*S17+1.993579e+00*S18+4.712812e+00*S19 \
V19_part3=V19_part2+1.080063e+01*S20+1.125224e+01*S21+6.773544e+00*S22+3.569312e+00*S23+1.005089e+01*S24+1.605102e+01*S25+1.659043e+00*S26+8.012115e+00*S27+8.148362e+00*S28+1.352925e+01*S29 \
V19=V19_part3+1.342689e+01*S30+1.146268e+01*S31+1.219032e+01*S32+4.533974e+00*S33+7.239029e+00*S34+1.455521e+01*S35+1.416593e+01*S36 \
V20_part1=4.200252e+00*S0+3.796446e+00*S1+3.328199e+00*S2+8.998533e+00*S3+5.272100e+00*S4+4.080515e+00*S5+3.239917e+00*S6+3.478093e+01*S7+2.462855e+00*S8+1.933770e+00*S9 \
V20_part2=V20_part1+7.194424e+00*S10+1.059705e+01*S11+1.050346e+01*S12+1.400711e+01*S13+7.476215e+00*S14+3.434202e+00*S15+4.686578e+00*S16+7.145367e+00*S17+1.125650e+01*S18+7.254425e+00*S19 \
V20_part3=V20_part2+1.120062e+01*S20+1.492410e+01*S21+1.695701e+01*S22+6.890498e+00*S23+1.197334e+01*S24+8.778336e+00*S25+5.990888e+00*S26+6.714826e+00*S27+1.011699e+01*S28+1.918733e+01*S29 \
V20=V20_part3+2.505166e+01*S30+1.258193e+01*S31+1.651052e+01*S32+1.480452e+01*S33+1.069515e+01*S34+2.167387e+01*S35+2.929427e+01*S36 \
V21_part1=2.745424e-01*S0+8.471682e+00*S1+(-2.337538e-02)*S2+3.154832e-01*S3+6.546138e-01*S4+2.414722e+01*S5+6.373414e+01*S6+(-2.405200e+03)*S7+4.201108e+01*S8+2.792896e+01*S9 \
V21_part2=V21_part1+3.070367e-01*S10+2.082462e-01*S11+3.752652e-01*S12+4.733818e-01*S13+5.720739e-02*S14+1.132745e-01*S15+7.468935e-01*S16+3.982257e+01*S17+1.505161e+00*S18+1.187522e+00*S19 \
V21_part3=V21_part2+2.024877e-01*S20+6.829275e-01*S21+9.011104e-01*S22+2.079706e+00*S23+2.711643e-01*S24+7.819213e+00*S25+1.448537e+00*S26+5.615862e-01*S27+1.077105e-01*S28+(-2.504431e+00)*S29 \
V21=V21_part3+(-3.631101e+00)*S30+9.322410e-02*S31+1.955827e-01*S32+3.296495e-01*S33+1.567833e+00*S34+2.261335e-01*S35+3.166740e-01*S36 \
V22_part1=1.056220e-01*S0+(-5.999912e-01)*S1+2.428859e+01*S2+1.720943e-01*S3+(-1.571102e-01)*S4+(-3.490036e+01)*S5+(-2.790947e-02)*S6+1.000000e+04*S7+(-4.012677e-01)*S8+(-1.018583e+01)*S9 \
V22_part2=V22_part1+(-7.333863e-01)*S10+(-2.347294e-01)*S11+(-1.193992e-01)*S12+(-2.427500e-01)*S13+1.668950e-01*S14+3.438934e+00*S15+1.598128e-01*S16+3.541002e+00*S17+(-3.924020e-01)*S18+(-5.206302e-01)*S19 \
V22_part3=V22_part2+(-2.742940e-02)*S20+(-4.722902e-02)*S21+(-3.724956e-01)*S22+3.005187e+00*S23+(-7.406536e-02)*S24+(-8.695194e-01)*S25+(-5.942707e-01)*S26+(-9.657643e-02)*S27+(-5.145079e-02)*S28+(-1.261233e-01)*S29 \
V22=V22_part3+3.024986e-01*S30+(-1.882240e+00)*S31+(-3.220154e-02)*S32+1.712208e-01*S33+3.921218e+00*S34+4.759271e-02*S35+3.555914e-03*S36 \
V23_part1=2.270685e-01*S0+(-8.618591e+00)*S1+(-6.897276e+00)*S2+(-1.874723e-01)*S3+7.908639e-03*S4+9.285995e-01*S5+(-5.552773e+01)*S6+(-6.585981e+02)*S7+(-4.128498e+01)*S8+(-1.213009e+01)*S9 \
V23_part2=V23_part1+9.467855e-01*S10+6.152360e-01*S11+4.131010e-02*S12+1.613675e-01*S13+3.943368e-01*S14+(-3.760529e-01)*S15+(-8.235820e-02)*S16+(-3.659931e+01)*S17+(-8.671235e-01)*S18+5.935648e-01*S19 \
V23_part3=V23_part2+2.905502e-01*S20+(-3.868636e-01)*S21+(-4.332675e-01)*S22+(-3.160281e+00)*S23+1.281822e-01*S24+(-6.742800e+00)*S25+(-8.821307e-01)*S26+(-1.954009e-01)*S27+4.256433e-01*S28+9.925283e+00*S29 \
V23=V23_part3+1.225032e+01*S30+3.534723e+00*S31+2.714212e-01*S32+(-5.221038e-01)*S33+(-3.642364e+00)*S34+2.150160e-01*S35+1.451284e-01*S36 \
V24_part1=(-9.490660e+01)*S0+0.000000e+00*S1+0.000000e+00*S2+2.465373e+00*S3+1.951070e+00*S4+1.812007e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V24_part2=V24_part1+0.000000e+00*S10+(-5.291126e+01)*S11+1.388469e+02*S12+(-1.920489e+02)*S13+2.620358e+02*S14+0.000000e+00*S15+4.484921e+01*S16+0.000000e+00*S17+0.000000e+00*S18+(-7.371476e+01)*S19 \
V24_part3=V24_part2+(-2.544525e+01)*S20+(-1.238242e+02)*S21+1.434239e+02*S22+1.007710e+01*S23+0.000000e+00*S24+0.000000e+00*S25+(-6.060881e+02)*S26+0.000000e+00*S27+1.212257e+01*S28+0.000000e+00*S29 \
V24=V24_part3+1.985649e+02*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+1.003806e+03*S36 \
V25_part1=7.854321e+02*S0+0.000000e+00*S1+0.000000e+00*S2+7.765238e+00*S3+2.176925e+00*S4+1.211421e+02*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V25_part2=V25_part1+0.000000e+00*S10+6.313866e+02*S11+4.995269e+02*S12+9.859367e+02*S13+3.557757e+02*S14+0.000000e+00*S15+1.623663e+02*S16+0.000000e+00*S17+0.000000e+00*S18+1.482748e+02*S19 \
V25_part3=V25_part2+8.833340e+01*S20+3.709645e+02*S21+1.449145e+02*S22+2.947820e+01*S23+0.000000e+00*S24+0.000000e+00*S25+1.547768e+03*S26+0.000000e+00*S27+1.504343e+02*S28+0.000000e+00*S29 \
V25=V25_part3+(-8.562169e+01)*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+(-6.115705e+02)*S36 \
V26_part1=2.623170e+01*S0+0.000000e+00*S1+0.000000e+00*S2+3.660103e+02*S3+1.437672e+00*S4+(-1.677367e+00)*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V26_part2=V26_part1+0.000000e+00*S10+1.073380e+02*S11+(-8.297399e+01)*S12+(-1.413169e+01)*S13+(-1.684656e+02)*S14+0.000000e+00*S15+(-2.393781e+01)*S16+0.000000e+00*S17+0.000000e+00*S18+1.960578e+01*S19 \
V26_part3=V26_part2+3.775141e+02*S20+4.456039e+02*S21+3.003157e+02*S22+8.543030e+01*S23+0.000000e+00*S24+0.000000e+00*S25+3.891186e+02*S26+0.000000e+00*S27+6.873966e+01*S28+0.000000e+00*S29 \
V26=V26_part3+(-2.210773e+01)*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+(-3.938299e+02)*S36 \
V27_part1=(-1.348800e+00)*S0+(-6.794009e-01)*S1+1.283603e-01*S2+(-1.376293e+00)*S3+(-7.898844e-01)*S4+(-2.217211e+00)*S5+1.450490e+00*S6+(-2.099578e+01)*S7+1.799126e+00*S8+1.755340e+00*S9 \
V27_part2=V27_part1+(-1.477880e+00)*S10+(-2.927744e+00)*S11+(-4.362218e+00)*S12+(-4.411092e+00)*S13+1.661563e+00*S14+1.358398e-01*S15+(-3.952204e-01)*S16+(-1.894300e+00)*S17+(-1.441525e+00)*S18+(-2.432473e+00)*S19 \
V27_part3=V27_part2+(-2.487202e+00)*S20+(-4.067601e+00)*S21+(-2.734630e+00)*S22+(-1.106972e+00)*S23+(-3.444585e+00)*S24+(-2.445748e+00)*S25+3.429513e+00*S26+(-7.807612e-02)*S27+(-9.679102e-01)*S28+(-4.886981e+00)*S29 \
V27=V27_part3+(-6.983367e+00)*S30+(-2.751444e+00)*S31+(-4.546702e+00)*S32+(-1.890784e-01)*S33+(-8.221871e-01)*S34+(-5.775420e+00)*S35+(-8.454188e+00)*S36 \
V28_part1=8.208389e+00*S0+4.954831e+00*S1+3.261913e+00*S2+2.482535e+00*S3+4.046035e+00*S4+6.889255e+00*S5+(-2.626578e-01)*S6+3.812878e+01*S7+(-2.206883e-01)*S8+3.831126e-01*S9 \
V28_part2=V28_part1+8.590157e+00*S10+8.965724e+00*S11+1.214614e+01*S12+9.207579e+00*S13+3.352810e+00*S14+2.431382e+00*S15+3.024453e+00*S16+4.601927e+00*S17+1.988308e+00*S18+4.958801e+00*S19 \
V28_part3=V28_part2+1.088370e+01*S20+1.123791e+01*S21+6.697657e+00*S22+3.705959e+00*S23+1.003761e+01*S24+1.642358e+01*S25+1.579996e+00*S26+7.975747e+00*S27+8.153180e+00*S28+1.363225e+01*S29 \
V28=V28_part3+1.351968e+01*S30+1.135403e+01*S31+1.215511e+01*S32+4.647235e+00*S33+6.823502e+00*S34+1.442116e+01*S35+1.437677e+01*S36 \
V29_part1=3.803344e+00*S0+3.142188e+00*S1+2.761568e+00*S2+8.606188e+00*S3+4.897572e+00*S4+8.675106e+00*S5+3.224978e+00*S6+3.385138e+01*S7+2.473925e+00*S8+1.909294e+00*S9 \
V29_part2=V29_part1+6.855074e+00*S10+1.037091e+01*S11+1.016544e+01*S12+1.386441e+01*S13+7.339525e+00*S14+3.166997e+00*S15+4.403787e+00*S16+6.551240e+00*S17+1.094238e+01*S18+6.900456e+00*S19 \
V29_part3=V29_part2+1.087047e+01*S20+1.502639e+01*S21+1.663402e+01*S22+6.633628e+00*S23+1.192517e+01*S24+9.378518e+00*S25+5.685302e+00*S26+6.878012e+00*S27+9.999010e+00*S28+1.888699e+01*S29 \
V29=V29_part3+2.467006e+01*S30+1.258495e+01*S31+1.672056e+01*S32+1.481629e+01*S33+1.033587e+01*S34+2.194752e+01*S35+2.936642e+01*S36 \
V30_part1=3.295310e-01*S0+8.216964e-01*S1+2.178590e+00*S2+4.541641e-01*S3+1.756402e-01*S4+2.536899e+03*S5+5.884991e+01*S6+(-2.375140e+03)*S7+4.368056e+01*S8+2.975449e+01*S9 \
V30_part2=V30_part1+2.815077e+00*S10+(-3.393844e-01)*S11+4.110278e+00*S12+(-7.059327e+00)*S13+2.213318e+00*S14+7.804800e-01*S15+3.399089e-02*S16+2.068746e+00*S17+1.257192e+00*S18+1.713662e+00*S19 \
V30_part3=V30_part2+1.543332e+00*S20+5.635855e-01*S21+9.032064e-01*S22+8.259004e-01*S23+(-3.458726e+00)*S24+5.356454e+01*S25+6.618472e-02*S26+1.064092e-01*S27+7.287797e-03*S28+(-2.946750e+00)*S29 \
V30=V30_part3+(-2.610355e+01)*S30+3.064283e-01*S31+1.988872e-02*S32+4.800537e-01*S33+(-6.288333e-02)*S34+(-4.349757e-01)*S35+(-5.859440e-01)*S36 \
V31_part1=1.086010e-01*S0+(-3.057809e-01)*S1+(-2.347825e-01)*S2+1.739102e-02*S3+(-2.576133e-01)*S4+(-2.783027e+02)*S5+(-8.800092e-02)*S6+1.000000e+04*S7+(-5.310722e-01)*S8+(-1.193368e+01)*S9 \
V31_part2=V31_part1+1.338291e+01*S10+(-7.469434e-01)*S11+1.363003e-01*S12+1.426992e-01*S13+(-1.686493e-01)*S14+(-1.860359e-01)*S15+9.929721e-02*S16+(-6.595812e-01)*S17+(-3.038391e-01)*S18+(-1.313970e-01)*S19 \
V31_part3=V31_part2+4.945008e+00*S20+(-1.861495e-01)*S21+(-2.909852e-01)*S22+5.109467e-02*S23+(-2.003011e+00)*S24+(-1.454681e+00)*S25+(-3.916140e-02)*S26+(-1.667875e-01)*S27+4.518589e-01*S28+2.676408e+02*S29 \
V31=V31_part3+6.087180e+01*S30+(-4.190330e-01)*S31+1.514451e+01*S32+1.156906e-01*S33+1.415778e+00*S34+(-7.516631e-01)*S35+(-2.521994e-01)*S36 \
V32_part1=1.990898e-01*S0+1.577529e-01*S1+(-1.108022e+00)*S2+(-1.478959e-01)*S3+8.352192e-01*S4+2.536899e+03*S5+(-4.988054e+01)*S6+(-7.316897e+02)*S7+(-4.308390e+01)*S8+(-1.266772e+01)*S9 \
V32_part2=V32_part1+(-9.001570e+00)*S10+3.901577e+00*S11+(-3.487174e+00)*S12+2.244370e+01*S13+(-1.572574e+00)*S14+(-1.819756e-01)*S15+1.783731e+00*S16+(-1.957009e-01)*S17+(-6.487942e-01)*S18+(-6.457900e-01)*S19 \
V32_part3=V32_part2+(-3.705078e+00)*S20+3.441711e-01*S21+(-4.978716e-01)*S22+3.901354e-01*S23+1.613665e+01*S24+(-5.010935e+01)*S25+1.107680e+00*S26+6.353395e-01*S27+4.672734e-01*S28+(-1.996259e+01)*S29 \
V32=V32_part3+(-1.794818e+01)*S30+7.401353e-01*S31+1.379203e+00*S32+(-8.077692e-01)*S33+1.230285e+00*S34+4.161456e+00*S35+3.765143e+00*S36 \
V33_part1=(-8.677525e+01)*S0+0.000000e+00*S1+1.053797e+02*S2+2.598984e+01*S3+(-3.016068e+01)*S4+(-3.084670e+00)*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V33_part2=V33_part1+0.000000e+00*S10+(-2.072342e+01)*S11+8.481381e+01*S12+(-4.719314e+02)*S13+(-5.316338e+01)*S14+5.620633e+01*S15+4.062637e+01*S16+0.000000e+00*S17+(-2.528685e+01)*S18+2.612739e+01*S19 \
V33_part3=V33_part2+(-9.540693e+00)*S20+(-1.758617e+02)*S21+(-1.061130e+02)*S22+1.111330e+01*S23+(-1.077518e+02)*S24+0.000000e+00*S25+2.900987e+02*S26+6.757793e+01*S27+1.983323e+01*S28+0.000000e+00*S29 \
V33=V33_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+(-1.179869e+01)*S34+3.032729e+02*S35+0.000000e+00*S36 \
V34_part1=7.292206e+02*S0+0.000000e+00*S1+1.290064e+02*S2+1.713298e+02*S3+6.570933e+01*S4+1.015490e+02*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V34_part2=V34_part1+0.000000e+00*S10+5.826061e+02*S11+5.487301e+02*S12+5.497516e+02*S13+1.025642e+02*S14+1.068195e+02*S15+1.523841e+02*S16+0.000000e+00*S17+1.656710e+02*S18+3.800496e+01*S19 \
V34_part3=V34_part2+1.114723e+02*S20+2.792796e+02*S21+5.245184e+02*S22+5.331688e+01*S23+7.764399e+02*S24+0.000000e+00*S25+3.006454e+02*S26+4.679066e+02*S27+8.807846e+01*S28+0.000000e+00*S29 \
V34=V34_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+2.713829e+02*S34+5.731818e+02*S35+0.000000e+00*S36 \
V35_part1=1.729657e+01*S0+0.000000e+00*S1+(-7.677300e+01)*S2+1.781860e+02*S3+(-9.227580e-02)*S4+(-1.832149e+00)*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V35_part2=V35_part1+0.000000e+00*S10+8.246882e+01*S11+(-4.034808e+01)*S12+7.354696e+02*S13+2.388921e+02*S14+(-1.348563e+01)*S15+(-2.725350e+01)*S16+0.000000e+00*S17+3.148873e+02*S18+1.053548e+02*S19 \
V35_part3=V35_part2+3.241336e+02*S20+5.151068e+02*S21+2.692683e+02*S22+6.048035e+01*S23+2.543550e+02*S24+0.000000e+00*S25+(-2.199213e+02)*S26+(-3.909942e+01)*S27+2.738194e+02*S28+0.000000e+00*S29 \
V35=V35_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+1.421961e+02*S34+(-1.276302e+02)*S35+0.000000e+00*S36 \
V36_part1=0.000000e+00*S0+(-1.843471e+00)*S1+(-4.187569e+00)*S2+(-1.912659e+00)*S3+(-5.382352e+00)*S4+0.000000e+00*S5+(-2.610170e+00)*S6+(-3.816326e+00)*S7+(-3.933830e+00)*S8+(-4.847996e+00)*S9 \
V36_part2=V36_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+(-1.718888e+01)*S14+(-2.443883e+00)*S15+(-2.728801e+00)*S16+(-2.619247e+00)*S17+(-2.668495e+00)*S18+(-4.235687e+00)*S19 \
V36_part3=V36_part2+0.000000e+00*S20+0.000000e+00*S21+(-6.094097e+00)*S22+(-1.826792e+00)*S23+0.000000e+00*S24+0.000000e+00*S25+(-1.441278e+01)*S26+(-1.701949e+01)*S27+(-4.064353e+00)*S28+0.000000e+00*S29 \
V36=V36_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+(-1.307794e+01)*S33+(-4.780297e+00)*S34+0.000000e+00*S35+0.000000e+00*S36 \
V37_part1=0.000000e+00*S0+3.527278e+00*S1+8.787077e+00*S2+7.392164e+00*S3+7.677591e+00*S4+0.000000e+00*S5+8.081902e+00*S6+6.396757e+00*S7+8.361358e+00*S8+8.892100e+00*S9 \
V37_part2=V37_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+1.657000e+01*S14+9.048048e+00*S15+7.741874e+00*S16+9.676086e+00*S17+8.935283e+00*S18+8.541199e+00*S19 \
V37_part3=V37_part2+0.000000e+00*S20+0.000000e+00*S21+8.754788e+00*S22+1.061375e+01*S23+0.000000e+00*S24+0.000000e+00*S25+1.449236e+01*S26+1.127465e+01*S27+1.188741e+01*S28+0.000000e+00*S29 \
V37=V37_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+1.664585e+01*S33+1.444816e+01*S34+0.000000e+00*S35+0.000000e+00*S36 \
V38_part1=0.000000e+00*S0+5.044306e+00*S1+4.650708e+00*S2+(-1.339252e+00)*S3+5.089548e+00*S4+0.000000e+00*S5+4.702094e+00*S6+8.199432e+00*S7+5.716939e+00*S8+5.871454e+00*S9 \
V38_part2=V38_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+1.379232e+01*S14+4.181287e+00*S15+5.367813e+00*S16+2.702096e+00*S17+3.423851e-01*S18+6.211660e+00*S19 \
V38_part3=V38_part2+0.000000e+00*S20+0.000000e+00*S21+6.528894e+00*S22+4.366643e+00*S23+0.000000e+00*S24+0.000000e+00*S25+1.895703e+01*S26+1.995251e+01*S27+7.122336e+00*S28+0.000000e+00*S29 \
V38=V38_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+1.222241e+01*S33+1.039142e+01*S34+0.000000e+00*S35+0.000000e+00*S36 \
V39_part1=(-1.079692e+00)*S0+0.000000e+00*S1+0.000000e+00*S2+(-2.207946e-02)*S3+0.000000e+00*S4+0.000000e+00*S5+3.802646e-03*S6+1.801888e-01*S7+(-7.738389e-03)*S8+1.929214e-03*S9 \
V39_part2=V39_part1+0.000000e+00*S10+0.000000e+00*S11+2.566094e-01*S12+5.246572e-02*S13+4.318674e-02*S14+7.542332e-02*S15+0.000000e+00*S16+(-7.084382e-04)*S17+0.000000e+00*S18+(-6.811524e-02)*S19 \
V39_part3=V39_part2+1.880290e-01*S20+(-4.656699e-01)*S21+1.329884e+02*S22+0.000000e+00*S23+2.087767e-01*S24+2.669216e-02*S25+(-6.504589e-01)*S26+(-8.126812e+02)*S27+4.671171e+00*S28+5.623942e-02*S29 \
V39=V39_part3+8.841193e-02*S30+1.055771e-01*S31+3.211340e-01*S32+1.000000e+04*S33+2.200993e-02*S34+1.030417e+00*S35+7.044844e+00*S36 \
V40_part1=5.049284e+01*S0+0.000000e+00*S1+0.000000e+00*S2+(-4.007321e-02)*S3+0.000000e+00*S4+0.000000e+00*S5+(-2.235188e-03)*S6+(-2.210272e-01)*S7+3.054233e-02*S8+1.042740e-03*S9 \
V40_part2=V40_part1+0.000000e+00*S10+0.000000e+00*S11+(-5.434270e-01)*S12+(-9.750840e-02)*S13+(-3.607366e-01)*S14+(-1.556609e-01)*S15+0.000000e+00*S16+(-2.502318e-02)*S17+0.000000e+00*S18+6.237983e-02*S19 \
V40_part3=V40_part2+(-4.561512e-01)*S20+(-1.128738e-01)*S21+2.022729e+01*S22+0.000000e+00*S23+3.739432e-03*S24+(-2.374633e-02)*S25+(-3.275251e-01)*S26+6.881582e+03*S27+3.432909e+02*S28+1.409880e-01*S29 \
V40=V40_part3+6.621809e-02*S30+7.373140e-01*S31+(-1.873766e-02)*S32+1.000000e+04*S33+4.607839e-02*S34+8.711488e-01*S35+6.426146e-01*S36 \
V41_part1=(-5.149193e+00)*S0+0.000000e+00*S1+0.000000e+00*S2+2.110985e-01*S3+0.000000e+00*S4+0.000000e+00*S5+4.313324e-03*S6+3.699712e-02*S7+(-8.143939e-03)*S8+9.470509e-03*S9 \
V41_part2=V41_part1+0.000000e+00*S10+0.000000e+00*S11+7.581803e-01*S12+4.712268e-01*S13+1.017031e+00*S14+1.200870e-01*S15+0.000000e+00*S16+6.829379e-02*S17+0.000000e+00*S18+6.685633e-02*S19 \
V41_part3=V41_part2+8.796091e-01*S20+2.081611e+00*S21+(-2.517405e+02)*S22+0.000000e+00*S23+(-5.368253e-03)*S24+1.254703e-01*S25+3.906469e+00*S26+(-3.822222e+03)*S27+(-1.664547e+02)*S28+(-7.961776e-05)*S29 \
V41=V41_part3+(-1.016127e-05)*S30+(-2.904984e-01)*S31+1.564699e-01*S32+1.000000e+04*S33+3.964014e-01*S34+(-1.754622e+00)*S35+(-1.285994e+01)*S36 \
V42_part1=0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+8.551674e+02*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+(-3.040733e+02)*S7+(-1.112989e+02)*S8+0.000000e+00*S9 \
V42_part2=V42_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+(-3.874375e+02)*S14+1.557944e+03*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V42_part3=V42_part2+0.000000e+00*S20+0.000000e+00*S21+3.105358e+02*S22+0.000000e+00*S23+0.000000e+00*S24+5.124522e+01*S25+0.000000e+00*S26+8.071851e+01*S27+(-3.261219e-01)*S28+0.000000e+00*S29 \
V42=V42_part3+0.000000e+00*S30+0.000000e+00*S31+(-8.509622e+01)*S32+(-3.238860e+02)*S33+2.011420e+02*S34+0.000000e+00*S35+(-3.708997e+02)*S36 \
V43_part1=0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+(-2.583615e+02)*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+1.877766e+03*S7+1.451968e+03*S8+0.000000e+00*S9 \
V43_part2=V43_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+1.160893e+03*S14+(-1.284427e+03)*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V43_part3=V43_part2+0.000000e+00*S20+0.000000e+00*S21+2.927902e+02*S22+0.000000e+00*S23+0.000000e+00*S24+6.043153e+02*S25+0.000000e+00*S26+6.315669e+02*S27+8.687170e-01*S28+0.000000e+00*S29 \
V43=V43_part3+0.000000e+00*S30+0.000000e+00*S31+1.078636e+03*S32+6.299099e+02*S33+(-8.412277e+01)*S34+0.000000e+00*S35+1.564009e+03*S36 \
V44_part1=0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+(-6.303731e+02)*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+4.822655e+01*S7+(-4.271205e+01)*S8+0.000000e+00*S9 \
V44_part2=V44_part1+0.000000e+00*S10+0.000000e+00*S11+0.000000e+00*S12+0.000000e+00*S13+(-8.396261e+01)*S14+(-1.204942e+03)*S15+0.000000e+00*S16+0.000000e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V44_part3=V44_part2+0.000000e+00*S20+0.000000e+00*S21+(-7.568017e+02)*S22+0.000000e+00*S23+0.000000e+00*S24+(-5.600971e+00)*S25+0.000000e+00*S26+3.908375e+01*S27+3.285730e+00*S28+0.000000e+00*S29 \
V44=V44_part3+0.000000e+00*S30+0.000000e+00*S31+2.328074e+02*S32+(-1.579206e+02)*S33+(-1.587955e+02)*S34+0.000000e+00*S35+1.382832e+02*S36 \
V45_part1=1.000000e+04*S0+1.406747e+03*S1+1.000000e+04*S2+(-9.505359e+00)*S3+3.384652e+01*S4+2.177364e+00*S5+1.161904e+01*S6+2.446349e+01*S7+6.684916e+00*S8+7.033781e+00*S9 \
V45_part2=V45_part1+6.566206e-01*S10+(-1.393843e+02)*S11+1.000000e+04*S12+(-3.333031e+03)*S13+8.924976e+03*S14+1.059606e+02*S15+(-3.710481e+00)*S16+(-8.700514e+02)*S17+1.095787e-01*S18+1.123330e+01*S19 \
V45_part3=V45_part2+(-3.332927e+03)*S20+(-1.242490e+01)*S21+(-5.264252e+01)*S22+3.581234e+02*S23+2.130240e+01*S24+6.140243e-01*S25+2.528431e+03*S26+5.601533e+01*S27+(-5.507342e-02)*S28+(-7.910659e+00)*S29 \
V45=V45_part3+(-8.151571e+00)*S30+2.949492e+03*S31+2.861389e-01*S32+2.931772e-02*S33+(-1.776117e+01)*S34+2.458509e-01*S35+3.304323e-01*S36 \
V46_part1=1.000000e+04*S0+4.059910e+02*S1+1.000000e+04*S2+2.697613e-01*S3+(-4.399303e+00)*S4+3.443277e+00*S5+(-1.043618e+01)*S6+(-2.054802e+00)*S7+(-6.381391e+00)*S8+(-5.434046e+00)*S9 \
V46_part2=V46_part1+(-6.383942e+02)*S10+(-2.515180e-01)*S11+1.000000e+04*S12+(-2.253796e-01)*S13+6.904671e+02*S14+2.196329e+01*S15+(-3.202465e+00)*S16+(-3.102552e+01)*S17+(-6.160904e+00)*S18+(-2.054763e+02)*S19 \
V46_part3=V46_part2+(-5.491215e-01)*S20+(-5.284241e-01)*S21+(-1.567319e-01)*S22+1.000000e+04*S23+(-2.402533e+01)*S24+(-7.362269e-01)*S25+1.956327e+01*S26+(-3.538781e-01)*S27+(-6.010036e-01)*S28+(-6.000479e-01)*S29 \
V46=V46_part3+(-4.843548e-01)*S30+1.000000e+04*S31+(-2.247076e-01)*S32+(-8.576527e-02)*S33+(-5.555097e+01)*S34+(-2.500211e-01)*S35+(-1.619931e-01)*S36 \
V47_part1=1.000000e+04*S0+1.000000e+04*S1+1.000000e+04*S2+2.857724e+01*S3+4.754167e+01*S4+8.621690e+00*S5+4.510004e+00*S6+(-5.762572e+00)*S7+2.543647e+00*S8+5.348566e-02*S9 \
V47_part2=V47_part1+7.963071e+02*S10+4.189183e+02*S11+1.000000e+04*S12+1.000000e+04*S13+7.488198e+02*S14+7.074896e+02*S15+1.991031e+01*S16+2.242500e+03*S17+2.105946e+01*S18+1.309545e+03*S19 \
V47_part3=V47_part2+1.000000e+04*S20+3.867216e+01*S21+1.589640e+02*S22+3.213089e+03*S23+(-8.143213e-01)*S24+3.246174e-01*S25+(-3.173953e+03)*S26+(-5.285587e+01)*S27+1.778916e+00*S28+2.526512e+01*S29 \
V47=V47_part3+2.632555e+01*S30+1.000000e+04*S31+(-4.652434e-02)*S32+8.619332e-01*S33+1.243342e+02*S34+1.249003e-01*S35+(-9.761809e-02)*S36 \
V48_part1=0.000000e+00*S0+0.000000e+00*S1+(-1.067619e+00)*S2+1.467007e+00*S3+(-7.987342e-01)*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V48_part2=V48_part1+(-2.506906e+00)*S10+(-1.483037e+00)*S11+0.000000e+00*S12+(-3.908782e+00)*S13+1.345058e+00*S14+(-3.840746e-01)*S15+3.654496e-01*S16+0.000000e+00*S17+(-5.102677e-01)*S18+7.887805e-02*S19 \
V48_part3=V48_part2+(-8.087859e-01)*S20+(-1.770566e+00)*S21+(-5.781052e+00)*S22+9.287514e-02*S23+0.000000e+00*S24+2.095280e-02*S25+0.000000e+00*S26+2.884197e-01*S27+0.000000e+00*S28+0.000000e+00*S29 \
V48=V48_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36 \
V49_part1=0.000000e+00*S0+0.000000e+00*S1+2.160678e+00*S2+(-1.021558e+00)*S3+1.000212e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V49_part2=V49_part1+9.293312e+00*S10+6.282793e+00*S11+0.000000e+00*S12+5.219223e+00*S13+6.201000e-01*S14+9.867818e-01*S15+4.268531e-01*S16+0.000000e+00*S17+5.485679e-01*S18+(-7.122422e-01)*S19 \
V49_part3=V49_part2+9.334145e+00*S20+8.131309e+00*S21+9.790304e+00*S22+7.171382e-01*S23+0.000000e+00*S24+1.617036e+01*S25+0.000000e+00*S26+4.899090e+00*S27+0.000000e+00*S28+0.000000e+00*S29 \
V49=V49_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36 \
V50_part1=0.000000e+00*S0+0.000000e+00*S1+7.879900e-01*S2+2.305071e-01*S3+1.281608e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V50_part2=V50_part1+2.963017e+00*S10+1.456867e+00*S11+0.000000e+00*S12+5.430153e+00*S13+8.738322e-01*S14+7.149754e-01*S15+3.705961e-03*S16+0.000000e+00*S17+1.358817e+00*S18+1.045914e+00*S19 \
V50_part3=V50_part2+3.685256e-01*S20+(-4.811877e-01)*S21+5.357852e+00*S22+8.310210e-01*S23+0.000000e+00*S24+(-3.151428e+00)*S25+0.000000e+00*S26+(-6.519574e-01)*S27+0.000000e+00*S28+0.000000e+00*S29 \
V50=V50_part3+0.000000e+00*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36 \
V51_part1=0.000000e+00*S0+1.521869e-01*S1+5.312893e-01*S2+6.101913e+00*S3+(-4.393149e+00)*S4+1.892049e+01*S5+(-2.306703e+03)*S6+1.000000e+04*S7+(-4.910109e+02)*S8+1.000000e+04*S9 \
V51_part2=V51_part1+1.453578e+00*S10+3.456730e+00*S11+1.000000e+04*S12+5.600292e+01*S13+1.000000e+04*S14+2.591136e+00*S15+(-2.988760e+00)*S16+1.665595e+00*S17+(-1.901391e+00)*S18+1.143263e+01*S19 \
V51_part3=V51_part2+1.000000e+04*S20+(-3.224594e+03)*S21+3.353736e+01*S22+(-1.004048e+00)*S23+(-1.432674e+00)*S24+(-2.872932e+02)*S25+0.000000e+00*S26+1.492068e-01*S27+1.113988e+02*S28+3.797765e+00*S29 \
V51=V51_part3+3.958812e+00*S30+9.830406e-01*S31+2.118726e+01*S32+1.000000e+04*S33+(-1.847833e+01)*S34+7.410173e+03*S35+8.593219e+03*S36 \
V52_part1=0.000000e+00*S0+(-2.169929e-01)*S1+(-4.796114e-01)*S2+4.606591e+00*S3+(-9.994440e-02)*S4+(-7.943725e+00)*S5+1.000000e+04*S6+1.000000e+04*S7+7.790320e+03*S8+1.000000e+04*S9 \
V52_part2=V52_part1+2.953331e-01*S10+4.433973e-02*S11+1.000000e+04*S12+1.133971e+01*S13+1.000000e+04*S14+(-3.835206e+00)*S15+(-2.585200e-01)*S16+(-1.343042e+00)*S17+4.666217e-01*S18+1.705279e+00*S19 \
V52_part3=V52_part2+2.473315e+01*S20+(-2.561590e-01)*S21+(-3.063403e+01)*S22+8.846435e-01*S23+(-4.585450e-01)*S24+1.680291e+03*S25+0.000000e+00*S26+1.993724e-01*S27+(-9.915526e-01)*S28+2.698272e-01*S29 \
V52=V52_part3+5.882317e-01*S30+2.860642e-01*S31+(-9.849851e+00)*S32+1.000000e+04*S33+9.163445e+01*S34+(-1.000000e+04)*S35+(-6.898712e+03)*S36 \
V53_part1=0.000000e+00*S0+1.240299e+00*S1+3.815784e-01*S2+2.325161e+00*S3+1.167450e+01*S4+(-6.597534e+00)*S5+(-9.137123e+02)*S6+9.999738e+03*S7+(-1.762166e+01)*S8+1.000000e+04*S9 \
V53_part2=V53_part1+(-1.562573e+00)*S10+(-3.494355e+00)*S11+1.000000e+04*S12+(-7.796335e+01)*S13+2.419131e+03*S14+(-2.585722e-01)*S15+1.295652e+01*S16+6.166304e-01*S17+8.219221e+00*S18+(-9.864122e+00)*S19 \
V53_part3=V53_part2+1.000000e+04*S20+9.676052e+03*S21+(-1.632726e+00)*S22+5.198010e+00*S23+5.516659e+00*S24+(-1.989800e+02)*S25+0.000000e+00*S26+(-1.739882e-01)*S27+(-2.079388e+02)*S28+(-6.796653e+00)*S29 \
V53=V53_part3+(-7.628539e+00)*S30+(-8.948014e-01)*S31+3.651177e-02*S32+1.867804e+03*S33+(-2.926507e-01)*S34+7.518786e+03*S35+(-1.449067e+03)*S36 \
V54_part1=4.141264e+00*S0+(-1.160762e+00)*S1+8.396574e-01*S2+(-2.149557e+00)*S3+1.714666e+00*S4+0.000000e+00*S5+6.167727e-02*S6+(-6.870121e-03)*S7+2.161311e-01*S8+(-2.359180e-02)*S9 \
V54_part2=V54_part1+5.334491e-01*S10+0.000000e+00*S11+(-4.297675e+00)*S12+0.000000e+00*S13+0.000000e+00*S14+1.267005e-01*S15+0.000000e+00*S16+(-1.028089e+00)*S17+(-2.559903e-01)*S18+(-7.651617e-01)*S19 \
V54_part3=V54_part2+0.000000e+00*S20+(-3.116802e-01)*S21+0.000000e+00*S22+0.000000e+00*S23+(-4.593741e+00)*S24+(-1.545840e+00)*S25+0.000000e+00*S26+0.000000e+00*S27+(-1.234647e+00)*S28+(-1.976535e+01)*S29 \
V54=V54_part3+(-3.640156e+01)*S30+(-3.686577e+00)*S31+0.000000e+00*S32+0.000000e+00*S33+9.641047e-01*S34+0.000000e+00*S35+0.000000e+00*S36 \
V55_part1=1.661025e+01*S0+6.603555e+00*S1+2.107679e+00*S2+3.678628e+00*S3+2.522001e+00*S4+0.000000e+00*S5+2.564157e-01*S6+3.721216e-01*S7+3.448727e-01*S8+6.308800e-01*S9 \
V55_part2=V55_part1+3.833781e+00*S10+0.000000e+00*S11+1.057467e+01*S12+0.000000e+00*S13+0.000000e+00*S14+2.735299e+00*S15+0.000000e+00*S16+3.431840e+00*S17+1.992309e+00*S18+3.142260e+00*S19 \
V55_part3=V55_part2+0.000000e+00*S20+6.938670e+00*S21+0.000000e+00*S22+0.000000e+00*S23+1.682854e+01*S24+3.517551e+00*S25+0.000000e+00*S26+0.000000e+00*S27+5.875751e+00*S28+3.442756e+01*S29 \
V55=V55_part3+3.184724e+01*S30+3.062457e+01*S31+0.000000e+00*S32+0.000000e+00*S33+1.030740e+01*S34+0.000000e+00*S35+0.000000e+00*S36 \
V56_part1=2.461740e+01*S0+(-1.288796e-01)*S1+(-6.054034e-01)*S2+2.001164e+00*S3+(-1.199426e+00)*S4+0.000000e+00*S5+(-2.980854e-03)*S6+(-8.531514e-02)*S7+(-2.236633e-02)*S8+1.398319e-01*S9 \
V56_part2=V56_part1+4.278348e-01*S10+0.000000e+00*S11+3.397689e+00*S12+0.000000e+00*S13+0.000000e+00*S14+6.905742e-01*S15+0.000000e+00*S16+1.679791e+00*S17+3.227647e+00*S18+2.771101e-01*S19 \
V56_part3=V56_part2+0.000000e+00*S20+(-1.249727e+00)*S21+0.000000e+00*S22+0.000000e+00*S23+8.253426e+00*S24+5.849351e+00*S25+0.000000e+00*S26+0.000000e+00*S27+3.078510e-01*S28+3.557055e+01*S29 \
V56=V56_part3+6.440067e+01*S30+3.406640e+00*S31+0.000000e+00*S32+0.000000e+00*S33+1.341180e+00*S34+0.000000e+00*S35+0.000000e+00*S36 \
V57_part1=7.275266e+02*S0+(-5.582366e+00)*S1+(-7.714828e-01)*S2+1.032621e+00*S3+1.220938e+01*S4+6.314584e+01*S5+1.000000e+04*S6+1.000000e+04*S7+(-1.638513e+03)*S8+1.000000e+04*S9 \
V57_part2=V57_part1+4.710287e-01*S10+5.958388e-01*S11+0.000000e+00*S12+1.066292e+00*S13+0.000000e+00*S14+7.445334e+03*S15+4.877325e+00*S16+4.997733e+02*S17+(-4.555214e+00)*S18+(-1.206243e+01)*S19 \
V57_part3=V57_part2+0.000000e+00*S20+3.818473e+02*S21+2.409681e+01*S22+(-4.814090e+00)*S23+5.903564e-02*S24+1.000000e+04*S25+(-2.379716e+02)*S26+9.976804e+03*S27+4.240738e+01*S28+1.213502e+00*S29 \
V57=V57_part3+1.339566e+00*S30+1.000000e+04*S31+0.000000e+00*S32+2.074897e+01*S33+1.659742e+01*S34+0.000000e+00*S35+0.000000e+00*S36 \
V58_part1=1.000000e+04*S0+(-2.709083e+01)*S1+(-2.989876e-01)*S2+1.487632e+02*S3+5.733154e-01*S4+(-7.436069e+01)*S5+(-1.923158e+03)*S6+1.000000e+04*S7+5.421692e+03*S8+1.000000e+04*S9 \
V58_part2=V58_part1+(-7.508700e-01)*S10+(-1.330491e-01)*S11+0.000000e+00*S12+(-2.664474e-01)*S13+0.000000e+00*S14+1.064767e+02*S15+(-4.177073e-01)*S16+4.596390e+01*S17+1.274435e+00*S18+(-2.660973e-01)*S19 \
V58_part3=V58_part2+0.000000e+00*S20+1.000000e+04*S21+2.039873e+00*S22+4.323020e+01*S23+(-2.432020e-02)*S24+1.000000e+04*S25+2.416565e-01*S26+9.977369e+03*S27+(-6.286928e-01)*S28+3.073524e-01*S29 \
V58=V58_part3+3.161779e-01*S30+1.000000e+04*S31+0.000000e+00*S32+(-7.607581e+00)*S33+3.735679e+00*S34+0.000000e+00*S35+0.000000e+00*S36 \
V59_part1=1.000000e+04*S0+1.548039e+02*S1+3.032672e+00*S2+(-1.599593e+02)*S3+(-1.065568e+01)*S4+(-1.295751e+01)*S5+(-2.753583e+03)*S6+1.000000e+04*S7+(-1.207048e+03)*S8+1.000000e+04*S9 \
V59_part2=V59_part1+2.923336e-01*S10+(-1.245831e-01)*S11+0.000000e+00*S12+(-1.041025e+00)*S13+0.000000e+00*S14+1.066170e+03*S15+(-4.010157e+00)*S16+(-5.049957e+02)*S17+1.610786e+01*S18+3.178789e+01*S19 \
V59_part3=V59_part2+0.000000e+00*S20+(-6.641462e+03)*S21+(-9.319773e+00)*S22+(-6.866598e+00)*S23+5.353961e-02*S24+1.000000e+04*S25+7.148264e+02*S26+1.782348e+03*S27+(-7.831359e+01)*S28+(-2.058009e+00)*S29 \
V59=V59_part3+(-2.306160e+00)*S30+(-2.812228e+02)*S31+0.000000e+00*S32+(-2.211372e+01)*S33+(-3.204632e+01)*S34+0.000000e+00*S35+0.000000e+00*S36 \
V60_part1=0.000000e+00*S0+(-9.918220e-01)*S1+0.000000e+00*S2+(-1.905877e+00)*S3+1.979985e+00*S4+0.000000e+00*S5+5.743158e-02*S6+(-6.262406e-03)*S7+2.042847e-01*S8+(-2.646636e-02)*S9 \
V60_part2=V60_part1+5.779478e-01*S10+0.000000e+00*S11+0.000000e+00*S12+(-7.962795e+00)*S13+9.464775e+00*S14+0.000000e+00*S15+0.000000e+00*S16+(-7.881092e-01)*S17+0.000000e+00*S18+(-1.634055e+00)*S19 \
V60_part3=V60_part2+0.000000e+00*S20+(-1.485657e-01)*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+(-5.691775e+00)*S25+1.533285e+00*S26+0.000000e+00*S27+0.000000e+00*S28+(-1.731576e+01)*S29 \
V60=V60_part3+(-2.809552e+01)*S30+(-1.194345e+00)*S31+0.000000e+00*S32+0.000000e+00*S33+(-2.970653e-02)*S34+1.366978e+03*S35+0.000000e+00*S36 \
V61_part1=0.000000e+00*S0+5.465575e+00*S1+0.000000e+00*S2+1.441057e+00*S3+1.590782e+00*S4+0.000000e+00*S5+2.625769e-01*S6+3.708175e-01*S7+3.572914e-01*S8+6.367742e-01*S9 \
V61_part2=V61_part1+3.811427e+00*S10+0.000000e+00*S11+0.000000e+00*S12+1.310909e+01*S13+1.256226e+02*S14+0.000000e+00*S15+0.000000e+00*S16+2.608657e+00*S17+0.000000e+00*S18+3.981672e+00*S19 \
V61_part3=V61_part2+0.000000e+00*S20+7.780548e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+7.447101e+00*S25+(-1.005833e+00)*S26+0.000000e+00*S27+0.000000e+00*S28+4.140480e+01*S29 \
V61=V61_part3+3.931555e+01*S30+1.365442e+01*S31+0.000000e+00*S32+0.000000e+00*S33+4.836030e+00*S34+1.000000e+04*S35+0.000000e+00*S36 \
V62_part1=0.000000e+00*S0+1.214249e-04*S1+0.000000e+00*S2+2.864284e+00*S3+(-1.185691e+00)*S4+0.000000e+00*S5+(-7.569455e-04)*S6+(-8.501353e-02)*S7+(-1.889844e-02)*S8+1.369399e-01*S9 \
V62_part2=V62_part1+3.574333e-01*S10+0.000000e+00*S11+0.000000e+00*S12+9.425203e+00*S13+1.522590e+02*S14+0.000000e+00*S15+0.000000e+00*S16+1.445361e+00*S17+0.000000e+00*S18+(-8.454761e-01)*S19 \
V62_part3=V62_part2+0.000000e+00*S20+(-2.915883e-02)*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+7.802089e+00*S25+(-5.269981e-01)*S26+0.000000e+00*S27+0.000000e+00*S28+2.615834e+01*S29 \
V62=V62_part3+4.145582e+01*S30+3.118931e+00*S31+0.000000e+00*S32+0.000000e+00*S33+1.952456e+00*S34+1.000000e+04*S35+0.000000e+00*S36 \
_P0=V0+V1*radius_+V2*w_ \
_P1=0.5*(_P0+sqrt(_P0*_P0+0.001)) \
_P2=1e-15*_P1 \
_P3=V3+V4*radius_+V5/w_ \
_P4=0.5*(_P3+sqrt(_P3*_P3+0.001)) \
_P5=V6+V7*radius_+V8*w_ \
_P6=0.5*(_P5+sqrt(_P5*_P5+0.001)) \
_P7=1e-09*_P6 \
_P8=1e-09*_P6 \
_P9=V9+V10*radius_+V11/w_ \
_P10=0.5*(_P9+sqrt(_P9*_P9+0.001)) \
_P11=V12+V13*radius_+V14*w_ \
_P12=0.5*(_P11+sqrt(_P11*_P11+0.001)) \
_P13=1e-09*_P12 \
_P14=V15+V16*radius_+V17*w_ \
_P15=0.5*(atan(2*_P14)/1.5708+1) \
_P16=0.7064*_P15 \
_P17=0.7064*_P15 \
_P18=V18+V19*radius_+V20*w_ \
_P19=0.5*(_P18+sqrt(_P18*_P18+0.001)) \
_P20=V21+V22*radius_+V23*w_ \
_P21=0.5*(_P20+sqrt(_P20*_P20+0.001)) \
_P22=V24+V25*radius_+V26*w_ \
_P23=0.5*(_P22+sqrt(_P22*_P22+0.001)) \
_P24=V27+V28*radius_+V29*w_ \
_P25=0.5*(_P24+sqrt(_P24*_P24+0.001)) \
_P26=V30+V31*radius_+V32*w_ \
_P27=0.5*(_P26+sqrt(_P26*_P26+0.001)) \
_P28=V33+V34*radius_+V35*w_ \
_P29=0.5*(_P28+sqrt(_P28*_P28+0.001)) \
_P30=V36+V37*radius_+V38*w_ \
_P31=0.5*(_P30+sqrt(_P30*_P30+0.001)) \
_P32=V39+V40*radius_+V41*w_ \
_P33=0.5*(_P32+sqrt(_P32*_P32+0.001)) \
_P34=V42+V43*radius_+V44*w_ \
_P35=0.5*(_P34+sqrt(_P34*_P34+0.001)) \
_P36=1e-14*_P19 \
_P37=100*_P21 \
_P38=1e-15*_P23 \
_P39=1e-14*_P25 \
_P40=100*_P27 \
_P41=1e-15*_P29 \
_P42=1e-14*_P31 \
_P43=100*_P33 \
_P44=1e-15*_P35 \
_P45=V45+V46*radius_+V47*w_ \
_P46=0.5*(_P45+sqrt(_P45*_P45+0.001)) \
_P47=V48+V49*radius_+V50*w_ \
_P48=0.5*(_P47+sqrt(_P47*_P47+0.001)) \
_P49=100*_P46 \
_P50=1e-13*_P48 \
_P51=V51+V52*radius_+V53*w_ \
_P52=0.5*(_P51+sqrt(_P51*_P51+0.001)) \
_P53=V54+V55*radius_+V56*w_ \
_P54=0.5*(_P53+sqrt(_P53*_P53+0.001)) \
_P55=100*_P52 \
_P56=1e-13*_P54 \
_P57=V57+V58*radius_+V59*w_ \
_P58=0.5*(_P57+sqrt(_P57*_P57+0.001)) \
_P59=V60+V61*radius_+V62*w_ \
_P60=0.5*(_P59+sqrt(_P59*_P59+0.001)) \
_P61=100*_P58 \
_P62=1e-13*_P60
cs (PLUS MINUS) capacitor c=_P2
rs1_1 (PLUS n1_1) resistor r=_P4*(1+drs_diff_ind_rf_pgs_psub_n) tc1=0.003
ls1_1 (n1_1 ni_1) inductor l=_P7*(1+dls_diff_ind_rf_pgs_psub_n)
rs2_1 (ni_1 n2_1) resistor r=_P4*(1+drs_diff_ind_rf_pgs_psub_n) tc1=0.003
ls2_1 (n2_1 MINUS) inductor l=_P8*(1+dls_diff_ind_rf_pgs_psub_n)
rs1_2 (PLUS n1_2) resistor r=_P10*(1+drs_diff_ind_rf_pgs_psub_n) tc1=0.003
ls1_2 (n1_2 MINUS) inductor l=_P13*(1+dls_diff_ind_rf_pgs_psub_n)
k1 mutual_inductor coupling=_P16 ind1=ls1_1 ind2=ls1_2
k2 mutual_inductor coupling=_P17 ind1=ls2_1 ind2=ls1_2
c_1_sub (PLUS _n1_1_sub) capacitor c=_P36
rs_1_sub (_n1_1_sub PSUB) resistor r=_P37
cs_1_sub (_n1_1_sub PSUB) capacitor c=_P38
c_2_sub (MINUS _n1_2_sub) capacitor c=_P39
rs_2_sub (_n1_2_sub PSUB) resistor r=_P40
cs_2_sub (_n1_2_sub PSUB) capacitor c=_P41
c_3_sub (ni_1 _n1_3_sub) capacitor c=_P42
rs_3_sub (_n1_3_sub PSUB) resistor r=_P43
cs_3_sub (_n1_3_sub PSUB) capacitor c=_P44
rx_1_2_sub (_n1_1_sub _n1_2_sub) resistor r=_P49
cx_1_2_sub (_n1_1_sub _n1_2_sub) capacitor c=_P50
rx_1_3_sub (_n1_1_sub _n1_3_sub) resistor r=_P55
cx_1_3_sub (_n1_1_sub _n1_3_sub) capacitor c=_P56
rx_2_3_sub (_n1_2_sub _n1_3_sub) resistor r=_P61
cx_2_3_sub (_n1_2_sub _n1_3_sub) capacitor c=_P62
ends diff_ind_rf_pgs_psub_n
