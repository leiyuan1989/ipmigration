.model nch5 nmos4 l=1 w=1 n=1
.model pch5 pmos4 l=1 w=1 n=1