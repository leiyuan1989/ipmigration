
****
.SUBCKT A2DFFQNX0P5MA10TR  VDD VSS VPW VNW QN   CK A B
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1010 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1016 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1036 QN S VSS VPW NCH W=0.28u L=0.06u
MNA1040 NIN A N1_13 VPW NCH W=0.3u L=0.06u
MNA106 NS S VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_13 B VSS VPW NCH W=0.3u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE020 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE024 NM NCLK NIN VPW NCH W=0.15u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.15u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1012 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1018 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.25u L=0.06u
MPA1038 QN S VDD VNW PCH W=0.37u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1043 NIN A VDD VNW PCH W=0.2u L=0.06u
MPA108 NS S VDD VNW PCH W=0.15u L=0.06u
MPA2 NIN B VDD VNW PCH W=0.2u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN022 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN026 NM BCLK NIN VNW PCH W=0.15u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.15u L=0.06u
.ENDS	A2DFFQNX0P5MA10TR

****
.SUBCKT A2DFFQNX1MA10TR  VDD VSS VPW VNW QN   CK A B
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1024 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.32u L=0.06u
MNA1036 QN S VSS VPW NCH W=0.53u L=0.06u
MNA1040 NIN A N1_13 VPW NCH W=0.45u L=0.06u
MNA108 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_13 B VSS VPW NCH W=0.45u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE012 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE016 NM NCLK NIN VPW NCH W=0.28u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.28u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1022 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1026 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.48u L=0.06u
MPA1038 QN S VDD VNW PCH W=0.7u L=0.06u
MPA104 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1043 NIN A VDD VNW PCH W=0.3u L=0.06u
MPA2 NIN B VDD VNW PCH W=0.3u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN014 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN018 NM BCLK NIN VNW PCH W=0.28u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	A2DFFQNX1MA10TR

****
.SUBCKT A2DFFQNX2MA10TR  VDD VSS VPW VNW QN   CK A B
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1028 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1036 QN S VSS VPW NCH W=1.06u L=0.06u
MNA1040 NIN A N1_13 VPW NCH W=0.58u L=0.06u
MNA108 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_13 B VSS VPW NCH W=0.58u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE012 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE016 NM NCLK NIN VPW NCH W=0.4u L=0.06u
MNOE020 S BCLK M VPW NCH W=0.4u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1026 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1030 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.6u L=0.06u
MPA1038 QN S VDD VNW PCH W=1.4u L=0.06u
MPA104 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1043 NIN A VDD VNW PCH W=0.4u L=0.06u
MPA2 NIN B VDD VNW PCH W=0.4u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN014 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN018 NM BCLK NIN VNW PCH W=0.4u L=0.06u
MPOEN022 S NCLK M VNW PCH W=0.4u L=0.06u
.ENDS	A2DFFQNX2MA10TR

****
.SUBCKT A2DFFQNX3MA10TR  VDD VSS VPW VNW QN   CK A B
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN A N1_13 VPW NCH W=0.58u L=0.06u
MNA1022 QN S VSS VPW NCH W=1.68u L=0.06u
MNA1026 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1030 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1034 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1038 M NM VSS VPW NCH W=0.58u L=0.06u
MNA108 N1_9 NS VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_13 B VSS VPW NCH W=0.58u L=0.06u
MNOE S BCLK M VPW NCH W=0.58u L=0.06u
MNOE012 S NCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE04 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE042 NM NCLK NIN VPW NCH W=0.45u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_11 NS VDD VNW PCH W=0.15u L=0.06u
MPA1019 NIN A VDD VNW PCH W=0.4u L=0.06u
MPA1024 QN S VDD VNW PCH W=2.1u L=0.06u
MPA1028 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1032 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1036 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1040 M NM VDD VNW PCH W=0.7u L=0.06u
MPA2 NIN B VDD VNW PCH W=0.4u L=0.06u
MPOEN S NCLK M VNW PCH W=0.58u L=0.06u
MPOEN014 S BCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN044 NM BCLK NIN VNW PCH W=0.45u L=0.06u
MPOEN06 NM NCLK P1 VNW PCH W=0.15u L=0.06u
.ENDS	A2DFFQNX3MA10TR

****
.SUBCKT A2DFFQX0P5MA10TR  VDD VSS VPW VNW Q   CK A B
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1028 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1036 NIN A N1_13 VPW NCH W=0.4u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1042 Q NS VSS VPW NCH W=0.31u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_13 B VSS VPW NCH W=0.4u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE016 S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE024 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE032 NM NCLK NIN VPW NCH W=0.15u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.25u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1030 M NM VDD VNW PCH W=0.25u L=0.06u
MPA1039 NIN A VDD VNW PCH W=0.2u L=0.06u
MPA1044 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA2 NIN B VDD VNW PCH W=0.2u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN018 S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN026 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN034 NM BCLK NIN VNW PCH W=0.15u L=0.06u
.ENDS	A2DFFQX0P5MA10TR


****
.SUBCKT A2DFFQX1MA10TR  VDD VSS VPW VNW Q   CK A B
MNA1 M NM VSS VPW NCH W=0.28u L=0.06u
MNA1010 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1014 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA102 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA1020 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 NS S VSS VPW NCH W=0.3u L=0.06u
MNA1040 NIN A N1_13 VPW NCH W=0.45u L=0.06u
MNA106 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA2 N1_13 B VSS VPW NCH W=0.45u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE024 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NIN VPW NCH W=0.28u L=0.06u
MNOE032 S BCLK M VPW NCH W=0.28u L=0.06u
MPA1 M NM VDD VNW PCH W=0.4u L=0.06u
MPA1012 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1016 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NS S VDD VNW PCH W=0.47u L=0.06u
MPA104 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA1043 NIN A VDD VNW PCH W=0.3u L=0.06u
MPA108 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA2 NIN B VDD VNW PCH W=0.3u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN026 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NIN VNW PCH W=0.28u L=0.06u
MPOEN034 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	A2DFFQX1MA10TR

****
.SUBCKT A2DFFQX2MA10TR  VDD VSS VPW VNW Q   CK A B
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1028 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1036 NIN A N1_13 VPW NCH W=0.58u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1042 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.43u L=0.06u
MNA2 N1_13 B VSS VPW NCH W=0.58u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE016 S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE024 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE032 NM NCLK NIN VPW NCH W=0.4u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1030 M NM VDD VNW PCH W=0.65u L=0.06u
MPA1039 NIN A VDD VNW PCH W=0.5u L=0.06u
MPA1044 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA2 NIN B VDD VNW PCH W=0.5u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN018 S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN026 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN034 NM BCLK NIN VNW PCH W=0.4u L=0.06u
.ENDS	A2DFFQX2MA10TR

****
.SUBCKT A2DFFQX3MA10TR  VDD VSS VPW VNW Q   CK A B
MNA1 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1010 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA1014 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1020 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 NS S VSS VPW NCH W=0.43u L=0.06u
MNA1040 NIN A N1_13 VPW NCH W=0.58u L=0.06u
MNA106 M NM VSS VPW NCH W=0.51u L=0.06u
MNA2 N1_13 B VSS VPW NCH W=0.58u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE024 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NIN VPW NCH W=0.45u L=0.06u
MNOE032 S BCLK M VPW NCH W=0.45u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1012 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1016 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NS S VDD VNW PCH W=0.7u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA1043 NIN A VDD VNW PCH W=0.5u L=0.06u
MPA108 M NM VDD VNW PCH W=0.77u L=0.06u
MPA2 NIN B VDD VNW PCH W=0.5u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN026 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NIN VNW PCH W=0.45u L=0.06u
MPOEN034 S NCLK M VNW PCH W=0.45u L=0.06u
.ENDS	A2DFFQX3MA10TR

****
.SUBCKT A2DFFQX4MA10TR  VDD VSS VPW VNW Q   CK A B
MNA1 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1010 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA1014 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1020 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 NS S VSS VPW NCH W=0.8u L=0.06u
MNA1040 NIN A N1_13 VPW NCH W=0.58u L=0.06u
MNA106 M NM VSS VPW NCH W=0.58u L=0.06u
MNA2 N1_13 B VSS VPW NCH W=0.58u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE024 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NIN VPW NCH W=0.45u L=0.06u
MNOE032 S BCLK M VPW NCH W=0.58u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1012 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA1016 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NS S VDD VNW PCH W=1u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPA1043 NIN A VDD VNW PCH W=0.5u L=0.06u
MPA108 M NM VDD VNW PCH W=0.7u L=0.06u
MPA2 NIN B VDD VNW PCH W=0.5u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN026 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NIN VNW PCH W=0.45u L=0.06u
MPOEN034 S NCLK M VNW PCH W=0.58u L=0.06u
.ENDS	A2DFFQX4MA10TR

****
.SUBCKT A2SDFFQNX0P5MA10TR  VDD VSS VPW VNW QN   CK A B SE SI
MN0 NMUX A N1 VPW NCH W=0.3u L=0.06u
MN1 N2 NSE VSS VPW NCH W=0.3u L=0.06u
MN2 N1 B N2 VPW NCH W=0.3u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1_15 NS VSS VPW NCH W=0.15u L=0.06u
MNA1021 N1_19 M VSS VPW NCH W=0.15u L=0.06u
MNA1038 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA104 N1_11 SI VSS VPW NCH W=0.15u L=0.06u
MNA1042 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1046 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1050 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1054 QN S VSS VPW NCH W=0.28u L=0.06u
MNOE NMUX SE N1_11 VPW NCH W=0.15u L=0.06u
MNOE016 S NCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE025 NM BCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE030 NM NCLK NMUX VPW NCH W=0.15u L=0.06u
MNOE034 S BCLK M VPW NCH W=0.15u L=0.06u
MP0 NMUX B P1 VNW PCH W=0.29u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.29u L=0.06u
MP2 NMUX A P1 VNW PCH W=0.29u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 P1_17 NS VDD VNW PCH W=0.15u L=0.06u
MPA1023 P1_21 M VDD VNW PCH W=0.15u L=0.06u
MPA1040 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1044 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1048 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1052 M NM VDD VNW PCH W=0.22u L=0.06u
MPA1056 QN S VDD VNW PCH W=0.37u L=0.06u
MPA106 P1_13 SI VDD VNW PCH W=0.15u L=0.06u
MPOEN NMUX NSE P1_13 VNW PCH W=0.15u L=0.06u
MPOEN018 S BCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN027 NM NCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN032 NM BCLK NMUX VNW PCH W=0.15u L=0.06u
MPOEN036 S NCLK M VNW PCH W=0.15u L=0.06u
.ENDS	A2SDFFQNX0P5MA10TR

****
.SUBCKT A2SDFFQNX1MA10TR  VDD VSS VPW VNW QN   CK A B SE SI
MN2 N1 B N2 VPW NCH W=0.5u L=0.06u
MN3 NMUX A N1 VPW NCH W=0.5u L=0.06u
MN4 N2 NSE VSS VPW NCH W=0.5u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_19 M VSS VPW NCH W=0.15u L=0.06u
MNA102 N1_11 SI VSS VPW NCH W=0.15u L=0.06u
MNA1038 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1042 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1046 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1050 M NM VSS VPW NCH W=0.32u L=0.06u
MNA1054 QN S VSS VPW NCH W=0.53u L=0.06u
MNA109 N1_15 NS VSS VPW NCH W=0.15u L=0.06u
MNOE NMUX SE N1_11 VPW NCH W=0.15u L=0.06u
MNOE013 S NCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE022 NM BCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MNOE034 S BCLK M VPW NCH W=0.28u L=0.06u
MP2 NMUX A P1 VNW PCH W=0.48u L=0.06u
MP3 P1 SE VDD VNW PCH W=0.48u L=0.06u
MP4 NMUX B P1 VNW PCH W=0.48u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1011 P1_17 NS VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_21 M VDD VNW PCH W=0.15u L=0.06u
MPA104 P1_13 SI VDD VNW PCH W=0.2u L=0.06u
MPA1040 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1044 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1048 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1052 M NM VDD VNW PCH W=0.48u L=0.06u
MPA1056 QN S VDD VNW PCH W=0.7u L=0.06u
MPOEN NMUX NSE P1_13 VNW PCH W=0.2u L=0.06u
MPOEN015 S BCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN024 NM NCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NMUX VNW PCH W=0.28u L=0.06u
MPOEN036 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	A2SDFFQNX1MA10TR

****
.SUBCKT A2SDFFQNX2MA10TR  VDD VSS VPW VNW QN   CK A B SE SI
MN2 N1 B N2 VPW NCH W=0.61u L=0.06u
MN3 NMUX A N1 VPW NCH W=0.61u L=0.06u
MN4 N2 NSE VSS VPW NCH W=0.61u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_19 M VSS VPW NCH W=0.15u L=0.06u
MNA102 N1_11 SI VSS VPW NCH W=0.15u L=0.06u
MNA1038 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1042 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1046 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1050 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1054 QN S VSS VPW NCH W=1.06u L=0.06u
MNA109 N1_15 NS VSS VPW NCH W=0.15u L=0.06u
MNOE NMUX SE N1_11 VPW NCH W=0.15u L=0.06u
MNOE013 S NCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE022 NM BCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MNOE034 S BCLK M VPW NCH W=0.4u L=0.06u
MP2 NMUX A P1 VNW PCH W=0.59u L=0.06u
MP3 P1 SE VDD VNW PCH W=0.59u L=0.06u
MP4 NMUX B P1 VNW PCH W=0.59u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1011 P1_17 NS VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_21 M VDD VNW PCH W=0.15u L=0.06u
MPA104 P1_13 SI VDD VNW PCH W=0.2u L=0.06u
MPA1040 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1044 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1048 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1052 M NM VDD VNW PCH W=0.56u L=0.06u
MPA1056 QN S VDD VNW PCH W=1.4u L=0.06u
MPOEN NMUX NSE P1_13 VNW PCH W=0.2u L=0.06u
MPOEN015 S BCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN024 NM NCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
MPOEN036 S NCLK M VNW PCH W=0.4u L=0.06u
.ENDS	A2SDFFQNX2MA10TR

****
.SUBCKT A2SDFFQNX3MA10TR  VDD VSS VPW VNW QN   CK A B SE SI
MN5 N1 B N2 VPW NCH W=0.61u L=0.06u
MN6 NMUX A N1 VPW NCH W=0.61u L=0.06u
MN7 N2 NSE VSS VPW NCH W=0.61u L=0.06u
MNA1 N1_11 M VSS VPW NCH W=0.15u L=0.06u
MNA1014 N1_15 NS VSS VPW NCH W=0.15u L=0.06u
MNA1022 QN S VSS VPW NCH W=1.59u L=0.06u
MNA1026 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1030 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA1038 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1042 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1046 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1050 M NM VSS VPW NCH W=0.58u L=0.06u
MNOE S BCLK M VPW NCH W=0.58u L=0.06u
MNOE010 NM BCLK N1_11 VPW NCH W=0.15u L=0.06u
MNOE018 S NCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE034 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE054 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MP5 NMUX A P1 VNW PCH W=0.59u L=0.06u
MP6 P1 SE VDD VNW PCH W=0.59u L=0.06u
MP7 NMUX B P1 VNW PCH W=0.59u L=0.06u
MPA1 P1_13 M VDD VNW PCH W=0.15u L=0.06u
MPA1016 P1_17 NS VDD VNW PCH W=0.15u L=0.06u
MPA1024 QN S VDD VNW PCH W=2.1u L=0.06u
MPA1028 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1032 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1040 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1044 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1048 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1052 M NM VDD VNW PCH W=0.7u L=0.06u
MPOEN S NCLK M VNW PCH W=0.58u L=0.06u
MPOEN012 NM NCLK P1_13 VNW PCH W=0.15u L=0.06u
MPOEN020 S BCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN036 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN056 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
.ENDS	A2SDFFQNX3MA10TR

****
.SUBCKT A2SDFFQX0P5MA10TR  VDD VSS VPW VNW Q   CK A B SE SI
MN0 NMUX A N1 VPW NCH W=0.3u L=0.06u
MN1 N2 NSE VSS VPW NCH W=0.3u L=0.06u
MN2 N1 B N2 VPW NCH W=0.3u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1013 N1_11 NS VSS VPW NCH W=0.15u L=0.06u
MNA1026 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1034 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1038 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1050 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1054 Q NS VSS VPW NCH W=0.31u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE017 S NCLK N1_11 VPW NCH W=0.15u L=0.06u
MNOE030 NM BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE042 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE046 NM NCLK NMUX VPW NCH W=0.15u L=0.06u
MP0 NMUX B P1 VNW PCH W=0.29u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.29u L=0.06u
MP2 NMUX A P1 VNW PCH W=0.29u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.24u L=0.06u
MPA1015 P1_13 NS VDD VNW PCH W=0.15u L=0.06u
MPA1028 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA1036 M NM VDD VNW PCH W=0.22u L=0.06u
MPA1040 P1_21 SI VDD VNW PCH W=0.15u L=0.06u
MPA1052 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1056 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN019 S BCLK P1_13 VNW PCH W=0.15u L=0.06u
MPOEN032 NM NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN044 NMUX NSE P1_21 VNW PCH W=0.15u L=0.06u
MPOEN048 NM BCLK NMUX VNW PCH W=0.15u L=0.06u
.ENDS	A2SDFFQX0P5MA10TR

****
.SUBCKT A2SDFFQX1MA10TR  VDD VSS VPW VNW Q   CK A B SE SI
MN5 N1 B N2 VPW NCH W=0.58u L=0.06u
MN6 NMUX A N1 VPW NCH W=0.58u L=0.06u
MN7 N2 NSE VSS VPW NCH W=0.58u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1010 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1020 N1_11 SI VSS VPW NCH W=0.15u L=0.06u
MNA1026 N1_15 NS VSS VPW NCH W=0.15u L=0.06u
MNA1034 N1_19 M VSS VPW NCH W=0.15u L=0.06u
MNA1050 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1054 NS S VSS VPW NCH W=0.3u L=0.06u
MNA106 M NM VSS VPW NCH W=0.28u L=0.06u
MNOE NMUX SE N1_11 VPW NCH W=0.15u L=0.06u
MNOE030 S NCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE038 NM BCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE042 NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MNOE046 S BCLK M VPW NCH W=0.28u L=0.06u
MP5 NMUX A P1 VNW PCH W=0.5u L=0.06u
MP6 P1 SE VDD VNW PCH W=0.5u L=0.06u
MP7 NMUX B P1 VNW PCH W=0.5u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1012 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA1022 P1_13 SI VDD VNW PCH W=0.2u L=0.06u
MPA1028 P1_17 NS VDD VNW PCH W=0.15u L=0.06u
MPA1036 P1_21 M VDD VNW PCH W=0.15u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1052 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1056 NS S VDD VNW PCH W=0.47u L=0.06u
MPA108 M NM VDD VNW PCH W=0.4u L=0.06u
MPOEN NMUX NSE P1_13 VNW PCH W=0.2u L=0.06u
MPOEN032 S BCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN040 NM NCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN044 NM BCLK NMUX VNW PCH W=0.28u L=0.06u
MPOEN048 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	A2SDFFQX1MA10TR

****
.SUBCKT A2SDFFQX2MA10TR  VDD VSS VPW VNW Q   CK A B SE SI
MN2 N1 B N2 VPW NCH W=0.62u L=0.06u
MN3 NMUX A N1 VPW NCH W=0.62u L=0.06u
MN4 N2 NSE VSS VPW NCH W=0.62u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1012 N1_11 NS VSS VPW NCH W=0.15u L=0.06u
MNA1026 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1034 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1038 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1050 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1054 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.44u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE016 S NCLK N1_11 VPW NCH W=0.15u L=0.06u
MNOE030 NM BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE042 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE046 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MP2 NMUX A P1 VNW PCH W=0.58u L=0.06u
MP3 P1 SE VDD VNW PCH W=0.58u L=0.06u
MP4 NMUX B P1 VNW PCH W=0.58u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1014 P1_13 NS VDD VNW PCH W=0.15u L=0.06u
MPA1028 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA1036 M NM VDD VNW PCH W=0.57u L=0.06u
MPA1040 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1052 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1056 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN018 S BCLK P1_13 VNW PCH W=0.15u L=0.06u
MPOEN032 NM NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN044 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN048 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
.ENDS	A2SDFFQX2MA10TR

****
.SUBCKT A2SDFFQX3MA10TR  VDD VSS VPW VNW Q   CK A B SE SI
MN5 N1 B N2 VPW NCH W=0.62u L=0.06u
MN6 NMUX A N1 VPW NCH W=0.62u L=0.06u
MN7 N2 NSE VSS VPW NCH W=0.62u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1010 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1020 N1_11 NS VSS VPW NCH W=0.15u L=0.06u
MNA1026 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1042 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1046 NS S VSS VPW NCH W=0.47u L=0.06u
MNA1050 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA106 M NM VSS VPW NCH W=0.51u L=0.06u
MNOE S NCLK N1_11 VPW NCH W=0.15u L=0.06u
MNOE030 NM BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE034 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE038 S BCLK M VPW NCH W=0.45u L=0.06u
MNOE054 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MP5 NMUX A P1 VNW PCH W=0.58u L=0.06u
MP6 P1 SE VDD VNW PCH W=0.58u L=0.06u
MP7 NMUX B P1 VNW PCH W=0.58u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1012 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1022 P1_13 NS VDD VNW PCH W=0.15u L=0.06u
MPA1028 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA1044 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1048 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1052 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA108 M NM VDD VNW PCH W=0.77u L=0.06u
MPOEN S BCLK P1_13 VNW PCH W=0.15u L=0.06u
MPOEN032 NM NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN036 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN040 S NCLK M VNW PCH W=0.45u L=0.06u
MPOEN056 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
.ENDS	A2SDFFQX3MA10TR

****
.SUBCKT A2SDFFQX4MA10TR  VDD VSS VPW VNW Q   CK A B SE SI
MN5 N1 B N2 VPW NCH W=0.62u L=0.06u
MN6 NMUX A N1 VPW NCH W=0.62u L=0.06u
MN7 N2 NSE VSS VPW NCH W=0.62u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1010 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1020 N1_11 NS VSS VPW NCH W=0.15u L=0.06u
MNA1026 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1042 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1046 NS S VSS VPW NCH W=0.8u L=0.06u
MNA1050 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA106 M NM VSS VPW NCH W=0.58u L=0.06u
MNOE S NCLK N1_11 VPW NCH W=0.15u L=0.06u
MNOE030 NM BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE034 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE038 S BCLK M VPW NCH W=0.58u L=0.06u
MNOE054 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MP5 NMUX A P1 VNW PCH W=0.58u L=0.06u
MP6 P1 SE VDD VNW PCH W=0.58u L=0.06u
MP7 NMUX B P1 VNW PCH W=0.58u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1012 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA1022 P1_13 NS VDD VNW PCH W=0.15u L=0.06u
MPA1028 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPA1044 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1048 NS S VDD VNW PCH W=1u L=0.06u
MPA1052 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA108 M NM VDD VNW PCH W=0.7u L=0.06u
MPOEN S BCLK P1_13 VNW PCH W=0.15u L=0.06u
MPOEN032 NM NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN036 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN040 S NCLK M VNW PCH W=0.58u L=0.06u
MPOEN056 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
.ENDS	A2SDFFQX4MA10TR

****
.SUBCKT ADDFX1MA10TR  VDD VSS VPW VNW CO S   A B CI
MN0 NCOUT CI N1 VPW NCH W=0.39u L=0.06u
MN1 N1 A VSS VPW NCH W=0.39u L=0.06u
MN10 NET49 A NET46 VPW NCH W=0.35u L=0.06u
MN11 NET46 B VSS VPW NCH W=0.35u L=0.06u
MN2 N1 B VSS VPW NCH W=0.39u L=0.06u
MN3 NET34 B VSS VPW NCH W=0.39u L=0.06u
MN4 NCOUT A NET34 VPW NCH W=0.39u L=0.06u
MN5 N2 A VSS VPW NCH W=0.35u L=0.06u
MN6 N2 CI VSS VPW NCH W=0.35u L=0.06u
MN7 NSUM NCOUT N2 VPW NCH W=0.35u L=0.06u
MN8 N2 B VSS VPW NCH W=0.35u L=0.06u
MN9 NSUM CI NET49 VPW NCH W=0.35u L=0.06u
MNA1 CO NCOUT VSS VPW NCH W=0.53u L=0.06u
MNA1022 S NSUM VSS VPW NCH W=0.53u L=0.06u
MP0 NCOUT CI P1 VNW PCH W=0.65u L=0.06u
MP1 P1 A VDD VNW PCH W=0.65u L=0.06u
MP10 NET87 A NET84 VNW PCH W=0.45u L=0.06u
MP11 NET84 B VDD VNW PCH W=0.45u L=0.06u
MP2 P1 B VDD VNW PCH W=0.65u L=0.06u
MP3 NCOUT A NET69 VNW PCH W=0.65u L=0.06u
MP4 NET69 B VDD VNW PCH W=0.65u L=0.06u
MP5 P2 A VDD VNW PCH W=0.45u L=0.06u
MP6 P2 CI VDD VNW PCH W=0.45u L=0.06u
MP7 NSUM NCOUT P2 VNW PCH W=0.45u L=0.06u
MP8 P2 B VDD VNW PCH W=0.45u L=0.06u
MP9 NSUM CI NET87 VNW PCH W=0.45u L=0.06u
MPA1 CO NCOUT VDD VNW PCH W=0.7u L=0.06u
MPA1024 S NSUM VDD VNW PCH W=0.7u L=0.06u
.ENDS	ADDFX1MA10TR

****
.SUBCKT ADDFX1P4MA10TR  VDD VSS VPW VNW CO S   A B CI
MN0 NCOUT CI N1 VPW NCH W=0.39u L=0.06u
MN1 N1 A VSS VPW NCH W=0.39u L=0.06u
MN10 NET111 A NET105 VPW NCH W=0.35u L=0.06u
MN11 NET105 B VSS VPW NCH W=0.35u L=0.06u
MN2 N1 B VSS VPW NCH W=0.39u L=0.06u
MN3 NET87 B VSS VPW NCH W=0.39u L=0.06u
MN4 NCOUT A NET87 VPW NCH W=0.39u L=0.06u
MN5 N2 A VSS VPW NCH W=0.35u L=0.06u
MN6 N2 CI VSS VPW NCH W=0.35u L=0.06u
MN7 NSUM NCOUT N2 VPW NCH W=0.35u L=0.06u
MN8 N2 B VSS VPW NCH W=0.35u L=0.06u
MN9 NSUM CI NET111 VPW NCH W=0.35u L=0.06u
MNA1 CO NCOUT VSS VPW NCH W=0.74u L=0.06u
MNA1022 S NSUM VSS VPW NCH W=0.74u L=0.06u
MP0 NCOUT CI P1 VNW PCH W=0.65u L=0.06u
MP1 P1 A VDD VNW PCH W=0.65u L=0.06u
MP10 NET68 A NET71 VNW PCH W=0.45u L=0.06u
MP11 NET71 B VDD VNW PCH W=0.45u L=0.06u
MP2 P1 B VDD VNW PCH W=0.65u L=0.06u
MP3 NCOUT A NET50 VNW PCH W=0.65u L=0.06u
MP4 NET50 B VDD VNW PCH W=0.65u L=0.06u
MP5 P2 A VDD VNW PCH W=0.45u L=0.06u
MP6 P2 CI VDD VNW PCH W=0.45u L=0.06u
MP7 NSUM NCOUT P2 VNW PCH W=0.45u L=0.06u
MP8 P2 B VDD VNW PCH W=0.45u L=0.06u
MP9 NSUM CI NET68 VNW PCH W=0.45u L=0.06u
MPA1 CO NCOUT VDD VNW PCH W=0.98u L=0.06u
MPA1024 S NSUM VDD VNW PCH W=0.98u L=0.06u
.ENDS	ADDFX1P4MA10TR

****
.SUBCKT ADDFX2MA10TR  VDD VSS VPW VNW CO S   A B CI
MN0 NCOUT CI N1 VPW NCH W=0.39u L=0.06u
MN1 N1 A VSS VPW NCH W=0.39u L=0.06u
MN10 NET111 A NET105 VPW NCH W=0.35u L=0.06u
MN11 NET105 B VSS VPW NCH W=0.35u L=0.06u
MN2 N1 B VSS VPW NCH W=0.39u L=0.06u
MN3 NET87 B VSS VPW NCH W=0.39u L=0.06u
MN4 NCOUT A NET87 VPW NCH W=0.39u L=0.06u
MN5 N2 A VSS VPW NCH W=0.35u L=0.06u
MN6 N2 CI VSS VPW NCH W=0.35u L=0.06u
MN7 NSUM NCOUT N2 VPW NCH W=0.35u L=0.06u
MN8 N2 B VSS VPW NCH W=0.35u L=0.06u
MN9 NSUM CI NET111 VPW NCH W=0.35u L=0.06u
MNA1 CO NCOUT VSS VPW NCH W=1.06u L=0.06u
MNA1022 S NSUM VSS VPW NCH W=1.06u L=0.06u
MP0 NCOUT CI P1 VNW PCH W=0.65u L=0.06u
MP1 P1 A VDD VNW PCH W=0.65u L=0.06u
MP10 NET68 A NET71 VNW PCH W=0.45u L=0.06u
MP11 NET71 B VDD VNW PCH W=0.45u L=0.06u
MP2 P1 B VDD VNW PCH W=0.65u L=0.06u
MP3 NCOUT A NET50 VNW PCH W=0.65u L=0.06u
MP4 NET50 B VDD VNW PCH W=0.65u L=0.06u
MP5 P2 A VDD VNW PCH W=0.45u L=0.06u
MP6 P2 CI VDD VNW PCH W=0.45u L=0.06u
MP7 NSUM NCOUT P2 VNW PCH W=0.45u L=0.06u
MP8 P2 B VDD VNW PCH W=0.45u L=0.06u
MP9 NSUM CI NET68 VNW PCH W=0.45u L=0.06u
MPA1 CO NCOUT VDD VNW PCH W=1.4u L=0.06u
MPA1024 S NSUM VDD VNW PCH W=1.4u L=0.06u
.ENDS	ADDFX2MA10TR

****
.SUBCKT ADDHX1MA10TR  VDD VSS VPW VNW CO S   A B
MNA1 NSUM NCOUT N1 VPW NCH W=0.4u L=0.06u
MNA1010 NCOUT A N1_4 VPW NCH W=0.42u L=0.06u
MNA1016 CO NCOUT VSS VPW NCH W=0.53u L=0.06u
MNA106 S NSUM VSS VPW NCH W=0.53u L=0.06u
MNA2 N1_4 B VSS VPW NCH W=0.42u L=0.06u
MNB1 N1 A VSS VPW NCH W=0.4u L=0.06u
MNB2 N1 B VSS VPW NCH W=0.4u L=0.06u
MPA1 NSUM NCOUT VDD VNW PCH W=0.29u L=0.06u
MPA1013 NCOUT A VDD VNW PCH W=0.46u L=0.06u
MPA1018 CO NCOUT VDD VNW PCH W=0.7u L=0.06u
MPA108 S NSUM VDD VNW PCH W=0.7u L=0.06u
MPA2 NCOUT B VDD VNW PCH W=0.46u L=0.06u
MPB1 NSUM A P1 VNW PCH W=0.4u L=0.06u
MPB2 P1 B VDD VNW PCH W=0.4u L=0.06u
.ENDS	ADDHX1MA10TR

****
.SUBCKT ADDHX1P4MA10TR  VDD VSS VPW VNW CO S   A B
MNA1 NSUM NCOUT N1 VPW NCH W=0.58u L=0.06u
MNA1010 NCOUT A N1_4 VPW NCH W=0.58u L=0.06u
MNA1016 CO NCOUT VSS VPW NCH W=0.74u L=0.06u
MNA106 S NSUM VSS VPW NCH W=0.74u L=0.06u
MNA2 N1_4 B VSS VPW NCH W=0.58u L=0.06u
MNB1 N1 A VSS VPW NCH W=0.58u L=0.06u
MNB2 N1 B VSS VPW NCH W=0.58u L=0.06u
MPA1 NSUM NCOUT VDD VNW PCH W=0.42u L=0.06u
MPA1013 NCOUT A VDD VNW PCH W=0.64u L=0.06u
MPA1018 CO NCOUT VDD VNW PCH W=0.98u L=0.06u
MPA108 S NSUM VDD VNW PCH W=0.98u L=0.06u
MPA2 NCOUT B VDD VNW PCH W=0.64u L=0.06u
MPB1 NSUM A P1 VNW PCH W=0.58u L=0.06u
MPB2 P1 B VDD VNW PCH W=0.58u L=0.06u
.ENDS	ADDHX1P4MA10TR

****
.SUBCKT ADDHX2MA10TR  VDD VSS VPW VNW CO S   A B
MNA1 NSUM NCOUT N1 VPW NCH W=0.58u L=0.06u
MNA1010 NCOUT A N1_4 VPW NCH W=0.58u L=0.06u
MNA1016 CO NCOUT VSS VPW NCH W=1.06u L=0.06u
MNA106 S NSUM VSS VPW NCH W=1.06u L=0.06u
MNA2 N1_4 B VSS VPW NCH W=0.58u L=0.06u
MNB1 N1 A VSS VPW NCH W=0.58u L=0.06u
MNB2 N1 B VSS VPW NCH W=0.58u L=0.06u
MPA1 NSUM NCOUT VDD VNW PCH W=0.42u L=0.06u
MPA1013 NCOUT A VDD VNW PCH W=0.64u L=0.06u
MPA1018 CO NCOUT VDD VNW PCH W=1.4u L=0.06u
MPA108 S NSUM VDD VNW PCH W=1.4u L=0.06u
MPA2 NCOUT B VDD VNW PCH W=0.64u L=0.06u
MPB1 NSUM A P1 VNW PCH W=0.58u L=0.06u
MPB2 P1 B VDD VNW PCH W=0.58u L=0.06u
.ENDS	ADDHX2MA10TR

****
.SUBCKT AND2X0P5MA10TR  VDD VSS VPW VNW Y   A B
MNA1 INT A N1 VPW NCH W=0.19u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.19u L=0.06u
MPA1 INT A VDD VNW PCH W=0.155u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA2 INT B VDD VNW PCH W=0.155u L=0.06u
.ENDS	AND2X0P5MA10TR

****
.SUBCKT AND2X0P7MA10TR  VDD VSS VPW VNW Y   A B
MNA1 INT A N1 VPW NCH W=0.235u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.37u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.235u L=0.06u
MPA1 INT A VDD VNW PCH W=0.195u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA2 INT B VDD VNW PCH W=0.195u L=0.06u
.ENDS	AND2X0P7MA10TR

****

****
.SUBCKT AND2X1MA10TR  VDD VSS VPW VNW Y   A B
MNA1 INT A N1 VPW NCH W=0.305u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.305u L=0.06u
MPA1 INT A VDD VNW PCH W=0.25u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA2 INT B VDD VNW PCH W=0.25u L=0.06u
.ENDS	AND2X1MA10TR

****
.SUBCKT AND2X1P4MA10TR  VDD VSS VPW VNW Y   A B
MNA1 INT A N1 VPW NCH W=0.44u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.74u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.44u L=0.06u
MPA1 INT A VDD VNW PCH W=0.36u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.98u L=0.06u
MPA2 INT B VDD VNW PCH W=0.36u L=0.06u
.ENDS	AND2X1P4MA10TR

****
.SUBCKT AND2X2MA10TR  VDD VSS VPW VNW Y   A B
MNA1 INT A N1 VPW NCH W=0.58u L=0.06u
MNA104 Y INT VSS VPW NCH W=1.06u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.58u L=0.06u
MPA1 INT A VDD VNW PCH W=0.475u L=0.06u
MPA106 Y INT VDD VNW PCH W=1.4u L=0.06u
MPA2 INT B VDD VNW PCH W=0.475u L=0.06u
.ENDS	AND2X2MA10TR

****

****

****

****

****
.SUBCKT AND3X0P5MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA102 INT A N2 VPW NCH W=0.335u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.335u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.335u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA105 INT A VDD VNW PCH W=0.205u L=0.06u
MPA2 INT B VDD VNW PCH W=0.205u L=0.06u
MPA3 INT C VDD VNW PCH W=0.205u L=0.06u
.ENDS	AND3X0P5MA10TR

****
.SUBCKT AND3X0P7MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MNA102 INT A N2 VPW NCH W=0.4u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.4u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.4u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA105 INT A VDD VNW PCH W=0.245u L=0.06u
MPA2 INT B VDD VNW PCH W=0.245u L=0.06u
MPA3 INT C VDD VNW PCH W=0.245u L=0.06u
.ENDS	AND3X0P7MA10TR

****
.SUBCKT AND3X11MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=5.83u L=0.06u
MNA102 INT A N2 VPW NCH W=4.94u L=0.06u
MNA2 N2 B N1 VPW NCH W=4.94u L=0.06u
MNA3 N1 C VSS VPW NCH W=4.94u L=0.06u
MPA1 Y INT VDD VNW PCH W=7.7u L=0.06u
MPA105 INT A VDD VNW PCH W=3.03u L=0.06u
MPA2 INT B VDD VNW PCH W=3.03u L=0.06u
MPA3 INT C VDD VNW PCH W=3.03u L=0.06u
.ENDS	AND3X11MA10TR

****
.SUBCKT AND3X1MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MNA102 INT A N2 VPW NCH W=0.505u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.505u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.505u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA105 INT A VDD VNW PCH W=0.31u L=0.06u
MPA2 INT B VDD VNW PCH W=0.31u L=0.06u
MPA3 INT C VDD VNW PCH W=0.31u L=0.06u
.ENDS	AND3X1MA10TR

****
.SUBCKT AND3X1P4MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=0.74u L=0.06u
MNA102 INT A N2 VPW NCH W=0.695u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.695u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.695u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.98u L=0.06u
MPA105 INT A VDD VNW PCH W=0.425u L=0.06u
MPA2 INT B VDD VNW PCH W=0.425u L=0.06u
MPA3 INT C VDD VNW PCH W=0.425u L=0.06u
.ENDS	AND3X1P4MA10TR

****

****

****
.SUBCKT AND3X4MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=2.12u L=0.06u
MNA102 INT A N2 VPW NCH W=1.74u L=0.06u
MNA2 N2 B N1 VPW NCH W=1.74u L=0.06u
MNA3 N1 C VSS VPW NCH W=1.74u L=0.06u
MPA1 Y INT VDD VNW PCH W=2.8u L=0.06u
MPA105 INT A VDD VNW PCH W=1.08u L=0.06u
MPA2 INT B VDD VNW PCH W=1.08u L=0.06u
MPA3 INT C VDD VNW PCH W=1.08u L=0.06u
.ENDS	AND3X4MA10TR

****
.SUBCKT AND3X6MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=3.18u L=0.06u
MNA102 INT A N2 VPW NCH W=2.64u L=0.06u
MNA2 N2 B N1 VPW NCH W=2.64u L=0.06u
MNA3 N1 C VSS VPW NCH W=2.64u L=0.06u
MPA1 Y INT VDD VNW PCH W=4.2u L=0.06u
MPA105 INT A VDD VNW PCH W=1.62u L=0.06u
MPA2 INT B VDD VNW PCH W=1.62u L=0.06u
MPA3 INT C VDD VNW PCH W=1.62u L=0.06u
.ENDS	AND3X6MA10TR

****
.SUBCKT AND3X8MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=4.24u L=0.06u
MNA102 INT A N2 VPW NCH W=3.48u L=0.06u
MNA2 N2 B N1 VPW NCH W=3.48u L=0.06u
MNA3 N1 C VSS VPW NCH W=3.48u L=0.06u
MPA1 Y INT VDD VNW PCH W=5.6u L=0.06u
MPA105 INT A VDD VNW PCH W=2.135u L=0.06u
MPA2 INT B VDD VNW PCH W=2.135u L=0.06u
MPA3 INT C VDD VNW PCH W=2.135u L=0.06u
.ENDS	AND3X8MA10TR

****
.SUBCKT AND4X0P5MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA102 INT A N3 VPW NCH W=0.485u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.485u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.485u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.485u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA105 INT A VDD VNW PCH W=0.245u L=0.06u
MPA2 INT B VDD VNW PCH W=0.245u L=0.06u
MPA3 INT C VDD VNW PCH W=0.245u L=0.06u
MPA4 INT D VDD VNW PCH W=0.245u L=0.06u
.ENDS	AND4X0P5MA10TR

****
.SUBCKT AND4X0P7MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MNA102 INT A N3 VPW NCH W=0.575u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.575u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.575u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.575u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA105 INT A VDD VNW PCH W=0.29u L=0.06u
MPA2 INT B VDD VNW PCH W=0.29u L=0.06u
MPA3 INT C VDD VNW PCH W=0.29u L=0.06u
MPA4 INT D VDD VNW PCH W=0.29u L=0.06u
.ENDS	AND4X0P7MA10TR

****
.SUBCKT AND4X1MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MNA102 INT A N3 VPW NCH W=0.72u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.72u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.72u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.72u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA105 INT A VDD VNW PCH W=0.365u L=0.06u
MPA2 INT B VDD VNW PCH W=0.365u L=0.06u
MPA3 INT C VDD VNW PCH W=0.365u L=0.06u
MPA4 INT D VDD VNW PCH W=0.365u L=0.06u
.ENDS	AND4X1MA10TR

****

****
.SUBCKT AND4X2MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y INT VSS VPW NCH W=1.06u L=0.06u
MNA102 INT A N3 VPW NCH W=1.35u L=0.06u
MNA2 N3 B N2 VPW NCH W=1.35u L=0.06u
MNA3 N2 C N1 VPW NCH W=1.35u L=0.06u
MNA4 N1 D VSS VPW NCH W=1.35u L=0.06u
MPA1 Y INT VDD VNW PCH W=1.4u L=0.06u
MPA105 INT A VDD VNW PCH W=0.685u L=0.06u
MPA2 INT B VDD VNW PCH W=0.685u L=0.06u
MPA3 INT C VDD VNW PCH W=0.685u L=0.06u
MPA4 INT D VDD VNW PCH W=0.685u L=0.06u
.ENDS	AND4X2MA10TR

****
.SUBCKT AND4X3MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y INT VSS VPW NCH W=1.59u L=0.06u
MNA102 INT A N3 VPW NCH W=1.915u L=0.06u
MNA2 N3 B N2 VPW NCH W=1.915u L=0.06u
MNA3 N2 C N1 VPW NCH W=1.915u L=0.06u
MNA4 N1 D VSS VPW NCH W=1.915u L=0.06u
MPA1 Y INT VDD VNW PCH W=2.1u L=0.06u
MPA105 INT A VDD VNW PCH W=0.97u L=0.06u
MPA2 INT B VDD VNW PCH W=0.97u L=0.06u
MPA3 INT C VDD VNW PCH W=0.97u L=0.06u
MPA4 INT D VDD VNW PCH W=0.97u L=0.06u
.ENDS	AND4X3MA10TR

****
.SUBCKT AND4X4MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y INT VSS VPW NCH W=2.12u L=0.06u
MNA102 INT A N3 VPW NCH W=2.545u L=0.06u
MNA2 N3 B N2 VPW NCH W=2.545u L=0.06u
MNA3 N2 C N1 VPW NCH W=2.545u L=0.06u
MNA4 N1 D VSS VPW NCH W=2.545u L=0.06u
MPA1 Y INT VDD VNW PCH W=2.8u L=0.06u
MPA105 INT A VDD VNW PCH W=1.29u L=0.06u
MPA2 INT B VDD VNW PCH W=1.29u L=0.06u
MPA3 INT C VDD VNW PCH W=1.29u L=0.06u
MPA4 INT D VDD VNW PCH W=1.29u L=0.06u
.ENDS	AND4X4MA10TR

****
.SUBCKT AND4X6MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y INT VSS VPW NCH W=3.18u L=0.06u
MNA102 INT A N3 VPW NCH W=3.74u L=0.06u
MNA2 N3 B N2 VPW NCH W=3.74u L=0.06u
MNA3 N2 C N1 VPW NCH W=3.74u L=0.06u
MNA4 N1 D VSS VPW NCH W=3.74u L=0.06u
MPA1 Y INT VDD VNW PCH W=4.2u L=0.06u
MPA105 INT A VDD VNW PCH W=1.9u L=0.06u
MPA2 INT B VDD VNW PCH W=1.9u L=0.06u
MPA3 INT C VDD VNW PCH W=1.9u L=0.06u
MPA4 INT D VDD VNW PCH W=1.9u L=0.06u
.ENDS	AND4X6MA10TR

****
.SUBCKT AND4X8MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y INT VSS VPW NCH W=4.24u L=0.06u
MNA102 INT A N3 VPW NCH W=5.09u L=0.06u
MNA2 N3 B N2 VPW NCH W=5.09u L=0.06u
MNA3 N2 C N1 VPW NCH W=5.09u L=0.06u
MNA4 N1 D VSS VPW NCH W=5.09u L=0.06u
MPA1 Y INT VDD VNW PCH W=5.6u L=0.06u
MPA105 INT A VDD VNW PCH W=2.58u L=0.06u
MPA2 INT B VDD VNW PCH W=2.58u L=0.06u
MPA3 INT C VDD VNW PCH W=2.58u L=0.06u
MPA4 INT D VDD VNW PCH W=2.58u L=0.06u
.ENDS	AND4X8MA10TR

****
.SUBCKT ANTENNA2A10TR  VDD VSS VPW VNW A
DD0 VPW A NDIO AREA=6E-08u PJ=1u
.ENDS	ANTENNA2A10TR

****
.SUBCKT AO1B2X0P5MA10TR  VDD VSS VPW VNW Y   A0N B0 B1
MNA1 INT B0 N1 VPW NCH W=0.15u L=0.06u
MNA104 Y INT N1_2 VPW NCH W=0.29u L=0.06u
MNA2 N1 B1 VSS VPW NCH W=0.15u L=0.06u
MNA206 N1_2 A0N VSS VPW NCH W=0.29u L=0.06u
MPA1 INT B0 VDD VNW PCH W=0.185u L=0.06u
MPA108 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA2 INT B1 VDD VNW PCH W=0.185u L=0.06u
MPA2010 Y A0N VDD VNW PCH W=0.35u L=0.06u
.ENDS	AO1B2X0P5MA10TR

****
.SUBCKT AO1B2X0P7MA10TR  VDD VSS VPW VNW Y   A0N B0 B1
MNA1 INT B0 N1 VPW NCH W=0.18u L=0.06u
MNA104 Y INT N1_2 VPW NCH W=0.405u L=0.06u
MNA2 N1 B1 VSS VPW NCH W=0.18u L=0.06u
MNA206 N1_2 A0N VSS VPW NCH W=0.405u L=0.06u
MPA1 INT B0 VDD VNW PCH W=0.22u L=0.06u
MPA108 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA2 INT B1 VDD VNW PCH W=0.22u L=0.06u
MPA2010 Y A0N VDD VNW PCH W=0.49u L=0.06u
.ENDS	AO1B2X0P7MA10TR

****
.SUBCKT AO1B2X1MA10TR  VDD VSS VPW VNW Y   A0N B0 B1
MNA1 INT B0 N1 VPW NCH W=0.24u L=0.06u
MNA104 Y INT N1_2 VPW NCH W=0.575u L=0.06u
MNA2 N1 B1 VSS VPW NCH W=0.24u L=0.06u
MNA206 N1_2 A0N VSS VPW NCH W=0.575u L=0.06u
MPA1 INT B0 VDD VNW PCH W=0.29u L=0.06u
MPA108 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA2 INT B1 VDD VNW PCH W=0.29u L=0.06u
MPA2010 Y A0N VDD VNW PCH W=0.7u L=0.06u
.ENDS	AO1B2X1MA10TR

****

****

****

****

****

****
.SUBCKT AO21BX0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 INT A0 N1 VPW NCH W=0.15u L=0.06u
MNA104 Y B0N N1_2 VPW NCH W=0.29u L=0.06u
MNA2 N1 A1 VSS VPW NCH W=0.15u L=0.06u
MNA206 N1_2 INT VSS VPW NCH W=0.29u L=0.06u
MPA1 INT A0 VDD VNW PCH W=0.185u L=0.06u
MPA108 Y B0N VDD VNW PCH W=0.35u L=0.06u
MPA2 INT A1 VDD VNW PCH W=0.185u L=0.06u
MPA2010 Y INT VDD VNW PCH W=0.35u L=0.06u
.ENDS	AO21BX0P5MA10TR

****
.SUBCKT AO21BX0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 INT A0 N1 VPW NCH W=0.18u L=0.06u
MNA104 Y B0N N1_2 VPW NCH W=0.405u L=0.06u
MNA2 N1 A1 VSS VPW NCH W=0.18u L=0.06u
MNA206 N1_2 INT VSS VPW NCH W=0.405u L=0.06u
MPA1 INT A0 VDD VNW PCH W=0.22u L=0.06u
MPA108 Y B0N VDD VNW PCH W=0.49u L=0.06u
MPA2 INT A1 VDD VNW PCH W=0.22u L=0.06u
MPA2010 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS	AO21BX0P7MA10TR

****
.SUBCKT AO21BX1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 INT A0 N1 VPW NCH W=0.24u L=0.06u
MNA104 Y B0N N1_2 VPW NCH W=0.575u L=0.06u
MNA2 N1 A1 VSS VPW NCH W=0.24u L=0.06u
MNA206 N1_2 INT VSS VPW NCH W=0.575u L=0.06u
MPA1 INT A0 VDD VNW PCH W=0.29u L=0.06u
MPA108 Y B0N VDD VNW PCH W=0.7u L=0.06u
MPA2 INT A1 VDD VNW PCH W=0.29u L=0.06u
MPA2010 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS	AO21BX1MA10TR

****

****

****

****

****

****
.SUBCKT AO21X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA106 INT B0 VSS VPW NCH W=0.15u L=0.06u
MNB1 INT A0 N1 VPW NCH W=0.25u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.25u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA108 INT B0 P1 VNW PCH W=0.365u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.365u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.365u L=0.06u
.ENDS	AO21X0P5MA10TR

****
.SUBCKT AO21X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MNA106 INT B0 VSS VPW NCH W=0.175u L=0.06u
MNB1 INT A0 N1 VPW NCH W=0.29u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.29u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA108 INT B0 P1 VNW PCH W=0.43u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.43u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.43u L=0.06u
.ENDS	AO21X0P7MA10TR

****
.SUBCKT AO21X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MNA106 INT B0 VSS VPW NCH W=0.23u L=0.06u
MNB1 INT A0 N1 VPW NCH W=0.38u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.38u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA108 INT B0 P1 VNW PCH W=0.56u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.56u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.56u L=0.06u
.ENDS	AO21X1MA10TR

****
.SUBCKT AO21X1P4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=0.74u L=0.06u
MNA106 INT B0 VSS VPW NCH W=0.31u L=0.06u
MNB1 INT A0 N1 VPW NCH W=0.515u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.515u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.98u L=0.06u
MPA108 INT B0 P1 VNW PCH W=0.76u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.76u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.76u L=0.06u
.ENDS	AO21X1P4MA10TR

****

****

****

****
.SUBCKT AO21X6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=3.18u L=0.06u
MNA106 INT B0 VSS VPW NCH W=1.245u L=0.06u
MNB1 INT A0 N1 VPW NCH W=2.06u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=2.06u L=0.06u
MPA1 Y INT VDD VNW PCH W=4.2u L=0.06u
MPA108 INT B0 P1 VNW PCH W=3.04u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=3.04u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=3.04u L=0.06u
.ENDS	AO21X6MA10TR

****
.SUBCKT AO22X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA106 INT B0 N1A VPW NCH W=0.255u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=0.255u L=0.06u
MNB1 INT A0 N1B VPW NCH W=0.255u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=0.255u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA109 INT B0 P1 VNW PCH W=0.385u L=0.06u
MPA2 INT B1 P1 VNW PCH W=0.385u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.385u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.385u L=0.06u
.ENDS	AO22X0P5MA10TR

****
.SUBCKT AO22X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MNA106 INT B0 N1A VPW NCH W=0.315u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=0.315u L=0.06u
MNB1 INT A0 N1B VPW NCH W=0.315u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=0.315u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA109 INT B0 P1 VNW PCH W=0.47u L=0.06u
MPA2 INT B1 P1 VNW PCH W=0.47u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.47u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.47u L=0.06u
.ENDS	AO22X0P7MA10TR

****
.SUBCKT AO22X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MNA106 INT B0 N1A VPW NCH W=0.4u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=0.4u L=0.06u
MNB1 INT A0 N1B VPW NCH W=0.4u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=0.4u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA109 INT B0 P1 VNW PCH W=0.6u L=0.06u
MPA2 INT B1 P1 VNW PCH W=0.6u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.6u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.6u L=0.06u
.ENDS	AO22X1MA10TR

****

****

****
.SUBCKT AO22X3MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y INT VSS VPW NCH W=1.59u L=0.06u
MNA106 INT B0 N1A VPW NCH W=1.08u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=1.08u L=0.06u
MNB1 INT A0 N1B VPW NCH W=1.08u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=1.08u L=0.06u
MPA1 Y INT VDD VNW PCH W=2.1u L=0.06u
MPA109 INT B0 P1 VNW PCH W=1.635u L=0.06u
MPA2 INT B1 P1 VNW PCH W=1.635u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=1.635u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=1.635u L=0.06u
.ENDS	AO22X3MA10TR

****
.SUBCKT AO22X4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y INT VSS VPW NCH W=2.12u L=0.06u
MNA106 INT B0 N1A VPW NCH W=1.395u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=1.395u L=0.06u
MNB1 INT A0 N1B VPW NCH W=1.395u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=1.395u L=0.06u
MPA1 Y INT VDD VNW PCH W=2.8u L=0.06u
MPA109 INT B0 P1 VNW PCH W=2.1u L=0.06u
MPA2 INT B1 P1 VNW PCH W=2.1u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.1u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.1u L=0.06u
.ENDS	AO22X4MA10TR

****
.SUBCKT AO22X6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y INT VSS VPW NCH W=3.18u L=0.06u
MNA106 INT B0 N1A VPW NCH W=2.15u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=2.15u L=0.06u
MNB1 INT A0 N1B VPW NCH W=2.15u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=2.15u L=0.06u
MPA1 Y INT VDD VNW PCH W=4.2u L=0.06u
MPA109 INT B0 P1 VNW PCH W=3.25u L=0.06u
MPA2 INT B1 P1 VNW PCH W=3.25u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=3.25u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=3.25u L=0.06u
.ENDS	AO22X6MA10TR

****
.SUBCKT AOI211X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 C0
MN0 Y C0 VSS VPW NCH W=0.15u L=0.06u
MN3 Y B0 VSS VPW NCH W=0.15u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.165u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.165u L=0.06u
MP1 Y C0 NET045 VNW PCH W=0.35u L=0.06u
MP2 NET045 B0 P1 VNW PCH W=0.35u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.35u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.35u L=0.06u
.ENDS	AOI211X0P5MA10TR

****
.SUBCKT AOI211X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 C0
MN0 Y C0 VSS VPW NCH W=0.15u L=0.06u
MN3 Y B0 VSS VPW NCH W=0.15u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.24u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.24u L=0.06u
MP1 Y C0 NET045 VNW PCH W=0.51u L=0.06u
MP2 NET045 B0 P1 VNW PCH W=0.51u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.51u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.51u L=0.06u
.ENDS	AOI211X0P7MA10TR

****
.SUBCKT AOI211X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 C0
MN0 Y C0 VSS VPW NCH W=0.205u L=0.06u
MN3 Y B0 VSS VPW NCH W=0.205u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.33u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.33u L=0.06u
MP1 Y C0 NET045 VNW PCH W=0.7u L=0.06u
MP2 NET045 B0 P1 VNW PCH W=0.7u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
.ENDS	AOI211X1MA10TR

****

****

****

****

****
.SUBCKT AOI21BX0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.15u L=0.06u
MNA106 Y NET28 VSS VPW NCH W=0.15u L=0.06u
MNB1 Y A0 N1 VPW NCH W=0.24u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.24u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.2u L=0.06u
MPA108 Y NET28 P1 VNW PCH W=0.37u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.37u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.37u L=0.06u
.ENDS	AOI21BX0P5MA10TR

****
.SUBCKT AOI21BX0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.15u L=0.06u
MNA106 Y NET28 VSS VPW NCH W=0.2u L=0.06u
MNB1 Y A0 N1 VPW NCH W=0.32u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.32u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.2u L=0.06u
MPA108 Y NET28 P1 VNW PCH W=0.49u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
.ENDS	AOI21BX0P7MA10TR

****
.SUBCKT AOI21BX1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.15u L=0.06u
MNA106 Y NET28 VSS VPW NCH W=0.285u L=0.06u
MNB1 Y A0 N1 VPW NCH W=0.455u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.2u L=0.06u
MPA108 Y NET28 P1 VNW PCH W=0.7u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
.ENDS	AOI21BX1MA10TR

****

****

****
.SUBCKT AOI21BX3MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.415u L=0.06u
MNA106 Y NET28 VSS VPW NCH W=0.855u L=0.06u
MNB1 Y A0 N1 VPW NCH W=1.365u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.365u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.55u L=0.06u
MPA108 Y NET28 P1 VNW PCH W=2.1u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.1u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.1u L=0.06u
.ENDS	AOI21BX3MA10TR

****
.SUBCKT AOI21BX4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.53u L=0.06u
MNA106 Y NET28 VSS VPW NCH W=1.14u L=0.06u
MNB1 Y A0 N1 VPW NCH W=1.82u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.82u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.7u L=0.06u
MPA108 Y NET28 P1 VNW PCH W=2.8u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.8u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.8u L=0.06u
.ENDS	AOI21BX4MA10TR

****
.SUBCKT AOI21BX6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.82u L=0.06u
MNA106 Y NET28 VSS VPW NCH W=1.71u L=0.06u
MNB1 Y A0 N1 VPW NCH W=2.73u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=2.73u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=1.08u L=0.06u
MPA108 Y NET28 P1 VNW PCH W=4.2u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=4.2u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=4.2u L=0.06u
.ENDS	AOI21BX6MA10TR

****
.SUBCKT AOI21BX8MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=1.06u L=0.06u
MNA106 Y NET28 VSS VPW NCH W=2.28u L=0.06u
MNB1 Y A0 N1 VPW NCH W=3.64u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=3.64u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=1.4u L=0.06u
MPA108 Y NET28 P1 VNW PCH W=5.6u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=5.6u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=5.6u L=0.06u
.ENDS	AOI21BX8MA10TR

****
.SUBCKT AOI21X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 VSS VPW NCH W=0.15u L=0.06u
MNB1 Y A0 N1 VPW NCH W=0.24u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.24u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.37u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.37u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.37u L=0.06u
.ENDS	AOI21X0P5MA10TR

****
.SUBCKT AOI21X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 VSS VPW NCH W=0.2u L=0.06u
MNB1 Y A0 N1 VPW NCH W=0.32u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.32u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.49u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
.ENDS	AOI21X0P7MA10TR

****
.SUBCKT AOI21X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 VSS VPW NCH W=0.285u L=0.06u
MNB1 Y A0 N1 VPW NCH W=0.455u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.7u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
.ENDS	AOI21X1MA10TR

****

****

****
.SUBCKT AOI21X3MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 VSS VPW NCH W=0.855u L=0.06u
MNB1 Y A0 N1 VPW NCH W=1.365u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.365u L=0.06u
MPA1 Y B0 P1 VNW PCH W=2.1u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.1u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.1u L=0.06u
.ENDS	AOI21X3MA10TR

****
.SUBCKT AOI21X4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 VSS VPW NCH W=1.14u L=0.06u
MNB1 Y A0 N1 VPW NCH W=1.82u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.82u L=0.06u
MPA1 Y B0 P1 VNW PCH W=2.8u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.8u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.8u L=0.06u
.ENDS	AOI21X4MA10TR

****
.SUBCKT AOI21X6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 VSS VPW NCH W=1.71u L=0.06u
MNB1 Y A0 N1 VPW NCH W=2.73u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=2.73u L=0.06u
MPA1 Y B0 P1 VNW PCH W=4.2u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=4.2u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=4.2u L=0.06u
.ENDS	AOI21X6MA10TR

****
.SUBCKT AOI21X8MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 VSS VPW NCH W=2.28u L=0.06u
MNB1 Y A0 N1 VPW NCH W=3.64u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=3.64u L=0.06u
MPA1 Y B0 P1 VNW PCH W=5.6u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=5.6u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=5.6u L=0.06u
.ENDS	AOI21X8MA10TR

****
.SUBCKT AOI221X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0
MN0 Y C0 VSS VPW NCH W=0.15u L=0.06u
MN2 NET26 B1 VSS VPW NCH W=0.165u L=0.06u
MN3 Y B0 NET26 VPW NCH W=0.165u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.165u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.165u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.35u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.35u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.35u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.35u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.35u L=0.06u
.ENDS	AOI221X0P5MA10TR

****
.SUBCKT AOI221X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0
MN0 Y C0 VSS VPW NCH W=0.15u L=0.06u
MN2 NET26 B1 VSS VPW NCH W=0.24u L=0.06u
MN3 Y B0 NET26 VPW NCH W=0.24u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.24u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.24u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.51u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.51u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.51u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.51u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.51u L=0.06u
.ENDS	AOI221X0P7MA10TR

****
.SUBCKT AOI221X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0
MN0 Y C0 VSS VPW NCH W=0.205u L=0.06u
MN2 NET26 B1 VSS VPW NCH W=0.33u L=0.06u
MN3 Y B0 NET26 VPW NCH W=0.33u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.33u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.33u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.7u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
.ENDS	AOI221X1MA10TR

****
.SUBCKT AOI221X1P4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0
MN0 Y C0 VSS VPW NCH W=0.29u L=0.06u
MN2 NET26 B1 VSS VPW NCH W=0.46u L=0.06u
MN3 Y B0 NET26 VPW NCH W=0.46u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.46u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.46u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.98u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.98u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.98u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.98u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.98u L=0.06u
.ENDS	AOI221X1P4MA10TR

****

****

****

****
.SUBCKT AOI222X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0 C1
MN0 Y C0 NET29 VPW NCH W=0.165u L=0.06u
MN1 NET29 C1 VSS VPW NCH W=0.165u L=0.06u
MN2 NET26 B1 VSS VPW NCH W=0.165u L=0.06u
MN3 Y B0 NET26 VPW NCH W=0.165u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.165u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.165u L=0.06u
MP0 Y C1 P2 VNW PCH W=0.35u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.35u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.35u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.35u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.35u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.35u L=0.06u
.ENDS	AOI222X0P5MA10TR

****
.SUBCKT AOI222X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0 C1
MN0 Y C0 NET29 VPW NCH W=0.23u L=0.06u
MN1 NET29 C1 VSS VPW NCH W=0.23u L=0.06u
MN2 NET26 B1 VSS VPW NCH W=0.23u L=0.06u
MN3 Y B0 NET26 VPW NCH W=0.23u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.23u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.23u L=0.06u
MP0 Y C1 P2 VNW PCH W=0.49u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.49u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.49u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.49u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.49u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.49u L=0.06u
.ENDS	AOI222X0P7MA10TR

****
.SUBCKT AOI222X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0 C1
MN0 Y C0 NET29 VPW NCH W=0.33u L=0.06u
MN1 NET29 C1 VSS VPW NCH W=0.33u L=0.06u
MN2 NET26 B1 VSS VPW NCH W=0.33u L=0.06u
MN3 Y B0 NET26 VPW NCH W=0.33u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.33u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.33u L=0.06u
MP0 Y C1 P2 VNW PCH W=0.7u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.7u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
.ENDS	AOI222X1MA10TR

****
.SUBCKT AOI222X1P4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0 C1
MN0 Y C0 NET29 VPW NCH W=0.46u L=0.06u
MN1 NET29 C1 VSS VPW NCH W=0.46u L=0.06u
MN2 NET26 B1 VSS VPW NCH W=0.46u L=0.06u
MN3 Y B0 NET26 VPW NCH W=0.46u L=0.06u
MN4 Y A0 NET17 VPW NCH W=0.46u L=0.06u
MN5 NET17 A1 VSS VPW NCH W=0.46u L=0.06u
MP0 Y C1 P2 VNW PCH W=0.98u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.98u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.98u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.98u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.98u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.98u L=0.06u
.ENDS	AOI222X1P4MA10TR

****

****

****

****
.SUBCKT AOI22X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1A VPW NCH W=0.24u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=0.24u L=0.06u
MNB1 Y A0 N1B VPW NCH W=0.24u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=0.24u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.37u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.37u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.37u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.37u L=0.06u
.ENDS	AOI22X0P5MA10TR

****
.SUBCKT AOI22X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1A VPW NCH W=0.32u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=0.32u L=0.06u
MNB1 Y A0 N1B VPW NCH W=0.32u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=0.32u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.49u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.49u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
.ENDS	AOI22X0P7MA10TR

****
.SUBCKT AOI22X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1A VPW NCH W=0.455u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=0.455u L=0.06u
MNB1 Y A0 N1B VPW NCH W=0.455u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=0.455u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.7u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.7u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
.ENDS	AOI22X1MA10TR

****

****

****
.SUBCKT AOI22X3MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1A VPW NCH W=1.365u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=1.365u L=0.06u
MNB1 Y A0 N1B VPW NCH W=1.365u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=1.365u L=0.06u
MPA1 Y B0 P1 VNW PCH W=2.1u L=0.06u
MPA2 Y B1 P1 VNW PCH W=2.1u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.1u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.1u L=0.06u
.ENDS	AOI22X3MA10TR

****
.SUBCKT AOI22X4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1A VPW NCH W=1.82u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=1.82u L=0.06u
MNB1 Y A0 N1B VPW NCH W=1.82u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=1.82u L=0.06u
MPA1 Y B0 P1 VNW PCH W=2.8u L=0.06u
MPA2 Y B1 P1 VNW PCH W=2.8u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.8u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.8u L=0.06u
.ENDS	AOI22X4MA10TR

****
.SUBCKT AOI22X6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1A VPW NCH W=2.73u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=2.73u L=0.06u
MNB1 Y A0 N1B VPW NCH W=2.73u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=2.73u L=0.06u
MPA1 Y B0 P1 VNW PCH W=4.2u L=0.06u
MPA2 Y B1 P1 VNW PCH W=4.2u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=4.2u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=4.2u L=0.06u
.ENDS	AOI22X6MA10TR

****
.SUBCKT AOI22X8MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1A VPW NCH W=3.64u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=3.64u L=0.06u
MNB1 Y A0 N1B VPW NCH W=3.64u L=0.06u
MNB2 N1B A1 VSS VPW NCH W=3.64u L=0.06u
MPA1 Y B0 P1 VNW PCH W=5.6u L=0.06u
MPA2 Y B1 P1 VNW PCH W=5.6u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=5.6u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=5.6u L=0.06u
.ENDS	AOI22X8MA10TR

****
.SUBCKT AOI2XB1X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.155u L=0.06u
MNA106 Y B0 VSS VPW NCH W=0.15u L=0.06u
MNB1 Y A0 N1 VPW NCH W=0.24u L=0.06u
MNB2 N1 INT VSS VPW NCH W=0.24u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.205u L=0.06u
MPA108 Y B0 P1 VNW PCH W=0.37u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.37u L=0.06u
MPB2 P1 INT VDD VNW PCH W=0.37u L=0.06u
.ENDS	AOI2XB1X0P5MA10TR

****
.SUBCKT AOI2XB1X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.155u L=0.06u
MNA106 Y B0 VSS VPW NCH W=0.2u L=0.06u
MNB1 Y A0 N1 VPW NCH W=0.32u L=0.06u
MNB2 N1 INT VSS VPW NCH W=0.32u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.205u L=0.06u
MPA108 Y B0 P1 VNW PCH W=0.49u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MPB2 P1 INT VDD VNW PCH W=0.49u L=0.06u
.ENDS	AOI2XB1X0P7MA10TR

****
.SUBCKT AOI2XB1X1MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.155u L=0.06u
MNA106 Y B0 VSS VPW NCH W=0.285u L=0.06u
MNB1 Y A0 N1 VPW NCH W=0.455u L=0.06u
MNB2 N1 INT VSS VPW NCH W=0.455u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.205u L=0.06u
MPA108 Y B0 P1 VNW PCH W=0.7u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MPB2 P1 INT VDD VNW PCH W=0.7u L=0.06u
.ENDS	AOI2XB1X1MA10TR

****

****

****
.SUBCKT AOI2XB1X3MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.455u L=0.06u
MNA106 Y B0 VSS VPW NCH W=0.855u L=0.06u
MNB1 Y A0 N1 VPW NCH W=1.365u L=0.06u
MNB2 N1 INT VSS VPW NCH W=1.365u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.6u L=0.06u
MPA108 Y B0 P1 VNW PCH W=2.1u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.1u L=0.06u
MPB2 P1 INT VDD VNW PCH W=2.1u L=0.06u
.ENDS	AOI2XB1X3MA10TR

****
.SUBCKT AOI2XB1X4MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.59u L=0.06u
MNA106 Y B0 VSS VPW NCH W=1.14u L=0.06u
MNB1 Y A0 N1 VPW NCH W=1.82u L=0.06u
MNB2 N1 INT VSS VPW NCH W=1.82u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.78u L=0.06u
MPA108 Y B0 P1 VNW PCH W=2.8u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.8u L=0.06u
MPB2 P1 INT VDD VNW PCH W=2.8u L=0.06u
.ENDS	AOI2XB1X4MA10TR

****
.SUBCKT AOI2XB1X6MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.89u L=0.06u
MNA106 Y B0 VSS VPW NCH W=1.71u L=0.06u
MNB1 Y A0 N1 VPW NCH W=2.73u L=0.06u
MNB2 N1 INT VSS VPW NCH W=2.73u L=0.06u
MPA1 INT A1N VDD VNW PCH W=1.18u L=0.06u
MPA108 Y B0 P1 VNW PCH W=4.2u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=4.2u L=0.06u
MPB2 P1 INT VDD VNW PCH W=4.2u L=0.06u
.ENDS	AOI2XB1X6MA10TR

****
.SUBCKT AOI2XB1X8MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=1.185u L=0.06u
MNA106 Y B0 VSS VPW NCH W=2.28u L=0.06u
MNB1 Y A0 N1 VPW NCH W=3.64u L=0.06u
MNB2 N1 INT VSS VPW NCH W=3.64u L=0.06u
MPA1 INT A1N VDD VNW PCH W=1.56u L=0.06u
MPA108 Y B0 P1 VNW PCH W=5.6u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=5.6u L=0.06u
MPB2 P1 INT VDD VNW PCH W=5.6u L=0.06u
.ENDS	AOI2XB1X8MA10TR

****
.SUBCKT AOI31X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0
MNA1 Y B0 VSS VPW NCH W=0.15u L=0.06u
MNB1 Y A0 N2 VPW NCH W=0.32u L=0.06u
MNB2 N2 A1 N1 VPW NCH W=0.32u L=0.06u
MNB3 N1 A2 VSS VPW NCH W=0.32u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.37u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.37u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.37u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=0.37u L=0.06u
.ENDS	AOI31X0P5MA10TR

****
.SUBCKT AOI31X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0
MNA1 Y B0 VSS VPW NCH W=0.19u L=0.06u
MNB1 Y A0 N2 VPW NCH W=0.405u L=0.06u
MNB2 N2 A1 N1 VPW NCH W=0.405u L=0.06u
MNB3 N1 A2 VSS VPW NCH W=0.405u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.465u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.465u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.465u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=0.465u L=0.06u
.ENDS	AOI31X0P7MA10TR

****
.SUBCKT AOI31X1MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0
MNA1 Y B0 VSS VPW NCH W=0.27u L=0.06u
MNB1 Y A0 N2 VPW NCH W=0.58u L=0.06u
MNB2 N2 A1 N1 VPW NCH W=0.58u L=0.06u
MNB3 N1 A2 VSS VPW NCH W=0.58u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.665u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.665u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.665u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=0.665u L=0.06u
.ENDS	AOI31X1MA10TR

****
.SUBCKT AOI31X1P4MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0
MNA1 Y B0 VSS VPW NCH W=0.38u L=0.06u
MNB1 Y A0 N2 VPW NCH W=0.81u L=0.06u
MNB2 N2 A1 N1 VPW NCH W=0.81u L=0.06u
MNB3 N1 A2 VSS VPW NCH W=0.81u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.93u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.93u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.93u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=0.93u L=0.06u
.ENDS	AOI31X1P4MA10TR

****
.SUBCKT AOI31X2MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0
MNA1 Y B0 VSS VPW NCH W=0.54u L=0.06u
MNB1 Y A0 N2 VPW NCH W=1.16u L=0.06u
MNB2 N2 A1 N1 VPW NCH W=1.16u L=0.06u
MNB3 N1 A2 VSS VPW NCH W=1.16u L=0.06u
MPA1 Y B0 P1 VNW PCH W=1.33u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=1.33u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=1.33u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=1.33u L=0.06u
.ENDS	AOI31X2MA10TR

****
.SUBCKT AOI31X3MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0
MNA1 Y B0 VSS VPW NCH W=0.81u L=0.06u
MNB1 Y A0 N2 VPW NCH W=1.74u L=0.06u
MNB2 N2 A1 N1 VPW NCH W=1.74u L=0.06u
MNB3 N1 A2 VSS VPW NCH W=1.74u L=0.06u
MPA1 Y B0 P1 VNW PCH W=1.995u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=1.995u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=1.995u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=1.995u L=0.06u
.ENDS	AOI31X3MA10TR

****
.SUBCKT AOI31X4MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0
MNA1 Y B0 VSS VPW NCH W=1.08u L=0.06u
MNB1 Y A0 N2 VPW NCH W=2.32u L=0.06u
MNB2 N2 A1 N1 VPW NCH W=2.32u L=0.06u
MNB3 N1 A2 VSS VPW NCH W=2.32u L=0.06u
MPA1 Y B0 P1 VNW PCH W=2.66u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.66u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.66u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=2.66u L=0.06u
.ENDS	AOI31X4MA10TR

****
.SUBCKT AOI31X6MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0
MNA1 Y B0 VSS VPW NCH W=1.62u L=0.06u
MNB1 Y A0 N2 VPW NCH W=3.48u L=0.06u
MNB2 N2 A1 N1 VPW NCH W=3.48u L=0.06u
MNB3 N1 A2 VSS VPW NCH W=3.48u L=0.06u
MPA1 Y B0 P1 VNW PCH W=3.99u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=3.99u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=3.99u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=3.99u L=0.06u
.ENDS	AOI31X6MA10TR

****
.SUBCKT AOI32X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0 B1
MNA1 Y B0 N1A VPW NCH W=0.22u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=0.22u L=0.06u
MNB1 Y A0 N2B VPW NCH W=0.29u L=0.06u
MNB2 N2B A1 N1B VPW NCH W=0.29u L=0.06u
MNB3 N1B A2 VSS VPW NCH W=0.29u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.335u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.335u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.335u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.335u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=0.335u L=0.06u
.ENDS	AOI32X0P5MA10TR

****
.SUBCKT AOI32X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0 B1
MNA1 Y B0 N1A VPW NCH W=0.305u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=0.305u L=0.06u
MNB1 Y A0 N2B VPW NCH W=0.405u L=0.06u
MNB2 N2B A1 N1B VPW NCH W=0.405u L=0.06u
MNB3 N1B A2 VSS VPW NCH W=0.405u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.465u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.465u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.465u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.465u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=0.465u L=0.06u
.ENDS	AOI32X0P7MA10TR

****
.SUBCKT AOI32X1MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0 B1
MNA1 Y B0 N1A VPW NCH W=0.435u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=0.435u L=0.06u
MNB1 Y A0 N2B VPW NCH W=0.58u L=0.06u
MNB2 N2B A1 N1B VPW NCH W=0.58u L=0.06u
MNB3 N1B A2 VSS VPW NCH W=0.58u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.665u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.665u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.665u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.665u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=0.665u L=0.06u
.ENDS	AOI32X1MA10TR

****

****

****
.SUBCKT AOI32X3MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0 B1
MNA1 Y B0 N1A VPW NCH W=1.305u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=1.305u L=0.06u
MNB1 Y A0 N2B VPW NCH W=1.74u L=0.06u
MNB2 N2B A1 N1B VPW NCH W=1.74u L=0.06u
MNB3 N1B A2 VSS VPW NCH W=1.74u L=0.06u
MPA1 Y B0 P1 VNW PCH W=1.995u L=0.06u
MPA2 Y B1 P1 VNW PCH W=1.995u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=1.995u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=1.995u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=1.995u L=0.06u
.ENDS	AOI32X3MA10TR

****
.SUBCKT AOI32X4MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0 B1
MNA1 Y B0 N1A VPW NCH W=1.74u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=1.74u L=0.06u
MNB1 Y A0 N2B VPW NCH W=2.32u L=0.06u
MNB2 N2B A1 N1B VPW NCH W=2.32u L=0.06u
MNB3 N1B A2 VSS VPW NCH W=2.32u L=0.06u
MPA1 Y B0 P1 VNW PCH W=2.66u L=0.06u
MPA2 Y B1 P1 VNW PCH W=2.66u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=2.66u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.66u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=2.66u L=0.06u
.ENDS	AOI32X4MA10TR

****
.SUBCKT AOI32X6MA10TR  VDD VSS VPW VNW Y   A0 A1 A2 B0 B1
MNA1 Y B0 N1A VPW NCH W=2.61u L=0.06u
MNA2 N1A B1 VSS VPW NCH W=2.61u L=0.06u
MNB1 Y A0 N2B VPW NCH W=3.48u L=0.06u
MNB2 N2B A1 N1B VPW NCH W=3.48u L=0.06u
MNB3 N1B A2 VSS VPW NCH W=3.48u L=0.06u
MPA1 Y B0 P1 VNW PCH W=3.99u L=0.06u
MPA2 Y B1 P1 VNW PCH W=3.99u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=3.99u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=3.99u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=3.99u L=0.06u
.ENDS	AOI32X6MA10TR

****
.SUBCKT BUFHX0P7MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.26u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.37u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.345u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.49u L=0.06u
.ENDS	BUFHX0P7MA10TR

****
.SUBCKT BUFHX0P8MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.29u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.425u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.38u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.56u L=0.06u
.ENDS	BUFHX0P8MA10TR

****
.SUBCKT BUFHX11MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=3.49u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=5.83u L=0.06u
MPA1 NET15 A VDD VNW PCH W=4.58u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=7.7u L=0.06u
.ENDS	BUFHX11MA10TR

****
.SUBCKT BUFHX13MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=4.07u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=6.89u L=0.06u
MPA1 NET15 A VDD VNW PCH W=5.38u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=9.1u L=0.06u
.ENDS	BUFHX13MA10TR

****
.SUBCKT BUFHX16MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=4.96u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=8.48u L=0.06u
MPA1 NET15 A VDD VNW PCH W=6.55u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=11.2u L=0.06u
.ENDS	BUFHX16MA10TR

****
.SUBCKT BUFHX1MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.34u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.53u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.45u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.7u L=0.06u
.ENDS	BUFHX1MA10TR

****
.SUBCKT BUFHX1P2MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.42u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.635u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.56u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.84u L=0.06u
.ENDS	BUFHX1P2MA10TR

****
.SUBCKT BUFHX1P4MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.48u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.74u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.63u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.98u L=0.06u
.ENDS	BUFHX1P4MA10TR

****
.SUBCKT BUFHX1P7MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.53u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.9u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.7u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=1.19u L=0.06u
.ENDS	BUFHX1P7MA10TR

****
.SUBCKT BUFHX2MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.64u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.06u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.84u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=1.4u L=0.06u
.ENDS	BUFHX2MA10TR

****
.SUBCKT BUFHX2P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.83u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.325u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.1u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=1.75u L=0.06u
.ENDS	BUFHX2P5MA10TR

****
.SUBCKT BUFHX3MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.96u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.59u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.27u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=2.1u L=0.06u
.ENDS	BUFHX3MA10TR

****
.SUBCKT BUFHX3P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.13u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.855u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.49u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=2.46u L=0.06u
.ENDS	BUFHX3P5MA10TR

****
.SUBCKT BUFHX4MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.26u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=2.12u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.66u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=2.8u L=0.06u
.ENDS	BUFHX4MA10TR

****
.SUBCKT BUFHX5MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.59u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=2.65u L=0.06u
MPA1 NET15 A VDD VNW PCH W=2.1u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=3.5u L=0.06u
.ENDS	BUFHX5MA10TR

****
.SUBCKT BUFHX6MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.91u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=3.18u L=0.06u
MPA1 NET15 A VDD VNW PCH W=2.49u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=4.2u L=0.06u
.ENDS	BUFHX6MA10TR

****
.SUBCKT BUFHX7P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=2.39u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=3.975u L=0.06u
MPA1 NET15 A VDD VNW PCH W=3.15u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=5.25u L=0.06u
.ENDS	BUFHX7P5MA10TR

****
.SUBCKT BUFHX9MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=2.85u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=4.77u L=0.06u
MPA1 NET15 A VDD VNW PCH W=3.76u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=6.3u L=0.06u
.ENDS	BUFHX9MA10TR

****
.SUBCKT BUFX0P7BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.255u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.29u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.49u L=0.06u
.ENDS	BUFX0P7BA10TR

****
.SUBCKT BUFX0P7MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.37u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.2u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.49u L=0.06u
.ENDS	BUFX0P7MA10TR

****
.SUBCKT BUFX0P8BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.29u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.29u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.56u L=0.06u
.ENDS	BUFX0P8BA10TR

****
.SUBCKT BUFX0P8MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.425u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.2u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.56u L=0.06u
.ENDS	BUFX0P8MA10TR

****
.SUBCKT BUFX11BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.21u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=3.96u L=0.06u
MPA1 NET15 A VDD VNW PCH W=2.345u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=7.7u L=0.06u
.ENDS	BUFX11BA10TR

****
.SUBCKT BUFX11MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.735u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=5.83u L=0.06u
MPA1 NET15 A VDD VNW PCH W=2.29u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=7.7u L=0.06u
.ENDS	BUFX11MA10TR

****
.SUBCKT BUFX13BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.42u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=4.68u L=0.06u
MPA1 NET15 A VDD VNW PCH W=2.755u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=9.1u L=0.06u
.ENDS	BUFX13BA10TR

****
.SUBCKT BUFX13MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=2.035u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=6.89u L=0.06u
MPA1 NET15 A VDD VNW PCH W=2.69u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=9.1u L=0.06u
.ENDS	BUFX13MA10TR

****
.SUBCKT BUFX16BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.73u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=5.76u L=0.06u
MPA1 NET15 A VDD VNW PCH W=3.35u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=11.2u L=0.06u
.ENDS	BUFX16BA10TR

****
.SUBCKT BUFX16MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=2.48u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=8.48u L=0.06u
MPA1 NET15 A VDD VNW PCH W=3.275u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=11.2u L=0.06u
.ENDS	BUFX16MA10TR

****
.SUBCKT BUFX1BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.36u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.29u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.7u L=0.06u
.ENDS	BUFX1BA10TR

****
.SUBCKT BUFX1MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.17u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.53u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.225u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.7u L=0.06u
.ENDS	BUFX1MA10TR

****
.SUBCKT BUFX1P2BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.43u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.29u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.84u L=0.06u
.ENDS	BUFX1P2BA10TR

****
.SUBCKT BUFX1P2MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.21u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.635u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.28u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.84u L=0.06u
.ENDS	BUFX1P2MA10TR

****
.SUBCKT BUFX1P4BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.165u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.505u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.325u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.98u L=0.06u
.ENDS	BUFX1P4BA10TR

****
.SUBCKT BUFX1P4MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.24u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.74u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.315u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=0.98u L=0.06u
.ENDS	BUFX1P4MA10TR

****
.SUBCKT BUFX1P7BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.195u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.61u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.375u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=1.19u L=0.06u
.ENDS	BUFX1P7BA10TR

****
.SUBCKT BUFX1P7MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.275u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.9u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.365u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=1.19u L=0.06u
.ENDS	BUFX1P7MA10TR

****
.SUBCKT BUFX2BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.22u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.72u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.43u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=1.4u L=0.06u
.ENDS	BUFX2BA10TR

****
.SUBCKT BUFX2MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.32u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.06u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.42u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=1.4u L=0.06u
.ENDS	BUFX2MA10TR

****
.SUBCKT BUFX2P5BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.29u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=0.9u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.565u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=1.75u L=0.06u
.ENDS	BUFX2P5BA10TR

****
.SUBCKT BUFX2P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.415u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.325u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.55u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=1.75u L=0.06u
.ENDS	BUFX2P5MA10TR

****
.SUBCKT BUFX3BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.335u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.08u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.65u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=2.1u L=0.06u
.ENDS	BUFX3BA10TR

****
.SUBCKT BUFX3MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.48u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.59u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.635u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=2.1u L=0.06u
.ENDS	BUFX3MA10TR

****
.SUBCKT BUFX3P5BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.395u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.26u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.765u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=2.46u L=0.06u
.ENDS	BUFX3P5BA10TR

****
.SUBCKT BUFX3P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.565u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.855u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.745u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=2.46u L=0.06u
.ENDS	BUFX3P5MA10TR

****
.SUBCKT BUFX4BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.44u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.44u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.855u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=2.8u L=0.06u
.ENDS	BUFX4BA10TR

****
.SUBCKT BUFX4MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.63u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=2.12u L=0.06u
MPA1 NET15 A VDD VNW PCH W=0.83u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=2.8u L=0.06u
.ENDS	BUFX4MA10TR

****
.SUBCKT BUFX5BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.555u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=1.8u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.08u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=3.5u L=0.06u
.ENDS	BUFX5BA10TR

****
.SUBCKT BUFX5MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.795u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=2.65u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.05u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=3.5u L=0.06u
.ENDS	BUFX5MA10TR

****
.SUBCKT BUFX6BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.655u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=2.16u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.275u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=4.2u L=0.06u
.ENDS	BUFX6BA10TR

****
.SUBCKT BUFX6MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.945u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=3.18u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.245u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=4.2u L=0.06u
.ENDS	BUFX6MA10TR

****
.SUBCKT BUFX7P5BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.835u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=2.7u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.615u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=5.25u L=0.06u
.ENDS	BUFX7P5BA10TR

****
.SUBCKT BUFX7P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.195u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=3.975u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.575u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=5.25u L=0.06u
.ENDS	BUFX7P5MA10TR

****
.SUBCKT BUFX9BA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=0.995u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=3.24u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.93u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=6.3u L=0.06u
.ENDS	BUFX9BA10TR

****
.SUBCKT BUFX9MA10TR  VDD VSS VPW VNW Y   A
MNA1 NET15 A VSS VPW NCH W=1.425u L=0.06u
MNA102 Y NET15 VSS VPW NCH W=4.77u L=0.06u
MPA1 NET15 A VDD VNW PCH W=1.88u L=0.06u
MPA104 Y NET15 VDD VNW PCH W=6.3u L=0.06u
.ENDS	BUFX9MA10TR

****
.SUBCKT BUFZX11MA10TR  VDD VSS VPW VNW Y   OE A
MN0 Y NET015 VSS VPW NCH W=6.05u L=0.06u
MN1 NET015 NEN VSS VPW NCH W=1.215u L=0.06u
MN2 NET015 A VSS VPW NCH W=2.9u L=0.06u
MN4 NET014 OE NET015 VPW NCH W=1.44u L=0.06u
MNA1 NEN OE VSS VPW NCH W=0.86u L=0.06u
MP0 Y NET014 VDD VNW PCH W=7.7u L=0.06u
MP1 NET014 OE VDD VNW PCH W=1.65u L=0.06u
MP3 NET014 A VDD VNW PCH W=4.2u L=0.06u
MP6 NET015 NEN NET014 VNW PCH W=2.1u L=0.06u
MPA1 NEN OE VDD VNW PCH W=1.14u L=0.06u
.ENDS	BUFZX11MA10TR

****
.SUBCKT BUFZX16MA10TR  VDD VSS VPW VNW Y   OE A
MN0 Y NET015 VSS VPW NCH W=8.8u L=0.06u
MN1 NET015 NEN VSS VPW NCH W=1.71u L=0.06u
MN2 NET015 A VSS VPW NCH W=4.06u L=0.06u
MN4 NET014 OE NET015 VPW NCH W=2.02u L=0.06u
MNA1 NEN OE VSS VPW NCH W=1.185u L=0.06u
MP0 Y NET014 VDD VNW PCH W=11.2u L=0.06u
MP1 NET014 OE VDD VNW PCH W=2.3u L=0.06u
MP3 NET014 A VDD VNW PCH W=5.895u L=0.06u
MP6 NET015 NEN NET014 VNW PCH W=2.95u L=0.06u
MPA1 NEN OE VDD VNW PCH W=1.575u L=0.06u
.ENDS	BUFZX16MA10TR

****
.SUBCKT BUFZX1MA10TR  VDD VSS VPW VNW Y   OE A
MN0 Y NET015 VSS VPW NCH W=0.55u L=0.06u
MN1 NET015 NEN VSS VPW NCH W=0.15u L=0.06u
MN2 NET015 A VSS VPW NCH W=0.36u L=0.06u
MN4 NET014 OE NET015 VPW NCH W=0.18u L=0.06u
MNA1 NEN OE VSS VPW NCH W=0.15u L=0.06u
MP0 Y NET014 VDD VNW PCH W=0.7u L=0.06u
MP1 NET014 OE VDD VNW PCH W=0.2u L=0.06u
MP3 NET014 A VDD VNW PCH W=0.52u L=0.06u
MP6 NET015 NEN NET014 VNW PCH W=0.26u L=0.06u
MPA1 NEN OE VDD VNW PCH W=0.2u L=0.06u
.ENDS	BUFZX1MA10TR

****
.SUBCKT BUFZX1P4MA10TR  VDD VSS VPW VNW Y   OE A
MN0 Y NET015 VSS VPW NCH W=0.77u L=0.06u
MN1 NET015 NEN VSS VPW NCH W=0.2u L=0.06u
MN2 NET015 A VSS VPW NCH W=0.49u L=0.06u
MN4 NET014 OE NET015 VPW NCH W=0.245u L=0.06u
MNA1 NEN OE VSS VPW NCH W=0.15u L=0.06u
MP0 Y NET014 VDD VNW PCH W=0.98u L=0.06u
MP1 NET014 OE VDD VNW PCH W=0.27u L=0.06u
MP3 NET014 A VDD VNW PCH W=0.7u L=0.06u
MP6 NET015 NEN NET014 VNW PCH W=0.35u L=0.06u
MPA1 NEN OE VDD VNW PCH W=0.2u L=0.06u
.ENDS	BUFZX1P4MA10TR

****
.SUBCKT BUFZX2MA10TR  VDD VSS VPW VNW Y   OE A
MN0 Y NET015 VSS VPW NCH W=1.1u L=0.06u
MN1 NET015 NEN VSS VPW NCH W=0.27u L=0.06u
MN2 NET015 A VSS VPW NCH W=0.67u L=0.06u
MN4 NET014 OE NET015 VPW NCH W=0.335u L=0.06u
MNA1 NEN OE VSS VPW NCH W=0.155u L=0.06u
MP0 Y NET014 VDD VNW PCH W=1.4u L=0.06u
MP1 NET014 OE VDD VNW PCH W=0.37u L=0.06u
MP3 NET014 A VDD VNW PCH W=0.95u L=0.06u
MP6 NET015 NEN NET014 VNW PCH W=0.475u L=0.06u
MPA1 NEN OE VDD VNW PCH W=0.205u L=0.06u
.ENDS	BUFZX2MA10TR

****
.SUBCKT BUFZX3MA10TR  VDD VSS VPW VNW Y   OE A
MN0 Y NET015 VSS VPW NCH W=1.65u L=0.06u
MN1 NET015 NEN VSS VPW NCH W=0.39u L=0.06u
MN2 NET015 A VSS VPW NCH W=0.97u L=0.06u
MN4 NET014 OE NET015 VPW NCH W=0.485u L=0.06u
MNA1 NEN OE VSS VPW NCH W=0.285u L=0.06u
MP0 Y NET014 VDD VNW PCH W=2.1u L=0.06u
MP1 NET014 OE VDD VNW PCH W=0.54u L=0.06u
MP3 NET014 A VDD VNW PCH W=1.38u L=0.06u
MP6 NET015 NEN NET014 VNW PCH W=0.69u L=0.06u
MPA1 NEN OE VDD VNW PCH W=0.38u L=0.06u
.ENDS	BUFZX3MA10TR

****
.SUBCKT BUFZX4MA10TR  VDD VSS VPW VNW Y   OE A
MN0 Y NET015 VSS VPW NCH W=2.2u L=0.06u
MN1 NET015 NEN VSS VPW NCH W=0.49u L=0.06u
MN2 NET015 A VSS VPW NCH W=1.215u L=0.06u
MN4 NET014 OE NET015 VPW NCH W=0.61u L=0.06u
MNA1 NEN OE VSS VPW NCH W=0.35u L=0.06u
MP0 Y NET014 VDD VNW PCH W=2.8u L=0.06u
MP1 NET014 OE VDD VNW PCH W=0.675u L=0.06u
MP3 NET014 A VDD VNW PCH W=1.725u L=0.06u
MP6 NET015 NEN NET014 VNW PCH W=0.86u L=0.06u
MPA1 NEN OE VDD VNW PCH W=0.47u L=0.06u
.ENDS	BUFZX4MA10TR

****
.SUBCKT BUFZX6MA10TR  VDD VSS VPW VNW Y   OE A
MN0 Y NET015 VSS VPW NCH W=3.3u L=0.06u
MN1 NET015 NEN VSS VPW NCH W=0.69u L=0.06u
MN2 NET015 A VSS VPW NCH W=1.72u L=0.06u
MN4 NET014 OE NET015 VPW NCH W=0.86u L=0.06u
MNA1 NEN OE VSS VPW NCH W=0.5u L=0.06u
MP0 Y NET014 VDD VNW PCH W=4.2u L=0.06u
MP1 NET014 OE VDD VNW PCH W=0.95u L=0.06u
MP3 NET014 A VDD VNW PCH W=2.42u L=0.06u
MP6 NET015 NEN NET014 VNW PCH W=1.21u L=0.06u
MPA1 NEN OE VDD VNW PCH W=0.66u L=0.06u
.ENDS	BUFZX6MA10TR

****
.SUBCKT BUFZX8MA10TR  VDD VSS VPW VNW Y   OE A
MN0 Y NET015 VSS VPW NCH W=4.4u L=0.06u
MN1 NET015 NEN VSS VPW NCH W=0.9u L=0.06u
MN2 NET015 A VSS VPW NCH W=2.24u L=0.06u
MN4 NET014 OE NET015 VPW NCH W=1.12u L=0.06u
MNA1 NEN OE VSS VPW NCH W=0.65u L=0.06u
MP0 Y NET014 VDD VNW PCH W=5.6u L=0.06u
MP1 NET014 OE VDD VNW PCH W=1.23u L=0.06u
MP3 NET014 A VDD VNW PCH W=3.15u L=0.06u
MP6 NET015 NEN NET014 VNW PCH W=1.575u L=0.06u
MPA1 NEN OE VDD VNW PCH W=0.86u L=0.06u
.ENDS	BUFZX8MA10TR

****
.SUBCKT DFFNQX1MA10TR  VDD VSS VPW VNW Q   CKN D
MNA1 NCLK_ CKN VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 NET86 D VSS VPW NCH W=0.2u L=0.06u
MNA1024 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.3u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.2u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.35u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.15u L=0.06u
MNOE016 S BCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK_ N1_9 VPW NCH W=0.15u L=0.06u
MNOE036 NM BCLK_ NET86 VPW NCH W=0.15u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.35u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 NET86 D VDD VNW PCH W=0.5u L=0.06u
MPA1026 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.45u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.25u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.45u L=0.06u
MPOEN018 S NCLK_ P1 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK_ P1_11 VNW PCH W=0.15u L=0.06u
MPOEN038 NM NCLK_ NET86 VNW PCH W=0.45u L=0.06u
.ENDS	DFFNQX1MA10TR

****
.SUBCKT DFFNQX2MA10TR  VDD VSS VPW VNW Q   CKN D
MNA1 NCLK_ CKN VSS VPW NCH W=0.16u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 NET80 D VSS VPW NCH W=0.3u L=0.06u
MNA1024 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.4u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.24u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.58u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.2u L=0.06u
MNOE016 S BCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK_ N1_9 VPW NCH W=0.15u L=0.06u
MNOE036 NM BCLK_ NET80 VPW NCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.32u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.58u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 NET80 D VDD VNW PCH W=0.7u L=0.06u
MPA1026 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.6u L=0.06u
MPA1042 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.3u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.6u L=0.06u
MPOEN018 S NCLK_ P1 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK_ P1_11 VNW PCH W=0.15u L=0.06u
MPOEN038 NM NCLK_ NET80 VNW PCH W=0.6u L=0.06u
.ENDS	DFFNQX2MA10TR

****
.SUBCKT DFFNQX3MA10TR  VDD VSS VPW VNW Q   CKN D
MNA1 NCLK_ CKN VSS VPW NCH W=0.18u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 NET85 D VSS VPW NCH W=0.3u L=0.06u
MNA1024 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.45u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.28u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA108 NS S VSS VPW NCH W=0.58u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.25u L=0.06u
MNOE016 S BCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK_ N1_9 VPW NCH W=0.15u L=0.06u
MNOE036 NM BCLK_ NET85 VPW NCH W=0.25u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.36u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.58u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 NET85 D VDD VNW PCH W=0.7u L=0.06u
MPA1026 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1042 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.34u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.7u L=0.06u
MPOEN018 S NCLK_ P1 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK_ P1_11 VNW PCH W=0.15u L=0.06u
MPOEN038 NM NCLK_ NET85 VNW PCH W=0.7u L=0.06u
.ENDS	DFFNQX3MA10TR

****
.SUBCKT DFFNRPQX1MA10TR  VDD VSS VPW VNW Q   CKN R D
MN2 NET47 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.15u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.15u L=0.06u
MNA1014 M R VSS VPW NCH W=0.2u L=0.06u
MNA1024 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 NIN D VSS VPW NCH W=0.2u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.2u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.36u L=0.06u
MNA2 M NM VSS VPW NCH W=0.2u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE032 NM BCLK_ NIN VPW NCH W=0.15u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.36u L=0.06u
MPA1017 M R P1 VNW PCH W=0.6u L=0.06u
MPA1026 P1_12 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NIN D VDD VNW PCH W=0.5u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.25u L=0.06u
MPA2 P1 NM VDD VNW PCH W=0.6u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.445u L=0.06u
MPOEN030 NM BCLK_ P1_12 VNW PCH W=0.15u L=0.06u
MPOEN034 NM NCLK_ NIN VNW PCH W=0.45u L=0.06u
.ENDS	DFFNRPQX1MA10TR

****
.SUBCKT DFFNRPQX2MA10TR  VDD VSS VPW VNW Q   CKN R D
MN2 NET47 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.15u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.16u L=0.06u
MNA1014 M R VSS VPW NCH W=0.3u L=0.06u
MNA1024 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.24u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.58u L=0.06u
MNA2 M NM VSS VPW NCH W=0.3u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.2u L=0.06u
MNOE028 NM NCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE032 NM BCLK_ NIN VPW NCH W=0.2u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.32u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.58u L=0.06u
MPA1017 M R P1 VNW PCH W=0.8u L=0.06u
MPA1026 P1_12 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1042 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.3u L=0.06u
MPA2 P1 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.6u L=0.06u
MPOEN030 NM BCLK_ P1_12 VNW PCH W=0.15u L=0.06u
MPOEN034 NM NCLK_ NIN VNW PCH W=0.6u L=0.06u
.ENDS	DFFNRPQX2MA10TR

****
.SUBCKT DFFNRPQX3MA10TR  VDD VSS VPW VNW Q   CKN R D
MN7 S R VSS VPW NCH W=0.15u L=0.06u
MN8 S BCLK_ NET49 VPW NCH W=0.15u L=0.06u
MN9 NET49 NS VSS VPW NCH W=0.15u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.18u L=0.06u
MNA1010 M R VSS VPW NCH W=0.3u L=0.06u
MNA102 BCLK_ NCLK_ VSS VPW NCH W=0.28u L=0.06u
MNA1020 NET0113 D VSS VPW NCH W=0.3u L=0.06u
MNA1025 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1039 NS S VSS VPW NCH W=0.58u L=0.06u
MNA106 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA2 M NM VSS VPW NCH W=0.3u L=0.06u
MNOE NM NCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE031 NM BCLK_ NET0113 VPW NCH W=0.25u L=0.06u
MNOE035 S NCLK_ M VPW NCH W=0.25u L=0.06u
MP10 NET69 NS NET63 VNW PCH W=0.2u L=0.06u
MP8 S NCLK_ NET69 VNW PCH W=0.2u L=0.06u
MP9 NET63 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.36u L=0.06u
MPA1013 M R P1 VNW PCH W=0.8u L=0.06u
MPA1022 NET0113 D VDD VNW PCH W=0.7u L=0.06u
MPA1027 P1_12 M VDD VNW PCH W=0.15u L=0.06u
MPA104 BCLK_ NCLK_ VDD VNW PCH W=0.34u L=0.06u
MPA1041 NS S VDD VNW PCH W=0.58u L=0.06u
MPA108 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA2 P1 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN NM BCLK_ P1_12 VNW PCH W=0.15u L=0.06u
MPOEN033 NM NCLK_ NET0113 VNW PCH W=0.7u L=0.06u
MPOEN037 S BCLK_ M VNW PCH W=0.65u L=0.06u
.ENDS	DFFNRPQX3MA10TR

****
.SUBCKT DFFNSQX1MA10TR  VDD VSS VPW VNW Q   CKN D SN
MN2 NET50 NS NET47 VPW NCH W=0.2u L=0.06u
MN3 NET47 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET50 VPW NCH W=0.2u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1030 NMUX D VSS VPW NCH W=0.2u L=0.06u
MNA1034 M SN N1_12 VPW NCH W=0.5u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.2u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.37u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.5u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.15u L=0.06u
MNOE022 NM NCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE026 NM BCLK_ NMUX VPW NCH W=0.15u L=0.06u
MP2 NET58 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.37u L=0.06u
MPA1020 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 NMUX D VDD VNW PCH W=0.5u L=0.06u
MPA1037 M SN VDD VNW PCH W=0.5u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.25u L=0.06u
MPA2 M NM VDD VNW PCH W=0.5u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.45u L=0.06u
MPOEN024 NM BCLK_ P1 VNW PCH W=0.15u L=0.06u
MPOEN028 NM NCLK_ NMUX VNW PCH W=0.45u L=0.06u
.ENDS	DFFNSQX1MA10TR

****
.SUBCKT DFFNSQX2MA10TR  VDD VSS VPW VNW Q   CKN D SN
MN2 NET50 NS NET47 VPW NCH W=0.2u L=0.06u
MN3 NET47 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET50 VPW NCH W=0.2u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.16u L=0.06u
MNA1018 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1030 NMUX D VSS VPW NCH W=0.3u L=0.06u
MNA1034 M SN N1_12 VPW NCH W=0.6u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.24u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.46u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.6u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.2u L=0.06u
MNOE022 NM NCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE026 NM BCLK_ NMUX VPW NCH W=0.2u L=0.06u
MP2 NET58 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.32u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.46u L=0.06u
MPA1020 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 NMUX D VDD VNW PCH W=0.7u L=0.06u
MPA1037 M SN VDD VNW PCH W=0.6u L=0.06u
MPA1042 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.3u L=0.06u
MPA2 M NM VDD VNW PCH W=0.6u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.6u L=0.06u
MPOEN024 NM BCLK_ P1 VNW PCH W=0.15u L=0.06u
MPOEN028 NM NCLK_ NMUX VNW PCH W=0.6u L=0.06u
.ENDS	DFFNSQX2MA10TR

****
.SUBCKT DFFNSQX3MA10TR  VDD VSS VPW VNW Q   CKN D SN
MN7 NET55 SN VSS VPW NCH W=0.2u L=0.06u
MN8 NET52 NS NET55 VPW NCH W=0.2u L=0.06u
MN9 S BCLK_ NET52 VPW NCH W=0.2u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.18u L=0.06u
MNA1015 NET0113 D VSS VPW NCH W=0.3u L=0.06u
MNA102 BCLK_ NCLK_ VSS VPW NCH W=0.28u L=0.06u
MNA1020 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1034 NS S VSS VPW NCH W=0.58u L=0.06u
MNA1038 M SN N1_12 VPW NCH W=0.6u L=0.06u
MNA106 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.6u L=0.06u
MNOE NM NCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE026 NM BCLK_ NET0113 VPW NCH W=0.25u L=0.06u
MNOE030 S NCLK_ M VPW NCH W=0.25u L=0.06u
MP5 NET66 NS VDD VNW PCH W=0.2u L=0.06u
MP8 S NCLK_ NET66 VNW PCH W=0.2u L=0.06u
MP9 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.36u L=0.06u
MPA1017 NET0113 D VDD VNW PCH W=0.7u L=0.06u
MPA1022 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1036 NS S VDD VNW PCH W=0.58u L=0.06u
MPA104 BCLK_ NCLK_ VDD VNW PCH W=0.34u L=0.06u
MPA1041 M SN VDD VNW PCH W=0.5u L=0.06u
MPA108 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA2 M NM VDD VNW PCH W=0.5u L=0.06u
MPOEN NM BCLK_ P1 VNW PCH W=0.15u L=0.06u
MPOEN028 NM NCLK_ NET0113 VNW PCH W=0.7u L=0.06u
MPOEN032 S BCLK_ M VNW PCH W=0.7u L=0.06u
.ENDS	DFFNSQX3MA10TR

****
.SUBCKT DFFNSRPQX1MA10TR  VDD VSS VPW VNW Q   CKN R D SN
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.3u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.3u L=0.06u
MN9 M R NET046 VPW NCH W=0.3u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.15u L=0.06u
MNA1027 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1039 NMUX D VSS VPW NCH W=0.2u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.2u L=0.06u
MNA1043 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.37u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.15u L=0.06u
MNOE031 NM NCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE035 NM BCLK_ NMUX VPW NCH W=0.15u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.45u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.45u L=0.06u
MP9 M SN VDD VNW PCH W=0.45u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.37u L=0.06u
MPA1029 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1041 NMUX D VDD VNW PCH W=0.5u L=0.06u
MPA1045 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.25u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.45u L=0.06u
MPOEN033 NM BCLK_ P1 VNW PCH W=0.15u L=0.06u
MPOEN037 NM NCLK_ NMUX VNW PCH W=0.45u L=0.06u
.ENDS	DFFNSRPQX1MA10TR

****
.SUBCKT DFFNSRPQX2MA10TR  VDD VSS VPW VNW Q   CKN R D SN
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.4u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.4u L=0.06u
MN9 M R NET046 VPW NCH W=0.4u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.21u L=0.06u
MNA1027 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1039 NMUX D VSS VPW NCH W=0.3u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.18u L=0.06u
MNA1043 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.47u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.2u L=0.06u
MNOE031 NM NCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE035 NM BCLK_ NMUX VPW NCH W=0.2u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.7u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.7u L=0.06u
MP9 M SN VDD VNW PCH W=0.7u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.47u L=0.06u
MPA1029 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1041 NMUX D VDD VNW PCH W=0.7u L=0.06u
MPA1045 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.36u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.6u L=0.06u
MPOEN033 NM BCLK_ P1 VNW PCH W=0.15u L=0.06u
MPOEN037 NM NCLK_ NMUX VNW PCH W=0.6u L=0.06u
.ENDS	DFFNSRPQX2MA10TR

****
.SUBCKT DFFNSRPQX3MA10TR  VDD VSS VPW VNW Q   CKN R D SN
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.4u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.4u L=0.06u
MN9 M R NET046 VPW NCH W=0.4u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.18u L=0.06u
MNA1026 NET0156 D VSS VPW NCH W=0.3u L=0.06u
MNA1031 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA104 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA1043 NS S VSS VPW NCH W=0.58u L=0.06u
MNA108 BCLK_ NCLK_ VSS VPW NCH W=0.28u L=0.06u
MNOE NM BCLK_ NET0156 VPW NCH W=0.25u L=0.06u
MNOE035 NM NCLK_ N1 VPW NCH W=0.15u L=0.06u
MNOE039 S NCLK_ M VPW NCH W=0.25u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.6u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.6u L=0.06u
MP9 M SN VDD VNW PCH W=0.6u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.36u L=0.06u
MPA1010 BCLK_ NCLK_ VDD VNW PCH W=0.34u L=0.06u
MPA1028 NET0156 D VDD VNW PCH W=0.7u L=0.06u
MPA1033 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1045 NS S VDD VNW PCH W=0.58u L=0.06u
MPA106 Q NS VDD VNW PCH W=2.1u L=0.06u
MPOEN NM NCLK_ NET0156 VNW PCH W=0.7u L=0.06u
MPOEN037 NM BCLK_ P1 VNW PCH W=0.15u L=0.06u
MPOEN041 S BCLK_ M VNW PCH W=0.7u L=0.06u
.ENDS	DFFNSRPQX3MA10TR

****
.SUBCKT DFFQNX0P5MA10TR  VDD VSS VPW VNW QN   CK D
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1010 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA1014 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1020 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1040 QN S VSS VPW NCH W=0.28u L=0.06u
MNA106 NS S VSS VPW NCH W=0.15u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE024 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NIN VPW NCH W=0.15u L=0.06u
MNOE032 S BCLK M VPW NCH W=0.15u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1012 NIN D VDD VNW PCH W=0.3u L=0.06u
MPA1016 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 M NM VDD VNW PCH W=0.25u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1042 QN S VDD VNW PCH W=0.37u L=0.06u
MPA108 NS S VDD VNW PCH W=0.15u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN026 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NIN VNW PCH W=0.15u L=0.06u
MPOEN034 S NCLK M VNW PCH W=0.15u L=0.06u
.ENDS	DFFQNX0P5MA10TR

****
.SUBCKT DFFQNX1MA10TR  VDD VSS VPW VNW QN   CK D
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1024 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.32u L=0.06u
MNA1036 QN S VSS VPW NCH W=0.53u L=0.06u
MNA1040 NET64 D VSS VPW NCH W=0.4u L=0.06u
MNA108 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE012 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE016 NM NCLK NET64 VPW NCH W=0.28u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.28u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1022 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1026 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.48u L=0.06u
MPA1038 QN S VDD VNW PCH W=0.7u L=0.06u
MPA104 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1042 NET64 D VDD VNW PCH W=0.4u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN014 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN018 NM BCLK NET64 VNW PCH W=0.28u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	DFFQNX1MA10TR

****
.SUBCKT DFFQNX2MA10TR  VDD VSS VPW VNW QN   CK D
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1028 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1036 QN S VSS VPW NCH W=1.06u L=0.06u
MNA1040 NET59 D VSS VPW NCH W=0.58u L=0.06u
MNA108 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE012 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE016 NM NCLK NET59 VPW NCH W=0.4u L=0.06u
MNOE020 S BCLK M VPW NCH W=0.4u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1026 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1030 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.6u L=0.06u
MPA1038 QN S VDD VNW PCH W=1.4u L=0.06u
MPA104 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1042 NET59 D VDD VNW PCH W=0.5u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN014 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN018 NM BCLK NET59 VNW PCH W=0.4u L=0.06u
MPOEN022 S NCLK M VNW PCH W=0.4u L=0.06u
.ENDS	DFFQNX2MA10TR

****
.SUBCKT DFFQNX3MA10TR  VDD VSS VPW VNW QN   CK D
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1028 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1036 QN S VSS VPW NCH W=1.62u L=0.06u
MNA1040 NET61 D VSS VPW NCH W=0.58u L=0.06u
MNA108 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE012 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE016 NM NCLK NET61 VPW NCH W=0.45u L=0.06u
MNOE020 S BCLK M VPW NCH W=0.58u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1026 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1030 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1038 QN S VDD VNW PCH W=2.1u L=0.06u
MPA104 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1042 NET61 D VDD VNW PCH W=0.5u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN014 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN018 NM BCLK NET61 VNW PCH W=0.45u L=0.06u
MPOEN022 S NCLK M VNW PCH W=0.58u L=0.06u
.ENDS	DFFQNX3MA10TR

****
.SUBCKT DFFQX0P5MA10TR  VDD VSS VPW VNW Q   CK D
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA1016 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.31u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE020 S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE036 NM NCLK NIN VPW NCH W=0.15u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.25u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.3u L=0.06u
MPA1018 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.22u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN022 S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN038 NM BCLK NIN VNW PCH W=0.15u L=0.06u
.ENDS	DFFQX0P5MA10TR

****
.SUBCKT DFFQX1MA10TR  VDD VSS VPW VNW Q   CK D
MNA1 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 NET88 D VSS VPW NCH W=0.4u L=0.06u
MNA1024 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.28u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA108 NS S VSS VPW NCH W=0.3u L=0.06u
MNOE S BCLK M VPW NCH W=0.28u L=0.06u
MNOE016 S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE036 NM NCLK NET88 VPW NCH W=0.28u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.48u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 NET88 D VDD VNW PCH W=0.4u L=0.06u
MPA1026 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.42u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPOEN S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN018 S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN038 NM BCLK NET88 VNW PCH W=0.28u L=0.06u
.ENDS	DFFQX1MA10TR

****
.SUBCKT DFFQX2MA10TR  VDD VSS VPW VNW Q   CK D
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 NET80 D VSS VPW NCH W=0.58u L=0.06u
MNA1024 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.4u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.46u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE016 S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE036 NM NCLK NET80 VPW NCH W=0.4u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 NET80 D VDD VNW PCH W=0.5u L=0.06u
MPA1026 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.6u L=0.06u
MPA1042 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN018 S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN038 NM BCLK NET80 VNW PCH W=0.4u L=0.06u
.ENDS	DFFQX2MA10TR

****
.SUBCKT DFFQX3MA10TR  VDD VSS VPW VNW Q   CK D
MNA1 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 NET85 D VSS VPW NCH W=0.58u L=0.06u
MNA1024 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.51u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA108 NS S VSS VPW NCH W=0.43u L=0.06u
MNOE S BCLK M VPW NCH W=0.45u L=0.06u
MNOE016 S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE036 NM NCLK NET85 VPW NCH W=0.45u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 NET85 D VDD VNW PCH W=0.5u L=0.06u
MPA1026 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.77u L=0.06u
MPA1042 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPOEN S NCLK M VNW PCH W=0.45u L=0.06u
MPOEN018 S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN038 NM BCLK NET85 VNW PCH W=0.45u L=0.06u
.ENDS	DFFQX3MA10TR

****
.SUBCKT DFFQX4MA10TR  VDD VSS VPW VNW Q   CK D
MNA1 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.15u L=0.06u
MNA1020 NET85 D VSS VPW NCH W=0.58u L=0.06u
MNA1024 N1_9 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.58u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1040 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA108 NS S VSS VPW NCH W=0.8u L=0.06u
MNOE S BCLK M VPW NCH W=0.58u L=0.06u
MNOE016 S NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_9 VPW NCH W=0.15u L=0.06u
MNOE036 NM NCLK NET85 VPW NCH W=0.45u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1010 NS S VDD VNW PCH W=1u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.15u L=0.06u
MPA1022 NET85 D VDD VNW PCH W=0.5u L=0.06u
MPA1026 P1_11 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1042 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPOEN S NCLK M VNW PCH W=0.58u L=0.06u
MPOEN018 S BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_11 VNW PCH W=0.15u L=0.06u
MPOEN038 NM BCLK NET85 VNW PCH W=0.45u L=0.06u
.ENDS	DFFQX4MA10TR

****
.SUBCKT DFFRPQNX0P5MA10TR  VDD VSS VPW VNW QN   CK R D
MN2 NET50 NET40 VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1010 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1020 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1034 QN S VSS VPW NCH W=0.28u L=0.06u
MNA1038 M NM VSS VPW NCH W=0.15u L=0.06u
MNA106 NET40 S VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.15u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NIN VPW NCH W=0.15u L=0.06u
MNOE030 S BCLK M VPW NCH W=0.15u L=0.06u
MP2 NET39 NET40 NET36 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET39 VNW PCH W=0.2u L=0.06u
MP5 NET36 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1012 NIN D VDD VNW PCH W=0.3u L=0.06u
MPA1022 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1036 QN S VDD VNW PCH W=0.37u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1041 M NM P1_12 VNW PCH W=0.45u L=0.06u
MPA108 NET40 S VDD VNW PCH W=0.15u L=0.06u
MPA2 P1_12 R VDD VNW PCH W=0.45u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN028 NM BCLK NIN VNW PCH W=0.15u L=0.06u
MPOEN032 S NCLK M VNW PCH W=0.15u L=0.06u
.ENDS	DFFRPQNX0P5MA10TR

****
.SUBCKT DFFRPQNX1MA10TR  VDD VSS VPW VNW QN   CK R D
MN2 NET53 NET37 VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET53 VPW NCH W=0.15u L=0.06u
MNA1 NET37 S VSS VPW NCH W=0.15u L=0.06u
MNA1022 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1026 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1030 QN S VSS VPW NCH W=0.53u L=0.06u
MNA1034 M R VSS VPW NCH W=0.32u L=0.06u
MNA1040 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA108 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA2 M NM VSS VPW NCH W=0.32u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE014 NM NCLK NIN VPW NCH W=0.28u L=0.06u
MNOE018 S BCLK M VPW NCH W=0.28u L=0.06u
MP2 NET36 NET37 NET39 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET36 VNW PCH W=0.2u L=0.06u
MP5 NET39 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NET37 S VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1024 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1028 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1032 QN S VDD VNW PCH W=0.7u L=0.06u
MPA1037 M R P1_12 VNW PCH W=0.68u L=0.06u
MPA1042 NIN D VDD VNW PCH W=0.4u L=0.06u
MPA2 P1_12 NM VDD VNW PCH W=0.68u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN016 NM BCLK NIN VNW PCH W=0.28u L=0.06u
MPOEN020 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	DFFRPQNX1MA10TR

****
.SUBCKT DFFRPQNX2MA10TR  VDD VSS VPW VNW QN   CK R D
MN2 NET53 NET37 VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET53 VPW NCH W=0.15u L=0.06u
MNA1 NET37 S VSS VPW NCH W=0.15u L=0.06u
MNA1022 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1026 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1030 QN S VSS VPW NCH W=1.16u L=0.06u
MNA1034 M R VSS VPW NCH W=0.4u L=0.06u
MNA1040 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA108 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA2 M NM VSS VPW NCH W=0.4u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE014 NM NCLK NIN VPW NCH W=0.4u L=0.06u
MNOE018 S BCLK M VPW NCH W=0.4u L=0.06u
MP2 NET36 NET37 NET39 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET36 VNW PCH W=0.2u L=0.06u
MP5 NET39 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NET37 S VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1024 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1028 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1032 QN S VDD VNW PCH W=1.4u L=0.06u
MPA1037 M R P1_12 VNW PCH W=0.8u L=0.06u
MPA1042 NIN D VDD VNW PCH W=0.6u L=0.06u
MPA2 P1_12 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN016 NM BCLK NIN VNW PCH W=0.4u L=0.06u
MPOEN020 S NCLK M VNW PCH W=0.4u L=0.06u
.ENDS	DFFRPQNX2MA10TR

****
.SUBCKT DFFRPQNX3MA10TR  VDD VSS VPW VNW QN   CK R D
MN2 NET53 NET37 VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET53 VPW NCH W=0.15u L=0.06u
MNA1 NET37 S VSS VPW NCH W=0.15u L=0.06u
MNA1022 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1026 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1030 QN S VSS VPW NCH W=1.74u L=0.06u
MNA1034 M R VSS VPW NCH W=0.4u L=0.06u
MNA1040 NET092 D VSS VPW NCH W=0.58u L=0.06u
MNA108 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA2 M NM VSS VPW NCH W=0.4u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE014 NM NCLK NET092 VPW NCH W=0.45u L=0.06u
MNOE018 S BCLK M VPW NCH W=0.5u L=0.06u
MP2 NET36 NET37 NET39 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET36 VNW PCH W=0.2u L=0.06u
MP5 NET39 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NET37 S VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1024 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1028 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1032 QN S VDD VNW PCH W=2.1u L=0.06u
MPA1037 M R P1_12 VNW PCH W=0.8u L=0.06u
MPA1042 NET092 D VDD VNW PCH W=0.5u L=0.06u
MPA2 P1_12 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN016 NM BCLK NET092 VNW PCH W=0.45u L=0.06u
MPOEN020 S NCLK M VNW PCH W=0.57u L=0.06u
.ENDS	DFFRPQNX3MA10TR

****
.SUBCKT DFFRPQX0P5MA10TR  VDD VSS VPW VNW Q   CK R D
MN2 NET63 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET63 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA1018 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1028 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.31u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.15u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE032 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE036 NM NCLK NIN VPW NCH W=0.15u L=0.06u
MP2 NET83 NS NET77 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET83 VNW PCH W=0.2u L=0.06u
MP5 NET77 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.22u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.3u L=0.06u
MPA1021 M NM P1 VNW PCH W=0.35u L=0.06u
MPA1030 P1_12 M VDD VNW PCH W=0.15u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA2 P1 R VDD VNW PCH W=0.35u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN034 NM NCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN038 NM BCLK NIN VNW PCH W=0.15u L=0.06u
.ENDS	DFFRPQX0P5MA10TR

****
.SUBCKT DFFRPQX1MA10TR  VDD VSS VPW VNW Q   CK R D
MN2 NET139 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET139 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1014 M R VSS VPW NCH W=0.28u L=0.06u
MNA1024 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 NET055 D VSS VPW NCH W=0.4u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA108 NS S VSS VPW NCH W=0.3u L=0.06u
MNA2 M NM VSS VPW NCH W=0.28u L=0.06u
MNOE S BCLK M VPW NCH W=0.28u L=0.06u
MNOE028 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE032 NM NCLK NET055 VPW NCH W=0.28u L=0.06u
MP2 NET129 NS NET123 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET129 VNW PCH W=0.2u L=0.06u
MP5 NET123 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.47u L=0.06u
MPA1017 M R P1 VNW PCH W=0.7u L=0.06u
MPA1026 P1_12 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NET055 D VDD VNW PCH W=0.4u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA2 P1 NM VDD VNW PCH W=0.7u L=0.06u
MPOEN S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN030 NM NCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN034 NM BCLK NET055 VNW PCH W=0.28u L=0.06u
.ENDS	DFFRPQX1MA10TR

****
.SUBCKT DFFRPQX2MA10TR  VDD VSS VPW VNW Q   CK R D
MN2 NET106 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET106 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1013 M R VSS VPW NCH W=0.4u L=0.06u
MNA1024 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 NET32 D VSS VPW NCH W=0.58u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.4u L=0.06u
MNA2 M NM VSS VPW NCH W=0.4u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE028 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE032 NM NCLK NET32 VPW NCH W=0.4u L=0.06u
MP2 NET102 NS NET96 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET102 VNW PCH W=0.2u L=0.06u
MP5 NET96 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.6u L=0.06u
MPA1016 M R P1 VNW PCH W=0.8u L=0.06u
MPA1026 P1_12 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NET32 D VDD VNW PCH W=0.5u L=0.06u
MPA1042 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA2 P1 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN030 NM NCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN034 NM BCLK NET32 VNW PCH W=0.4u L=0.06u
.ENDS	DFFRPQX2MA10TR

****
.SUBCKT DFFRPQX3MA10TR  VDD VSS VPW VNW Q   CK R D
MN2 NET140 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET140 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1010 M R VSS VPW NCH W=0.43u L=0.06u
MNA1020 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 NS S VSS VPW NCH W=0.53u L=0.06u
MNA1036 NET055 D VSS VPW NCH W=0.58u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA105 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA2 M NM VSS VPW NCH W=0.43u L=0.06u
MNOE S BCLK M VPW NCH W=0.45u L=0.06u
MNOE024 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NET055 VPW NCH W=0.45u L=0.06u
MP2 NET118 NS NET124 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET118 VNW PCH W=0.2u L=0.06u
MP5 NET124 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1013 M R P1 VNW PCH W=0.85u L=0.06u
MPA1022 P1_12 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 NS S VDD VNW PCH W=0.68u L=0.06u
MPA1038 NET055 D VDD VNW PCH W=0.5u L=0.06u
MPA1042 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA107 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA2 P1 NM VDD VNW PCH W=0.85u L=0.06u
MPOEN S NCLK M VNW PCH W=0.45u L=0.06u
MPOEN026 NM NCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NET055 VNW PCH W=0.45u L=0.06u
.ENDS	DFFRPQX3MA10TR

****
.SUBCKT DFFRPQX4MA10TR  VDD VSS VPW VNW Q   CK R D
MN2 NET134 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET134 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1014 M R VSS VPW NCH W=0.43u L=0.06u
MNA1024 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 NET056 D VSS VPW NCH W=0.58u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1040 Q NS VSS VPW NCH W=2.28u L=0.06u
MNA108 NS S VSS VPW NCH W=0.9u L=0.06u
MNA2 M NM VSS VPW NCH W=0.43u L=0.06u
MNOE S BCLK M VPW NCH W=0.55u L=0.06u
MNOE028 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE032 NM NCLK NET056 VPW NCH W=0.45u L=0.06u
MP2 NET124 NS NET118 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET124 VNW PCH W=0.2u L=0.06u
MP5 NET118 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.9u L=0.06u
MPA1017 M R P1 VNW PCH W=0.85u L=0.06u
MPA1026 P1_12 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NET056 D VDD VNW PCH W=0.5u L=0.06u
MPA1042 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPA2 P1 NM VDD VNW PCH W=0.85u L=0.06u
MPOEN S NCLK M VNW PCH W=0.55u L=0.06u
MPOEN030 NM NCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN034 NM BCLK NET056 VNW PCH W=0.45u L=0.06u
.ENDS	DFFRPQX4MA10TR

****
.SUBCKT DFFSQNX0P5MA10TR  VDD VSS VPW VNW QN   CK D SN
MN2 NET65 NS NET59 VPW NCH W=0.15u L=0.06u
MN3 NET59 SN VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET65 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1010 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1020 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1034 QN S VSS VPW NCH W=0.28u L=0.06u
MNA1038 M NM N1_12 VPW NCH W=0.3u L=0.06u
MNA106 NS S VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_12 SN VSS VPW NCH W=0.3u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NIN VPW NCH W=0.15u L=0.06u
MNOE030 S BCLK M VPW NCH W=0.15u L=0.06u
MP2 NET45 NS VDD VNW PCH W=0.15u L=0.06u
MP3 S BCLK NET45 VNW PCH W=0.15u L=0.06u
MP4 S SN VDD VNW PCH W=0.15u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1012 NIN D VDD VNW PCH W=0.3u L=0.06u
MPA1022 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1036 QN S VDD VNW PCH W=0.37u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1041 M NM VDD VNW PCH W=0.3u L=0.06u
MPA108 NS S VDD VNW PCH W=0.15u L=0.06u
MPA2 M SN VDD VNW PCH W=0.3u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN028 NM BCLK NIN VNW PCH W=0.15u L=0.06u
MPOEN032 S NCLK M VNW PCH W=0.15u L=0.06u
.ENDS	DFFSQNX0P5MA10TR

****
.SUBCKT DFFSQNX1MA10TR  VDD VSS VPW VNW QN   CK D SN
MN2 NET50 NS NET53 VPW NCH W=0.2u L=0.06u
MN3 NET53 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.2u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1026 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1030 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1034 QN S VSS VPW NCH W=0.53u L=0.06u
MNA1038 M SN N1_12 VPW NCH W=0.58u L=0.06u
MNA108 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.58u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE018 NM NCLK NIN VPW NCH W=0.28u L=0.06u
MNOE022 S BCLK M VPW NCH W=0.28u L=0.06u
MP2 NET42 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET42 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1010 NIN D VDD VNW PCH W=0.4u L=0.06u
MPA1014 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1028 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1032 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1036 QN S VDD VNW PCH W=0.7u L=0.06u
MPA1041 M SN VDD VNW PCH W=0.45u L=0.06u
MPA2 M NM VDD VNW PCH W=0.45u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN020 NM BCLK NIN VNW PCH W=0.28u L=0.06u
MPOEN024 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	DFFSQNX1MA10TR

****
.SUBCKT DFFSQNX2MA10TR  VDD VSS VPW VNW QN   CK D SN
MN2 NET50 NS NET53 VPW NCH W=0.2u L=0.06u
MN3 NET53 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.2u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1022 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1026 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1030 QN S VSS VPW NCH W=1.02u L=0.06u
MNA1034 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA1038 M SN N1_12 VPW NCH W=0.6u L=0.06u
MNA108 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.6u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE014 NM NCLK NIN VPW NCH W=0.4u L=0.06u
MNOE018 S BCLK M VPW NCH W=0.4u L=0.06u
MP2 NET42 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET42 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1024 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1028 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1032 QN S VDD VNW PCH W=1.4u L=0.06u
MPA1036 NIN D VDD VNW PCH W=0.5u L=0.06u
MPA1041 M SN VDD VNW PCH W=0.6u L=0.06u
MPA2 M NM VDD VNW PCH W=0.6u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN016 NM BCLK NIN VNW PCH W=0.4u L=0.06u
MPOEN020 S NCLK M VNW PCH W=0.39u L=0.06u
.ENDS	DFFSQNX2MA10TR

****
.SUBCKT DFFSQNX3MA10TR  VDD VSS VPW VNW QN   CK D SN
MN2 NET50 NS NET53 VPW NCH W=0.2u L=0.06u
MN3 NET53 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.2u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1026 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1030 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1034 QN S VSS VPW NCH W=1.59u L=0.06u
MNA1038 M SN N1_12 VPW NCH W=0.6u L=0.06u
MNA108 NET089 D VSS VPW NCH W=0.58u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.6u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE018 NM NCLK NET089 VPW NCH W=0.45u L=0.06u
MNOE022 S BCLK M VPW NCH W=0.54u L=0.06u
MP2 NET42 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET42 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1010 NET089 D VDD VNW PCH W=0.5u L=0.06u
MPA1014 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1028 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1032 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1036 QN S VDD VNW PCH W=2.1u L=0.06u
MPA1041 M SN VDD VNW PCH W=0.58u L=0.06u
MPA2 M NM VDD VNW PCH W=0.58u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN020 NM BCLK NET089 VNW PCH W=0.45u L=0.06u
MPOEN024 S NCLK M VNW PCH W=0.53u L=0.06u
.ENDS	DFFSQNX3MA10TR

****
.SUBCKT DFFSQX0P5MA10TR  VDD VSS VPW VNW Q   CK D SN
MN2 NET69 NS NET72 VPW NCH W=0.15u L=0.06u
MN3 NET72 SN VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET69 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA1022 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1034 M NM N1_12 VPW NCH W=0.25u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.31u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_12 SN VSS VPW NCH W=0.25u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE026 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE030 NM NCLK NIN VPW NCH W=0.15u L=0.06u
MP2 NET83 NS VDD VNW PCH W=0.15u L=0.06u
MP3 S BCLK NET83 VNW PCH W=0.15u L=0.06u
MP4 S SN VDD VNW PCH W=0.15u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.25u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.3u L=0.06u
MPA1024 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1037 M NM VDD VNW PCH W=0.25u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA2 M SN VDD VNW PCH W=0.25u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN028 NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN032 NM BCLK NIN VNW PCH W=0.15u L=0.06u
.ENDS	DFFSQX0P5MA10TR

****
.SUBCKT DFFSQX1MA10TR  VDD VSS VPW VNW Q   CK D SN
MN2 NET44 NS NET47 VPW NCH W=0.2u L=0.06u
MN3 NET47 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET44 VPW NCH W=0.2u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1018 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1030 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA1034 M SN N1_12 VPW NCH W=0.4u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA108 NS S VSS VPW NCH W=0.28u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.4u L=0.06u
MNOE S BCLK M VPW NCH W=0.28u L=0.06u
MNOE022 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NIN VPW NCH W=0.28u L=0.06u
MP2 NET58 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET58 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.52u L=0.06u
MPA1020 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 NIN D VDD VNW PCH W=0.4u L=0.06u
MPA1037 M SN VDD VNW PCH W=0.45u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA2 M NM VDD VNW PCH W=0.45u L=0.06u
MPOEN S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN024 NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN028 NM BCLK NIN VNW PCH W=0.28u L=0.06u
.ENDS	DFFSQX1MA10TR

****
.SUBCKT DFFSQX2MA10TR  VDD VSS VPW VNW Q   CK D SN
MN2 NET50 NS NET47 VPW NCH W=0.2u L=0.06u
MN3 NET47 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.2u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1018 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1030 NMUX D VSS VPW NCH W=0.58u L=0.06u
MNA1034 M SN N1_12 VPW NCH W=0.6u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.43u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.6u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE022 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MP2 NET58 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET58 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1020 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 NMUX D VDD VNW PCH W=0.5u L=0.06u
MPA1037 M SN VDD VNW PCH W=0.6u L=0.06u
MPA1042 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA2 M NM VDD VNW PCH W=0.6u L=0.06u
MPOEN S NCLK M VNW PCH W=0.39u L=0.06u
MPOEN024 NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN028 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
.ENDS	DFFSQX2MA10TR

****
.SUBCKT DFFSQX3MA10TR  VDD VSS VPW VNW Q   CK D SN
MN7 S NCLK NET49 VPW NCH W=0.2u L=0.06u
MN8 NET52 SN VSS VPW NCH W=0.2u L=0.06u
MN9 NET49 NS NET52 VPW NCH W=0.2u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1016 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA102 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA1030 NS S VSS VPW NCH W=0.45u L=0.06u
MNA1034 NET0105 D VSS VPW NCH W=0.58u L=0.06u
MNA1038 M SN N1_12 VPW NCH W=0.66u L=0.06u
MNA106 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.66u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE022 NM NCLK NET0105 VPW NCH W=0.45u L=0.06u
MNOE026 S BCLK M VPW NCH W=0.44u L=0.06u
MP7 NET66 NS VDD VNW PCH W=0.2u L=0.06u
MP8 S BCLK NET66 VNW PCH W=0.2u L=0.06u
MP9 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1018 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1036 NET0105 D VDD VNW PCH W=0.5u L=0.06u
MPA104 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1041 M SN VDD VNW PCH W=0.62u L=0.06u
MPA108 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA2 M NM VDD VNW PCH W=0.62u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN024 NM BCLK NET0105 VNW PCH W=0.45u L=0.06u
MPOEN028 S NCLK M VNW PCH W=0.44u L=0.06u
.ENDS	DFFSQX3MA10TR

****
.SUBCKT DFFSQX4MA10TR  VDD VSS VPW VNW Q   CK D SN
MN10 NET55 SN VSS VPW NCH W=0.2u L=0.06u
MN11 NET52 NS NET55 VPW NCH W=0.2u L=0.06u
MN12 S NCLK NET52 VPW NCH W=0.2u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1013 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1021 NET0105 D VSS VPW NCH W=0.58u L=0.06u
MNA1025 NS S VSS VPW NCH W=0.8u L=0.06u
MNA1029 M SN N1_12 VPW NCH W=0.66u L=0.06u
MNA103 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1035 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA2 N1_12 NM VSS VPW NCH W=0.66u L=0.06u
MNOE NM NCLK NET0105 VPW NCH W=0.45u L=0.06u
MNOE017 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE09 S BCLK M VPW NCH W=0.54u L=0.06u
MP10 NET66 NS VDD VNW PCH W=0.2u L=0.06u
MP11 S BCLK NET66 VNW PCH W=0.2u L=0.06u
MP12 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1015 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1023 NET0105 D VDD VNW PCH W=0.5u L=0.06u
MPA1027 NS S VDD VNW PCH W=1u L=0.06u
MPA1032 M SN VDD VNW PCH W=0.62u L=0.06u
MPA1037 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA105 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPA2 M NM VDD VNW PCH W=0.62u L=0.06u
MPOEN NM BCLK NET0105 VNW PCH W=0.45u L=0.06u
MPOEN011 S NCLK M VNW PCH W=0.53u L=0.06u
MPOEN019 NM NCLK P1 VNW PCH W=0.15u L=0.06u
.ENDS	DFFSQX4MA10TR

****
.SUBCKT DFFSRPQX0P5MA10TR  VDD VSS VPW VNW Q   CK R D SN
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.2u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.2u L=0.06u
MN9 M R NET046 VPW NCH W=0.2u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA1031 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1043 Q NS VSS VPW NCH W=0.31u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE035 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE039 NM NCLK NIN VPW NCH W=0.15u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.35u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.35u L=0.06u
MP9 M SN VDD VNW PCH W=0.35u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.25u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.3u L=0.06u
MPA1033 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1045 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.22u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN037 NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN041 NM BCLK NIN VNW PCH W=0.15u L=0.06u
.ENDS	DFFSRPQX0P5MA10TR

****
.SUBCKT DFFSRPQX1MA10TR  VDD VSS VPW VNW Q   CK R D SN
MN12 M NM NET79 VPW NCH W=0.32u L=0.06u
MN13 NET79 SN VSS VPW NCH W=0.32u L=0.06u
MN14 M R NET79 VPW NCH W=0.32u L=0.06u
MN15 S R NET64 VPW NCH W=0.2u L=0.06u
MN16 NET70 SN VSS VPW NCH W=0.2u L=0.06u
MN17 S NCLK NET61 VPW NCH W=0.2u L=0.06u
MN18 NET64 SN VSS VPW NCH W=0.2u L=0.06u
MN19 NET61 NS NET70 VPW NCH W=0.2u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1021 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1025 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA1029 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1037 NS S VSS VPW NCH W=0.28u L=0.06u
MNA1041 NIN D VSS VPW NCH W=0.4u L=0.06u
MNOE NM NCLK NIN VPW NCH W=0.28u L=0.06u
MNOE015 S BCLK M VPW NCH W=0.28u L=0.06u
MNOE033 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MP12 M NM NET108 VNW PCH W=0.6u L=0.06u
MP13 NET108 R VDD VNW PCH W=0.6u L=0.06u
MP14 M SN VDD VNW PCH W=0.6u L=0.06u
MP15 S BCLK NET99 VNW PCH W=0.2u L=0.06u
MP16 NET90 R VDD VNW PCH W=0.2u L=0.06u
MP17 S SN VDD VNW PCH W=0.2u L=0.06u
MP18 NET99 NS NET90 VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1023 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1027 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA1031 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1039 NS S VDD VNW PCH W=0.62u L=0.06u
MPA1043 NIN D VDD VNW PCH W=0.4u L=0.06u
MPOEN NM BCLK NIN VNW PCH W=0.28u L=0.06u
MPOEN017 S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN035 NM NCLK P1 VNW PCH W=0.15u L=0.06u
.ENDS	DFFSRPQX1MA10TR

****
.SUBCKT DFFSRPQX2MA10TR  VDD VSS VPW VNW Q   CK R D SN
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.4u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.4u L=0.06u
MN9 M R NET046 VPW NCH W=0.4u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1027 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1039 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1043 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.35u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE031 NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE035 NM NCLK NIN VPW NCH W=0.4u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.7u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.7u L=0.06u
MP9 M SN VDD VNW PCH W=0.7u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1029 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1041 NIN D VDD VNW PCH W=0.5u L=0.06u
MPA1045 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN033 NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN037 NM BCLK NIN VNW PCH W=0.4u L=0.06u
.ENDS	DFFSRPQX2MA10TR

****
.SUBCKT DFFSRPQX3MA10TR  VDD VSS VPW VNW Q   CK R D SN
MN15 S R NET67 VPW NCH W=0.2u L=0.06u
MN16 NET70 SN VSS VPW NCH W=0.2u L=0.06u
MN17 S NCLK NET79 VPW NCH W=0.2u L=0.06u
MN18 NET67 SN VSS VPW NCH W=0.2u L=0.06u
MN19 NET79 NS NET70 VPW NCH W=0.2u L=0.06u
MN20 M NM NET88 VPW NCH W=0.4u L=0.06u
MN21 NET88 SN VSS VPW NCH W=0.4u L=0.06u
MN22 M R NET88 VPW NCH W=0.4u L=0.06u
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1022 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1026 NS S VSS VPW NCH W=0.45u L=0.06u
MNA1030 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA1034 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1043 NET0155 D VSS VPW NCH W=0.58u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE014 NM NCLK NET0155 VPW NCH W=0.45u L=0.06u
MNOE018 S BCLK M VPW NCH W=0.4u L=0.06u
MP15 S BCLK NET96 VNW PCH W=0.2u L=0.06u
MP16 NET105 R VDD VNW PCH W=0.2u L=0.06u
MP17 S SN VDD VNW PCH W=0.2u L=0.06u
MP18 NET96 NS NET105 VNW PCH W=0.2u L=0.06u
MP19 M NM NET108 VNW PCH W=0.7u L=0.06u
MP20 NET108 R VDD VNW PCH W=0.7u L=0.06u
MP21 M SN VDD VNW PCH W=0.7u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1024 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA1028 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1032 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1036 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1045 NET0155 D VDD VNW PCH W=0.5u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN016 NM BCLK NET0155 VNW PCH W=0.45u L=0.06u
MPOEN020 S NCLK M VNW PCH W=0.4u L=0.06u
.ENDS	DFFSRPQX3MA10TR

****
.SUBCKT DFFSRPQX4MA10TR  VDD VSS VPW VNW Q   CK R D SN
MN12 S R NET73 VPW NCH W=0.2u L=0.06u
MN13 NET79 SN VSS VPW NCH W=0.2u L=0.06u
MN14 S NCLK NET70 VPW NCH W=0.2u L=0.06u
MN15 NET73 SN VSS VPW NCH W=0.2u L=0.06u
MN16 NET70 NS NET79 VPW NCH W=0.2u L=0.06u
MN17 M NM NET64 VPW NCH W=0.4u L=0.06u
MN18 NET64 SN VSS VPW NCH W=0.4u L=0.06u
MN19 M R NET64 VPW NCH W=0.4u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1014 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1019 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1033 NS S VSS VPW NCH W=0.8u L=0.06u
MNA1037 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA1041 NET0155 D VSS VPW NCH W=0.58u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE025 NM NCLK NET0155 VPW NCH W=0.45u L=0.06u
MNOE029 S BCLK M VPW NCH W=0.4u L=0.06u
MP12 S BCLK NET108 VNW PCH W=0.2u L=0.06u
MP13 NET99 R VDD VNW PCH W=0.2u L=0.06u
MP14 S SN VDD VNW PCH W=0.2u L=0.06u
MP15 NET108 NS NET99 VNW PCH W=0.2u L=0.06u
MP16 M NM NET96 VNW PCH W=0.7u L=0.06u
MP17 NET96 R VDD VNW PCH W=0.7u L=0.06u
MP18 M SN VDD VNW PCH W=0.7u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1016 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPA1021 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1035 NS S VDD VNW PCH W=1u L=0.06u
MPA1039 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA1043 NET0155 D VDD VNW PCH W=0.5u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN027 NM BCLK NET0155 VNW PCH W=0.45u L=0.06u
MPOEN031 S NCLK M VNW PCH W=0.4u L=0.06u
.ENDS	DFFSRPQX4MA10TR

****
.SUBCKT DFFYQX1MA10TR  VDD VSS VPW VNW Q   CK D
MNA1 NCLK CK VSS VPW NCH W=0.29u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.4u L=0.06u
MNA1020 N1_9 M VSS VPW NCH W=0.4u L=0.06u
MNA1028 M NM VSS VPW NCH W=0.32u L=0.06u
MNA1036 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1040 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.32u L=0.06u
MNOE S BCLK M VPW NCH W=0.28u L=0.06u
MNOE016 S NCLK N1 VPW NCH W=0.4u L=0.06u
MNOE024 NM BCLK N1_9 VPW NCH W=0.4u L=0.06u
MNOE032 NM NCLK NIN VPW NCH W=0.28u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.36u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.5u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.4u L=0.06u
MPA1022 P1_11 M VDD VNW PCH W=0.4u L=0.06u
MPA1030 M NM VDD VNW PCH W=0.5u L=0.06u
MPA1038 NIN D VDD VNW PCH W=0.4u L=0.06u
MPA1042 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPOEN S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN018 S BCLK P1 VNW PCH W=0.4u L=0.06u
MPOEN026 NM NCLK P1_11 VNW PCH W=0.4u L=0.06u
MPOEN034 NM BCLK NIN VNW PCH W=0.28u L=0.06u
.ENDS	DFFYQX1MA10TR

****
.SUBCKT DFFYQX2MA10TR  VDD VSS VPW VNW Q   CK D
MNA1 NCLK CK VSS VPW NCH W=0.42u L=0.06u
MNA1012 N1 NS VSS VPW NCH W=0.4u L=0.06u
MNA1020 N1_9 M VSS VPW NCH W=0.4u L=0.06u
MNA1028 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1036 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.35u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.53u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE016 S NCLK N1 VPW NCH W=0.4u L=0.06u
MNOE024 NM BCLK N1_9 VPW NCH W=0.4u L=0.06u
MNOE032 NM NCLK NIN VPW NCH W=0.4u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.52u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1014 P1 NS VDD VNW PCH W=0.4u L=0.06u
MPA1022 P1_11 M VDD VNW PCH W=0.4u L=0.06u
MPA1030 M NM VDD VNW PCH W=0.6u L=0.06u
MPA1038 NIN D VDD VNW PCH W=0.5u L=0.06u
MPA1042 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.7u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN018 S BCLK P1 VNW PCH W=0.4u L=0.06u
MPOEN026 NM NCLK P1_11 VNW PCH W=0.4u L=0.06u
MPOEN034 NM BCLK NIN VNW PCH W=0.4u L=0.06u
.ENDS	DFFYQX2MA10TR

****
.SUBCKT DFFYQX3MA10TR  VDD VSS VPW VNW Q   CK D
MNA1 N1 NS VSS VPW NCH W=0.4u L=0.06u
MNA1024 NS S VSS VPW NCH W=0.4u L=0.06u
MNA1028 NCLK CK VSS VPW NCH W=0.3u L=0.06u
MNA1032 BCLK NCLK VSS VPW NCH W=0.26u L=0.06u
MNA1036 M NM VSS VPW NCH W=0.38u L=0.06u
MNA104 NET85 D VSS VPW NCH W=0.58u L=0.06u
MNA1040 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA108 N1_9 M VSS VPW NCH W=0.4u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.4u L=0.06u
MNOE012 NM BCLK N1_9 VPW NCH W=0.4u L=0.06u
MNOE016 NM NCLK NET85 VPW NCH W=0.45u L=0.06u
MNOE020 S BCLK M VPW NCH W=0.45u L=0.06u
MPA1 P1 NS VDD VNW PCH W=0.4u L=0.06u
MPA1010 P1_11 M VDD VNW PCH W=0.4u L=0.06u
MPA1026 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1030 NCLK CK VDD VNW PCH W=0.37u L=0.06u
MPA1034 BCLK NCLK VDD VNW PCH W=0.52u L=0.06u
MPA1038 M NM VDD VNW PCH W=0.76u L=0.06u
MPA1042 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA106 NET85 D VDD VNW PCH W=0.5u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.4u L=0.06u
MPOEN014 NM NCLK P1_11 VNW PCH W=0.4u L=0.06u
MPOEN018 NM BCLK NET85 VNW PCH W=0.45u L=0.06u
MPOEN022 S NCLK M VNW PCH W=0.45u L=0.06u
.ENDS	DFFYQX3MA10TR

****
.SUBCKT DFFYQX4MA10TR  VDD VSS VPW VNW Q   CK D
MNA1 N1 NS VSS VPW NCH W=0.4u L=0.06u
MNA1020 NS S VSS VPW NCH W=1.05u L=0.06u
MNA1024 NCLK CK VSS VPW NCH W=0.38u L=0.06u
MNA1028 BCLK NCLK VSS VPW NCH W=0.35u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.45u L=0.06u
MNA1036 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA104 N1_9 M VSS VPW NCH W=0.4u L=0.06u
MNA1040 NET85 D VSS VPW NCH W=0.58u L=0.06u
MNOE S NCLK N1 VPW NCH W=0.4u L=0.06u
MNOE012 NM NCLK NET85 VPW NCH W=0.45u L=0.06u
MNOE016 S BCLK M VPW NCH W=0.57u L=0.06u
MNOE08 NM BCLK N1_9 VPW NCH W=0.4u L=0.06u
MPA1 P1 NS VDD VNW PCH W=0.4u L=0.06u
MPA1022 NS S VDD VNW PCH W=1.25u L=0.06u
MPA1026 NCLK CK VDD VNW PCH W=0.47u L=0.06u
MPA1030 BCLK NCLK VDD VNW PCH W=0.7u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1038 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA1042 NET85 D VDD VNW PCH W=0.5u L=0.06u
MPA106 P1_11 M VDD VNW PCH W=0.4u L=0.06u
MPOEN S BCLK P1 VNW PCH W=0.4u L=0.06u
MPOEN010 NM NCLK P1_11 VNW PCH W=0.4u L=0.06u
MPOEN014 NM BCLK NET85 VNW PCH W=0.45u L=0.06u
MPOEN018 S NCLK M VNW PCH W=0.57u L=0.06u
.ENDS	DFFYQX4MA10TR

****
.SUBCKT DLY2X0P5MA10TR  VDD VSS VPW VNW Y   A
MN0 VSS NET15 VSS VPW NCH W=0.18u L=0.06u
MNA1 Y NET15 VSS VPW NCH W=0.265u L=0.06u
MNA104 N1 A VSS VPW NCH W=0.15u L=0.06u
MNOE NET15 A N1 VPW NCH W=0.15u L=0.06u
MP0 VDD NET15 VDD VNW PCH W=0.22u L=0.06u
MPA1 Y NET15 VDD VNW PCH W=0.35u L=0.06u
MPA106 P1 A VDD VNW PCH W=0.22u L=0.06u
MPOEN NET15 A P1 VNW PCH W=0.22u L=0.06u
.ENDS	DLY2X0P5MA10TR

****
.SUBCKT DLY4X0P5MA10TR  VDD VSS VPW VNW Y   A
MN0 VSS NBIN VSS VPW NCH W=0.185u L=0.06u
MNA1 N1 BIN VSS VPW NCH W=0.15u L=0.06u
MNA1010 N1_5 A VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_9 NIN VSS VPW NCH W=0.15u L=0.06u
MNA106 Y NBIN VSS VPW NCH W=0.265u L=0.06u
MNOE NBIN BIN N1 VPW NCH W=0.15u L=0.06u
MNOE014 NIN A N1_5 VPW NCH W=0.15u L=0.06u
MNOE022 BIN NIN N1_9 VPW NCH W=0.15u L=0.06u
MP0 VDD NBIN VDD VNW PCH W=0.22u L=0.06u
MPA1 P1 BIN VDD VNW PCH W=0.22u L=0.06u
MPA1012 P1_7 A VDD VNW PCH W=0.22u L=0.06u
MPA1020 P1_11 NIN VDD VNW PCH W=0.22u L=0.06u
MPA108 Y NBIN VDD VNW PCH W=0.35u L=0.06u
MPOEN NBIN BIN P1 VNW PCH W=0.22u L=0.06u
MPOEN016 NIN A P1_7 VNW PCH W=0.22u L=0.06u
MPOEN024 BIN NIN P1_11 VNW PCH W=0.22u L=0.06u
.ENDS	DLY4X0P5MA10TR

****
.SUBCKT EDFFQNX0P5MA10TR  VDD VSS VPW VNW QN   CK E D
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 NEN E VSS VPW NCH W=0.2u L=0.06u
MNA1016 NFB NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1024 NET59 D VSS VPW NCH W=0.25u L=0.06u
MNA1032 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1036 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 N1_13 NS VSS VPW NCH W=0.15u L=0.06u
MNA1048 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1052 QN S VSS VPW NCH W=0.28u L=0.06u
MNA1060 NET75 NFB VSS VPW NCH W=0.25u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE020 NENMUX E NET59 VPW NCH W=0.25u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.15u L=0.06u
MNOE044 S NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE056 NENMUX NEN NET75 VPW NCH W=0.25u L=0.06u
MNOE08 NM NCLK NENMUX VPW NCH W=0.15u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 NEN E VDD VNW PCH W=0.27u L=0.06u
MPA1018 NFB NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 NET59 D VDD VNW PCH W=0.3u L=0.06u
MPA1034 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1038 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA104 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1042 P1_15 NS VDD VNW PCH W=0.15u L=0.06u
MPA1050 M NM VDD VNW PCH W=0.2u L=0.06u
MPA1054 QN S VDD VNW PCH W=0.37u L=0.06u
MPA1062 NET75 NFB VDD VNW PCH W=0.3u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 NM BCLK NENMUX VNW PCH W=0.15u L=0.06u
MPOEN022 NENMUX NEN NET59 VNW PCH W=0.25u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN046 S BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN058 NENMUX E NET75 VNW PCH W=0.25u L=0.06u
.ENDS	EDFFQNX0P5MA10TR

****
.SUBCKT EDFFQNX1MA10TR  VDD VSS VPW VNW QN   CK E D
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 NEN E VSS VPW NCH W=0.27u L=0.06u
MNA1016 FB NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1024 NIN D VSS VPW NCH W=0.28u L=0.06u
MNA1032 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1036 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1040 N1_13 NS VSS VPW NCH W=0.15u L=0.06u
MNA1048 M NM VSS VPW NCH W=0.32u L=0.06u
MNA1052 QN S VSS VPW NCH W=0.53u L=0.06u
MNA1060 NFB FB VSS VPW NCH W=0.28u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE020 NENMUX E NIN VPW NCH W=0.28u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.28u L=0.06u
MNOE044 S NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE056 NENMUX NEN NFB VPW NCH W=0.28u L=0.06u
MNOE08 NM NCLK NENMUX VPW NCH W=0.28u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 NEN E VDD VNW PCH W=0.36u L=0.06u
MPA1018 FB NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 NIN D VDD VNW PCH W=0.36u L=0.06u
MPA1034 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1038 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA104 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1042 P1_15 NS VDD VNW PCH W=0.15u L=0.06u
MPA1050 M NM VDD VNW PCH W=0.48u L=0.06u
MPA1054 QN S VDD VNW PCH W=0.7u L=0.06u
MPA1062 NFB FB VDD VNW PCH W=0.36u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 NM BCLK NENMUX VNW PCH W=0.28u L=0.06u
MPOEN022 NENMUX NEN NIN VNW PCH W=0.28u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN046 S BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN058 NENMUX E NFB VNW PCH W=0.28u L=0.06u
.ENDS	EDFFQNX1MA10TR

****
.SUBCKT EDFFQNX2MA10TR  VDD VSS VPW VNW QN   CK E D
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 NEN E VSS VPW NCH W=0.32u L=0.06u
MNA1016 FB NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1024 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA1032 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1036 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1040 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1044 N1_13 NS VSS VPW NCH W=0.15u L=0.06u
MNA1052 QN S VSS VPW NCH W=1.06u L=0.06u
MNA1060 NFB FB VSS VPW NCH W=0.4u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE020 NENMUX E NIN VPW NCH W=0.4u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.4u L=0.06u
MNOE048 S NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE056 NENMUX NEN NFB VPW NCH W=0.4u L=0.06u
MNOE08 NM NCLK NENMUX VPW NCH W=0.4u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 NEN E VDD VNW PCH W=0.43u L=0.06u
MPA1018 FB NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 NIN D VDD VNW PCH W=0.52u L=0.06u
MPA1034 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1038 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA104 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1042 M NM VDD VNW PCH W=0.6u L=0.06u
MPA1046 P1_15 NS VDD VNW PCH W=0.15u L=0.06u
MPA1054 QN S VDD VNW PCH W=1.4u L=0.06u
MPA1062 NFB FB VDD VNW PCH W=0.52u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 NM BCLK NENMUX VNW PCH W=0.4u L=0.06u
MPOEN022 NENMUX NEN NIN VNW PCH W=0.4u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN050 S BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN058 NENMUX E NFB VNW PCH W=0.4u L=0.06u
.ENDS	EDFFQNX2MA10TR

****
.SUBCKT EDFFQNX3MA10TR  VDD VSS VPW VNW QN   CK E D
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 NEN E VSS VPW NCH W=0.32u L=0.06u
MNA1016 FB NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1024 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1036 N1_13 NS VSS VPW NCH W=0.15u L=0.06u
MNA1044 QN S VSS VPW NCH W=1.59u L=0.06u
MNA1052 NFB FB VSS VPW NCH W=0.4u L=0.06u
MNA1056 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1060 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE020 NENMUX E NIN VPW NCH W=0.4u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.4u L=0.06u
MNOE040 S NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE048 NENMUX NEN NFB VPW NCH W=0.4u L=0.06u
MNOE08 NM NCLK NENMUX VPW NCH W=0.45u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 NEN E VDD VNW PCH W=0.43u L=0.06u
MPA1018 FB NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 NIN D VDD VNW PCH W=0.6u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1038 P1_15 NS VDD VNW PCH W=0.15u L=0.06u
MPA104 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1046 QN S VDD VNW PCH W=2.1u L=0.06u
MPA1054 NFB FB VDD VNW PCH W=0.6u L=0.06u
MPA1058 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1062 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 NM BCLK NENMUX VNW PCH W=0.45u L=0.06u
MPOEN022 NENMUX NEN NIN VNW PCH W=0.4u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.58u L=0.06u
MPOEN042 S BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN050 NENMUX E NFB VNW PCH W=0.4u L=0.06u
.ENDS	EDFFQNX3MA10TR

****
.SUBCKT EDFFQX0P5MA10TR  VDD VSS VPW VNW Q   CK E D
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA1012 NEN E VSS VPW NCH W=0.2u L=0.06u
MNA1016 NFB S VSS VPW NCH W=0.2u L=0.06u
MNA102 N1 NM VSS VPW NCH W=0.15u L=0.06u
MNA1024 NET0128 D VSS VPW NCH W=0.2u L=0.06u
MNA1032 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1036 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 NM M VSS VPW NCH W=0.15u L=0.06u
MNA1044 N1_13 S VSS VPW NCH W=0.15u L=0.06u
MNA1052 NET144 NENMUX VSS VPW NCH W=0.2u L=0.06u
MNA1056 Q NS VSS VPW NCH W=0.28u L=0.06u
MNOE M BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE020 NENMUX E NET0128 VPW NCH W=0.2u L=0.06u
MNOE028 NS BCLK NM VPW NCH W=0.15u L=0.06u
MNOE048 NS NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE060 NENMUX NEN NFB VPW NCH W=0.2u L=0.06u
MNOE08 M NCLK NET144 VPW NCH W=0.15u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1014 NEN E VDD VNW PCH W=0.27u L=0.06u
MPA1018 NFB S VDD VNW PCH W=0.3u L=0.06u
MPA1026 NET0128 D VDD VNW PCH W=0.4u L=0.06u
MPA1034 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1038 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA104 P1 NM VDD VNW PCH W=0.15u L=0.06u
MPA1042 NM M VDD VNW PCH W=0.2u L=0.06u
MPA1046 P1_15 S VDD VNW PCH W=0.15u L=0.06u
MPA1054 NET144 NENMUX VDD VNW PCH W=0.2u L=0.06u
MPA1058 Q NS VDD VNW PCH W=0.37u L=0.06u
MPOEN M NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 M BCLK NET144 VNW PCH W=0.15u L=0.06u
MPOEN022 NENMUX NEN NET0128 VNW PCH W=0.3u L=0.06u
MPOEN030 NS NCLK NM VNW PCH W=0.15u L=0.06u
MPOEN050 NS BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN062 NENMUX E NFB VNW PCH W=0.3u L=0.06u
.ENDS	EDFFQX0P5MA10TR

****
.SUBCKT EDFFQX1MA10TR  VDD VSS VPW VNW Q   CK E D
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA1012 NFB S VSS VPW NCH W=0.2u L=0.06u
MNA102 N1 NM VSS VPW NCH W=0.15u L=0.06u
MNA1024 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1028 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1032 NM M VSS VPW NCH W=0.32u L=0.06u
MNA1036 N1_13 S VSS VPW NCH W=0.15u L=0.06u
MNA1044 NET144 NENMUX VSS VPW NCH W=0.28u L=0.06u
MNA1048 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA1056 NIN D VSS VPW NCH W=0.2u L=0.06u
MNA1060 NEN E VSS VPW NCH W=0.26u L=0.06u
MNOE M BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE016 NENMUX NEN NFB VPW NCH W=0.2u L=0.06u
MNOE020 NS BCLK NM VPW NCH W=0.28u L=0.06u
MNOE040 NS NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE052 NENMUX E NIN VPW NCH W=0.2u L=0.06u
MNOE08 M NCLK NET144 VPW NCH W=0.28u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1014 NFB S VDD VNW PCH W=0.4u L=0.06u
MPA1026 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1030 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1034 NM M VDD VNW PCH W=0.48u L=0.06u
MPA1038 P1_15 S VDD VNW PCH W=0.15u L=0.06u
MPA104 P1 NM VDD VNW PCH W=0.15u L=0.06u
MPA1046 NET144 NENMUX VDD VNW PCH W=0.28u L=0.06u
MPA1050 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA1058 NIN D VDD VNW PCH W=0.4u L=0.06u
MPA1062 NEN E VDD VNW PCH W=0.34u L=0.06u
MPOEN M NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 M BCLK NET144 VNW PCH W=0.28u L=0.06u
MPOEN018 NENMUX E NFB VNW PCH W=0.3u L=0.06u
MPOEN022 NS NCLK NM VNW PCH W=0.28u L=0.06u
MPOEN042 NS BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN054 NENMUX NEN NIN VNW PCH W=0.3u L=0.06u
.ENDS	EDFFQX1MA10TR

****
.SUBCKT EDFFQX2MA10TR  VDD VSS VPW VNW Q   CK E D
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA1012 NEN E VSS VPW NCH W=0.31u L=0.06u
MNA1016 NFB S VSS VPW NCH W=0.3u L=0.06u
MNA102 N1 NM VSS VPW NCH W=0.15u L=0.06u
MNA1024 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA1032 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1036 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1040 NM M VSS VPW NCH W=0.4u L=0.06u
MNA1044 N1_13 S VSS VPW NCH W=0.15u L=0.06u
MNA1052 MUX NENMUX VSS VPW NCH W=0.4u L=0.06u
MNA1056 Q NS VSS VPW NCH W=1.06u L=0.06u
MNOE M BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE020 NENMUX E NIN VPW NCH W=0.3u L=0.06u
MNOE028 NS BCLK NM VPW NCH W=0.4u L=0.06u
MNOE048 NS NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE060 NENMUX NEN NFB VPW NCH W=0.3u L=0.06u
MNOE08 M NCLK MUX VPW NCH W=0.4u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1014 NEN E VDD VNW PCH W=0.41u L=0.06u
MPA1018 NFB S VDD VNW PCH W=0.5u L=0.06u
MPA1026 NIN D VDD VNW PCH W=0.5u L=0.06u
MPA1034 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1038 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA104 P1 NM VDD VNW PCH W=0.15u L=0.06u
MPA1042 NM M VDD VNW PCH W=0.6u L=0.06u
MPA1046 P1_15 S VDD VNW PCH W=0.15u L=0.06u
MPA1054 MUX NENMUX VDD VNW PCH W=0.4u L=0.06u
MPA1058 Q NS VDD VNW PCH W=1.4u L=0.06u
MPOEN M NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 M BCLK MUX VNW PCH W=0.4u L=0.06u
MPOEN022 NENMUX NEN NIN VNW PCH W=0.45u L=0.06u
MPOEN030 NS NCLK NM VNW PCH W=0.4u L=0.06u
MPOEN050 NS BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN062 NENMUX E NFB VNW PCH W=0.45u L=0.06u
.ENDS	EDFFQX2MA10TR

****
.SUBCKT EDFFQX3MA10TR  VDD VSS VPW VNW Q   CK E D
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA1012 NEN E VSS VPW NCH W=0.31u L=0.06u
MNA102 N1 NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NFB S VSS VPW NCH W=0.3u L=0.06u
MNA1028 NIN D VSS VPW NCH W=0.3u L=0.06u
MNA1032 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1036 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1040 N1_13 S VSS VPW NCH W=0.15u L=0.06u
MNA1048 MUX NENMUX VSS VPW NCH W=0.45u L=0.06u
MNA1056 Q NS VSS VPW NCH W=1.65u L=0.06u
MNA1060 NM M VSS VPW NCH W=0.58u L=0.06u
MNOE M BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE016 NS BCLK NM VPW NCH W=0.4u L=0.06u
MNOE024 NENMUX E NIN VPW NCH W=0.3u L=0.06u
MNOE044 NS NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE052 NENMUX NEN NFB VPW NCH W=0.3u L=0.06u
MNOE08 M NCLK MUX VPW NCH W=0.45u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1014 NEN E VDD VNW PCH W=0.41u L=0.06u
MPA1022 NFB S VDD VNW PCH W=0.6u L=0.06u
MPA1030 NIN D VDD VNW PCH W=0.6u L=0.06u
MPA1034 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1038 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA104 P1 NM VDD VNW PCH W=0.15u L=0.06u
MPA1042 P1_15 S VDD VNW PCH W=0.15u L=0.06u
MPA1050 MUX NENMUX VDD VNW PCH W=0.45u L=0.06u
MPA1058 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1062 NM M VDD VNW PCH W=0.7u L=0.06u
MPOEN M NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 M BCLK MUX VNW PCH W=0.45u L=0.06u
MPOEN018 NS NCLK NM VNW PCH W=0.58u L=0.06u
MPOEN026 NENMUX NEN NIN VNW PCH W=0.45u L=0.06u
MPOEN046 NS BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN054 NENMUX E NFB VNW PCH W=0.45u L=0.06u
.ENDS	EDFFQX3MA10TR

****
.SUBCKT ESDFFQNX0P5MA10TR  VDD VSS VPW VNW QN   CK E D SE SI
MNA1 S NS VSS VPW NCH W=0.17u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1024 NFB S VSS VPW NCH W=0.2u L=0.06u
MNA1032 NET0135 D VSS VPW NCH W=0.2u L=0.06u
MNA1040 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1044 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1048 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1052 NM M VSS VPW NCH W=0.15u L=0.06u
MNA1056 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET144 NSEMUX VSS VPW NCH W=0.15u L=0.06u
MNA1068 QN S VSS VPW NCH W=0.31u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.15u L=0.06u
MNOE028 NENMUX E NET0135 VPW NCH W=0.2u L=0.06u
MNOE036 NS BCLK NM VPW NCH W=0.15u L=0.06u
MNOE060 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE072 NSEMUX NSE NENMUX VPW NCH W=0.2u L=0.06u
MNOE076 NENMUX NEN NFB VPW NCH W=0.2u L=0.06u
MPA1 S NS VDD VNW PCH W=0.34u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NEN E VDD VNW PCH W=0.2u L=0.06u
MPA1026 NFB S VDD VNW PCH W=0.3u L=0.06u
MPA1034 NET0135 D VDD VNW PCH W=0.4u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1046 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1050 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1054 NM M VDD VNW PCH W=0.22u L=0.06u
MPA1058 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1066 NET144 NSEMUX VDD VNW PCH W=0.15u L=0.06u
MPA1070 QN S VDD VNW PCH W=0.37u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.15u L=0.06u
MPOEN030 NENMUX NEN NET0135 VNW PCH W=0.25u L=0.06u
MPOEN038 NS NCLK NM VNW PCH W=0.15u L=0.06u
MPOEN062 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN074 NSEMUX SE NENMUX VNW PCH W=0.25u L=0.06u
MPOEN078 NENMUX E NFB VNW PCH W=0.25u L=0.06u
.ENDS	ESDFFQNX0P5MA10TR

****
.SUBCKT ESDFFQNX1MA10TR  VDD VSS VPW VNW QN   CK E D SE SI
MNA1 S NS VSS VPW NCH W=0.27u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.26u L=0.06u
MNA1024 NFB S VSS VPW NCH W=0.2u L=0.06u
MNA1032 NET0135 D VSS VPW NCH W=0.2u L=0.06u
MNA1040 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1044 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1048 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1052 NM M VSS VPW NCH W=0.32u L=0.06u
MNA1056 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET144 NSEMUX VSS VPW NCH W=0.32u L=0.06u
MNA1068 QN S VSS VPW NCH W=0.58u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.28u L=0.06u
MNOE028 NENMUX E NET0135 VPW NCH W=0.2u L=0.06u
MNOE036 NS BCLK NM VPW NCH W=0.28u L=0.06u
MNOE060 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE072 NSEMUX NSE NENMUX VPW NCH W=0.2u L=0.06u
MNOE076 NENMUX NEN NFB VPW NCH W=0.2u L=0.06u
MPA1 S NS VDD VNW PCH W=0.54u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NEN E VDD VNW PCH W=0.34u L=0.06u
MPA1026 NFB S VDD VNW PCH W=0.4u L=0.06u
MPA1034 NET0135 D VDD VNW PCH W=0.4u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1046 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1050 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1054 NM M VDD VNW PCH W=0.48u L=0.06u
MPA1058 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1066 NET144 NSEMUX VDD VNW PCH W=0.32u L=0.06u
MPA1070 QN S VDD VNW PCH W=0.7u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.28u L=0.06u
MPOEN030 NENMUX NEN NET0135 VNW PCH W=0.3u L=0.06u
MPOEN038 NS NCLK NM VNW PCH W=0.28u L=0.06u
MPOEN062 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN074 NSEMUX SE NENMUX VNW PCH W=0.3u L=0.06u
MPOEN078 NENMUX E NFB VNW PCH W=0.3u L=0.06u
.ENDS	ESDFFQNX1MA10TR

****
.SUBCKT ESDFFQNX2MA10TR  VDD VSS VPW VNW QN   CK E D SE SI
MNA1 S NS VSS VPW NCH W=0.3u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.31u L=0.06u
MNA1024 NFB S VSS VPW NCH W=0.3u L=0.06u
MNA1032 NET0135 D VSS VPW NCH W=0.3u L=0.06u
MNA1040 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1044 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1048 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1052 NM M VSS VPW NCH W=0.4u L=0.06u
MNA1056 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET144 NSEMUX VSS VPW NCH W=0.4u L=0.06u
MNA1068 QN S VSS VPW NCH W=1.06u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.4u L=0.06u
MNOE028 NENMUX E NET0135 VPW NCH W=0.3u L=0.06u
MNOE036 NS BCLK NM VPW NCH W=0.4u L=0.06u
MNOE060 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE072 NSEMUX NSE NENMUX VPW NCH W=0.3u L=0.06u
MNOE076 NENMUX NEN NFB VPW NCH W=0.3u L=0.06u
MPA1 S NS VDD VNW PCH W=0.7u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NEN E VDD VNW PCH W=0.41u L=0.06u
MPA1026 NFB S VDD VNW PCH W=0.6u L=0.06u
MPA1034 NET0135 D VDD VNW PCH W=0.6u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1046 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1050 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1054 NM M VDD VNW PCH W=0.65u L=0.06u
MPA1058 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1066 NET144 NSEMUX VDD VNW PCH W=0.4u L=0.06u
MPA1070 QN S VDD VNW PCH W=1.4u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.4u L=0.06u
MPOEN030 NENMUX NEN NET0135 VNW PCH W=0.45u L=0.06u
MPOEN038 NS NCLK NM VNW PCH W=0.4u L=0.06u
MPOEN062 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN074 NSEMUX SE NENMUX VNW PCH W=0.45u L=0.06u
MPOEN078 NENMUX E NFB VNW PCH W=0.45u L=0.06u
.ENDS	ESDFFQNX2MA10TR

****
.SUBCKT ESDFFQNX3MA10TR  VDD VSS VPW VNW QN   CK E D SE SI
MNA1 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1012 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNA1028 NEN E VSS VPW NCH W=0.31u L=0.06u
MNA1032 NFB S VSS VPW NCH W=0.3u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1040 NET0135 D VSS VPW NCH W=0.3u L=0.06u
MNA1044 NM M VSS VPW NCH W=0.51u L=0.06u
MNA1052 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1056 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET144 NSEMUX VSS VPW NCH W=0.45u L=0.06u
MNA1076 QN S VSS VPW NCH W=1.74u L=0.06u
MNA108 S NS VSS VPW NCH W=0.43u L=0.06u
MNOE NS BCLK NM VPW NCH W=0.4u L=0.06u
MNOE016 NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE024 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE036 NENMUX E NET0135 VPW NCH W=0.3u L=0.06u
MNOE048 M NCLK NET144 VPW NCH W=0.45u L=0.06u
MNOE060 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE068 NSEMUX NSE NENMUX VPW NCH W=0.3u L=0.06u
MNOE072 NENMUX NEN NFB VPW NCH W=0.3u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1010 S NS VDD VNW PCH W=0.7u L=0.06u
MPA1014 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1022 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1030 NEN E VDD VNW PCH W=0.41u L=0.06u
MPA1034 NFB S VDD VNW PCH W=0.6u L=0.06u
MPA1042 NET0135 D VDD VNW PCH W=0.6u L=0.06u
MPA1046 NM M VDD VNW PCH W=0.77u L=0.06u
MPA1054 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1058 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA1066 NET144 NSEMUX VDD VNW PCH W=0.45u L=0.06u
MPA1078 QN S VDD VNW PCH W=2.1u L=0.06u
MPOEN NS NCLK NM VNW PCH W=0.45u L=0.06u
MPOEN018 NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN026 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN038 NENMUX NEN NET0135 VNW PCH W=0.45u L=0.06u
MPOEN050 M BCLK NET144 VNW PCH W=0.45u L=0.06u
MPOEN062 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN070 NSEMUX SE NENMUX VNW PCH W=0.45u L=0.06u
MPOEN074 NENMUX E NFB VNW PCH W=0.45u L=0.06u
.ENDS	ESDFFQNX3MA10TR

****
.SUBCKT ESDFFQX0P5MA10TR  VDD VSS VPW VNW Q   CK E D SE SI
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.19u L=0.06u
MNA1024 NFB S VSS VPW NCH W=0.2u L=0.06u
MNA1032 NET0128 D VSS VPW NCH W=0.2u L=0.06u
MNA1040 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1044 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1048 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1052 NM M VSS VPW NCH W=0.15u L=0.06u
MNA1056 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET144 NSEMUX VSS VPW NCH W=0.2u L=0.06u
MNA1068 Q NS VSS VPW NCH W=0.28u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.15u L=0.06u
MNOE028 NENMUX E NET0128 VPW NCH W=0.2u L=0.06u
MNOE036 NS BCLK NM VPW NCH W=0.15u L=0.06u
MNOE060 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE072 NSEMUX NSE NENMUX VPW NCH W=0.2u L=0.06u
MNOE076 NENMUX NEN NFB VPW NCH W=0.2u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NEN E VDD VNW PCH W=0.26u L=0.06u
MPA1026 NFB S VDD VNW PCH W=0.3u L=0.06u
MPA1034 NET0128 D VDD VNW PCH W=0.4u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.25u L=0.06u
MPA1042 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1046 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1050 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1054 NM M VDD VNW PCH W=0.2u L=0.06u
MPA1058 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1066 NET144 NSEMUX VDD VNW PCH W=0.2u L=0.06u
MPA1070 Q NS VDD VNW PCH W=0.37u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.25u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.15u L=0.06u
MPOEN030 NENMUX NEN NET0128 VNW PCH W=0.25u L=0.06u
MPOEN038 NS NCLK NM VNW PCH W=0.15u L=0.06u
MPOEN062 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN074 NSEMUX SE NENMUX VNW PCH W=0.25u L=0.06u
MPOEN078 NENMUX E NFB VNW PCH W=0.25u L=0.06u
.ENDS	ESDFFQX0P5MA10TR

****
.SUBCKT ESDFFQX1MA10TR  VDD VSS VPW VNW Q   CK E D SE SI
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.27u L=0.06u
MNA1024 NFB S VSS VPW NCH W=0.22u L=0.06u
MNA1032 NET0135 D VSS VPW NCH W=0.22u L=0.06u
MNA1040 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1044 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1048 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1052 NM M VSS VPW NCH W=0.32u L=0.06u
MNA1056 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET144 NSEMUX VSS VPW NCH W=0.28u L=0.06u
MNA1068 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.28u L=0.06u
MNOE028 NENMUX E NET0135 VPW NCH W=0.22u L=0.06u
MNOE036 NS BCLK NM VPW NCH W=0.28u L=0.06u
MNOE060 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE072 NSEMUX NSE NENMUX VPW NCH W=0.22u L=0.06u
MNOE076 NENMUX NEN NFB VPW NCH W=0.22u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NEN E VDD VNW PCH W=0.36u L=0.06u
MPA1026 NFB S VDD VNW PCH W=0.44u L=0.06u
MPA1034 NET0135 D VDD VNW PCH W=0.44u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1046 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1050 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1054 NM M VDD VNW PCH W=0.48u L=0.06u
MPA1058 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1066 NET144 NSEMUX VDD VNW PCH W=0.28u L=0.06u
MPA1070 Q NS VDD VNW PCH W=0.7u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.28u L=0.06u
MPOEN030 NENMUX NEN NET0135 VNW PCH W=0.33u L=0.06u
MPOEN038 NS NCLK NM VNW PCH W=0.28u L=0.06u
MPOEN062 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN074 NSEMUX SE NENMUX VNW PCH W=0.33u L=0.06u
MPOEN078 NENMUX E NFB VNW PCH W=0.33u L=0.06u
.ENDS	ESDFFQX1MA10TR

****
.SUBCKT ESDFFQX2MA10TR  VDD VSS VPW VNW Q   CK E D SE SI
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.24u L=0.06u
MNA1024 NFB S VSS VPW NCH W=0.3u L=0.06u
MNA1032 NET0135 D VSS VPW NCH W=0.3u L=0.06u
MNA1040 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1044 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1048 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1052 NM M VSS VPW NCH W=0.4u L=0.06u
MNA1056 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET144 NSEMUX VSS VPW NCH W=0.4u L=0.06u
MNA1068 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.4u L=0.06u
MNOE028 NENMUX E NET0135 VPW NCH W=0.3u L=0.06u
MNOE036 NS BCLK NM VPW NCH W=0.4u L=0.06u
MNOE060 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE072 NSEMUX NSE NENMUX VPW NCH W=0.3u L=0.06u
MNOE076 NENMUX NEN NFB VPW NCH W=0.3u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NEN E VDD VNW PCH W=0.31u L=0.06u
MPA1026 NFB S VDD VNW PCH W=0.6u L=0.06u
MPA1034 NET0135 D VDD VNW PCH W=0.6u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1046 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1050 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1054 NM M VDD VNW PCH W=0.6u L=0.06u
MPA1058 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1066 NET144 NSEMUX VDD VNW PCH W=0.4u L=0.06u
MPA1070 Q NS VDD VNW PCH W=1.4u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.4u L=0.06u
MPOEN030 NENMUX NEN NET0135 VNW PCH W=0.45u L=0.06u
MPOEN038 NS NCLK NM VNW PCH W=0.4u L=0.06u
MPOEN062 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN074 NSEMUX SE NENMUX VNW PCH W=0.45u L=0.06u
MPOEN078 NENMUX E NFB VNW PCH W=0.45u L=0.06u
.ENDS	ESDFFQX2MA10TR

****
.SUBCKT ESDFFQX3MA10TR  VDD VSS VPW VNW Q   CK E D SE SI
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.24u L=0.06u
MNA1024 NFB S VSS VPW NCH W=0.3u L=0.06u
MNA1032 NET0135 D VSS VPW NCH W=0.3u L=0.06u
MNA1040 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1044 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1048 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1052 NM M VSS VPW NCH W=0.5u L=0.06u
MNA1056 NET144 NSEMUX VSS VPW NCH W=0.45u L=0.06u
MNA1060 Q NS VSS VPW NCH W=1.59u L=0.06u
MNA1072 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.45u L=0.06u
MNOE028 NENMUX E NET0135 VPW NCH W=0.3u L=0.06u
MNOE036 NS BCLK NM VPW NCH W=0.4u L=0.06u
MNOE064 NSEMUX NSE NENMUX VPW NCH W=0.3u L=0.06u
MNOE068 NENMUX NEN NFB VPW NCH W=0.3u L=0.06u
MNOE076 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NEN E VDD VNW PCH W=0.31u L=0.06u
MPA1026 NFB S VDD VNW PCH W=0.6u L=0.06u
MPA1034 NET0135 D VDD VNW PCH W=0.6u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1046 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1050 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1054 NM M VDD VNW PCH W=0.7u L=0.06u
MPA1058 NET144 NSEMUX VDD VNW PCH W=0.45u L=0.06u
MPA1062 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1074 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.45u L=0.06u
MPOEN030 NENMUX NEN NET0135 VNW PCH W=0.45u L=0.06u
MPOEN038 NS NCLK NM VNW PCH W=0.58u L=0.06u
MPOEN066 NSEMUX SE NENMUX VNW PCH W=0.45u L=0.06u
MPOEN070 NENMUX E NFB VNW PCH W=0.45u L=0.06u
MPOEN078 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
.ENDS	ESDFFQX3MA10TR

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****
.SUBCKT INVX0P5BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.18u L=0.06u
MPA1 Y A VDD VNW PCH W=0.35u L=0.06u
.ENDS	INVX0P5BA10TR

****
.SUBCKT INVX0P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.265u L=0.06u
MPA1 Y A VDD VNW PCH W=0.35u L=0.06u
.ENDS	INVX0P5MA10TR

****
.SUBCKT INVX0P6BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.215u L=0.06u
MPA1 Y A VDD VNW PCH W=0.42u L=0.06u
.ENDS	INVX0P6BA10TR

****
.SUBCKT INVX0P6MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.32u L=0.06u
MPA1 Y A VDD VNW PCH W=0.42u L=0.06u
.ENDS	INVX0P6MA10TR

****
.SUBCKT INVX0P7BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.255u L=0.06u
MPA1 Y A VDD VNW PCH W=0.49u L=0.06u
.ENDS	INVX0P7BA10TR

****
.SUBCKT INVX0P7MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.37u L=0.06u
MPA1 Y A VDD VNW PCH W=0.49u L=0.06u
.ENDS	INVX0P7MA10TR

****
.SUBCKT INVX0P8BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.29u L=0.06u
MPA1 Y A VDD VNW PCH W=0.56u L=0.06u
.ENDS	INVX0P8BA10TR

****
.SUBCKT INVX0P8MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.425u L=0.06u
MPA1 Y A VDD VNW PCH W=0.56u L=0.06u
.ENDS	INVX0P8MA10TR

****
.SUBCKT INVX11BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=3.96u L=0.06u
MPA1 Y A VDD VNW PCH W=7.7u L=0.06u
.ENDS	INVX11BA10TR

****
.SUBCKT INVX11MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=5.83u L=0.06u
MPA1 Y A VDD VNW PCH W=7.7u L=0.06u
.ENDS	INVX11MA10TR

****
.SUBCKT INVX13BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=4.68u L=0.06u
MPA1 Y A VDD VNW PCH W=9.1u L=0.06u
.ENDS	INVX13BA10TR

****
.SUBCKT INVX13MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=6.89u L=0.06u
MPA1 Y A VDD VNW PCH W=9.1u L=0.06u
.ENDS	INVX13MA10TR

****
.SUBCKT INVX16BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=5.76u L=0.06u
MPA1 Y A VDD VNW PCH W=11.2u L=0.06u
.ENDS	INVX16BA10TR

****
.SUBCKT INVX16MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=8.48u L=0.06u
MPA1 Y A VDD VNW PCH W=11.2u L=0.06u
.ENDS	INVX16MA10TR


****
.SUBCKT INVX1BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.36u L=0.06u
MPA1 Y A VDD VNW PCH W=0.7u L=0.06u
.ENDS	INVX1BA10TR


****
.SUBCKT INVX1MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.53u L=0.06u
MPA1 Y A VDD VNW PCH W=0.7u L=0.06u
.ENDS	INVX1MA10TR

****
.SUBCKT INVX1P2BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.43u L=0.06u
MPA1 Y A VDD VNW PCH W=0.84u L=0.06u
.ENDS	INVX1P2BA10TR

****
.SUBCKT INVX1P2MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.635u L=0.06u
MPA1 Y A VDD VNW PCH W=0.84u L=0.06u
.ENDS	INVX1P2MA10TR

****
.SUBCKT INVX1P4BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.505u L=0.06u
MPA1 Y A VDD VNW PCH W=0.98u L=0.06u
.ENDS	INVX1P4BA10TR

****
.SUBCKT INVX1P4MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.74u L=0.06u
MPA1 Y A VDD VNW PCH W=0.98u L=0.06u
.ENDS	INVX1P4MA10TR

****
.SUBCKT INVX1P7BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.61u L=0.06u
MPA1 Y A VDD VNW PCH W=1.19u L=0.06u
.ENDS	INVX1P7BA10TR

****
.SUBCKT INVX1P7MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.9u L=0.06u
MPA1 Y A VDD VNW PCH W=1.19u L=0.06u
.ENDS	INVX1P7MA10TR

****
.SUBCKT INVX2BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.72u L=0.06u
MPA1 Y A VDD VNW PCH W=1.4u L=0.06u
.ENDS	INVX2BA10TR

****
.SUBCKT INVX2MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=1.06u L=0.06u
MPA1 Y A VDD VNW PCH W=1.4u L=0.06u
.ENDS	INVX2MA10TR

****
.SUBCKT INVX2P5BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=0.9u L=0.06u
MPA1 Y A VDD VNW PCH W=1.75u L=0.06u
.ENDS	INVX2P5BA10TR

****
.SUBCKT INVX2P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=1.325u L=0.06u
MPA1 Y A VDD VNW PCH W=1.75u L=0.06u
.ENDS	INVX2P5MA10TR

****
.SUBCKT INVX3BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=1.08u L=0.06u
MPA1 Y A VDD VNW PCH W=2.1u L=0.06u
.ENDS	INVX3BA10TR

****
.SUBCKT INVX3MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=1.59u L=0.06u
MPA1 Y A VDD VNW PCH W=2.1u L=0.06u
.ENDS	INVX3MA10TR

****
.SUBCKT INVX3P5BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=1.26u L=0.06u
MPA1 Y A VDD VNW PCH W=2.45u L=0.06u
.ENDS	INVX3P5BA10TR

****
.SUBCKT INVX3P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=1.855u L=0.06u
MPA1 Y A VDD VNW PCH W=2.45u L=0.06u
.ENDS	INVX3P5MA10TR

****
.SUBCKT INVX4BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=1.44u L=0.06u
MPA1 Y A VDD VNW PCH W=2.8u L=0.06u
.ENDS	INVX4BA10TR

****
.SUBCKT INVX4MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=2.12u L=0.06u
MPA1 Y A VDD VNW PCH W=2.8u L=0.06u
.ENDS	INVX4MA10TR

****
.SUBCKT INVX5BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=1.8u L=0.06u
MPA1 Y A VDD VNW PCH W=3.5u L=0.06u
.ENDS	INVX5BA10TR

****
.SUBCKT INVX5MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=2.65u L=0.06u
MPA1 Y A VDD VNW PCH W=3.5u L=0.06u
.ENDS	INVX5MA10TR

****
.SUBCKT INVX6BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=2.16u L=0.06u
MPA1 Y A VDD VNW PCH W=4.2u L=0.06u
.ENDS	INVX6BA10TR

****
.SUBCKT INVX6MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=3.18u L=0.06u
MPA1 Y A VDD VNW PCH W=4.2u L=0.06u
.ENDS	INVX6MA10TR

****
.SUBCKT INVX7P5BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=2.7u L=0.06u
MPA1 Y A VDD VNW PCH W=5.25u L=0.06u
.ENDS	INVX7P5BA10TR

****
.SUBCKT INVX7P5MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=3.975u L=0.06u
MPA1 Y A VDD VNW PCH W=5.25u L=0.06u
.ENDS	INVX7P5MA10TR

****
.SUBCKT INVX9BA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=3.24u L=0.06u
MPA1 Y A VDD VNW PCH W=6.3u L=0.06u
.ENDS	INVX9BA10TR

****
.SUBCKT INVX9MA10TR  VDD VSS VPW VNW Y   A
MNA1 Y A VSS VPW NCH W=4.77u L=0.06u
MPA1 Y A VDD VNW PCH W=6.3u L=0.06u
.ENDS	INVX9MA10TR

****
.SUBCKT LATNQNX0P5MA10TR  VDD VSS VPW VNW QN   GN D
MNA1 M NM VSS VPW NCH W=0.21u L=0.06u
MNA1012 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.15u L=0.06u
MNA1020 QN M VSS VPW NCH W=0.27u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.15u L=0.06u
MNOE08 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.25u L=0.06u
MPA1014 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.25u L=0.06u
MPA1022 QN M VDD VNW PCH W=0.35u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.15u L=0.06u
MPOEN010 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNQNX0P5MA10TR

****
.SUBCKT LATNQNX1MA10TR  VDD VSS VPW VNW QN   GN D
MNA1 M NM VSS VPW NCH W=0.27u L=0.06u
MNA1012 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.32u L=0.06u
MNA1020 QN M VSS VPW NCH W=0.53u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.28u L=0.06u
MNOE08 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.35u L=0.06u
MPA1014 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.48u L=0.06u
MPA1022 QN M VDD VNW PCH W=0.7u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.28u L=0.06u
MPOEN010 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNQNX1MA10TR

****
.SUBCKT LATNQNX2MA10TR  VDD VSS VPW VNW QN   GN D
MNA1 M NM VSS VPW NCH W=0.51u L=0.06u
MNA1012 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA1020 QN M VSS VPW NCH W=1.06u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.4u L=0.06u
MNOE08 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.61u L=0.06u
MPA1014 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.6u L=0.06u
MPA1022 QN M VDD VNW PCH W=1.4u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.4u L=0.06u
MPOEN010 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNQNX2MA10TR

****
.SUBCKT LATNQNX3MA10TR  VDD VSS VPW VNW QN   GN D
MNA1 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1012 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.45u L=0.06u
MNA1020 QN M VSS VPW NCH W=1.59u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.45u L=0.06u
MNOE08 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1014 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1022 QN M VDD VNW PCH W=2.1u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.45u L=0.06u
MPOEN010 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNQNX3MA10TR

****
.SUBCKT LATNQNX4MA10TR  VDD VSS VPW VNW QN   GN D
MNA1 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1012 NCLK_ GN VSS VPW NCH W=0.18u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA1020 QN M VSS VPW NCH W=2.12u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.58u L=0.06u
MNOE08 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1014 NCLK_ GN VDD VNW PCH W=0.23u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1022 QN M VDD VNW PCH W=2.8u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.58u L=0.06u
MPOEN010 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNQNX4MA10TR

****
.SUBCKT LATNQX0P5MA10TR  VDD VSS VPW VNW Q   GN D
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.15u L=0.06u
MNA1020 Q NM VSS VPW NCH W=0.29u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.15u L=0.06u
MNOE08 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.25u L=0.06u
MPA1022 Q NM VDD VNW PCH W=0.35u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.15u L=0.06u
MPOEN010 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNQX0P5MA10TR

****
.SUBCKT LATNQX1MA10TR  VDD VSS VPW VNW Q   GN D
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.32u L=0.06u
MNA1020 Q NM VSS VPW NCH W=0.58u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.28u L=0.06u
MNOE08 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.48u L=0.06u
MPA1022 Q NM VDD VNW PCH W=0.7u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.28u L=0.06u
MPOEN010 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNQX1MA10TR

****
.SUBCKT LATNQX2MA10TR  VDD VSS VPW VNW Q   GN D
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.47u L=0.06u
MNA1020 Q NM VSS VPW NCH W=1.16u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.4u L=0.06u
MNOE08 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1022 Q NM VDD VNW PCH W=1.4u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.4u L=0.06u
MPOEN010 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNQX2MA10TR

****
.SUBCKT LATNQX3MA10TR  VDD VSS VPW VNW Q   GN D
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ GN VSS VPW NCH W=0.18u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA1020 Q NM VSS VPW NCH W=1.74u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.58u L=0.06u
MNOE08 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ GN VDD VNW PCH W=0.23u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1022 Q NM VDD VNW PCH W=2.1u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.58u L=0.06u
MPOEN010 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNQX3MA10TR

****
.SUBCKT LATNRPQNX0P5MA10TR  VDD VSS VPW VNW QN   GN R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.21u L=0.06u
MNA1022 QN M VSS VPW NCH W=0.27u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.21u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.15u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.25u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.44u L=0.06u
MPA1024 QN M VDD VNW PCH W=0.35u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.44u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.15u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNRPQNX0P5MA10TR

****
.SUBCKT LATNRPQNX1MA10TR  VDD VSS VPW VNW QN   GN R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.32u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.37u L=0.06u
MNA1022 QN M VSS VPW NCH W=0.58u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.37u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.28u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.48u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.65u L=0.06u
MPA1024 QN M VDD VNW PCH W=0.7u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.65u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.28u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNRPQNX1MA10TR

****
.SUBCKT LATNRPQNX2MA10TR  VDD VSS VPW VNW QN   GN R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.5u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.38u L=0.06u
MNA1022 QN M VSS VPW NCH W=1.16u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.38u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.4u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.6u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.7u L=0.06u
MPA1024 QN M VDD VNW PCH W=1.4u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.7u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.4u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNRPQNX2MA10TR

****
.SUBCKT LATNRPQNX3MA10TR  VDD VSS VPW VNW QN   GN R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.45u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.3u L=0.06u
MNA1022 QN M VSS VPW NCH W=1.74u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.3u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.45u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.7u L=0.06u
MPA1024 QN M VDD VNW PCH W=2.1u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.7u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.45u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNRPQNX3MA10TR

****
.SUBCKT LATNRPQNX4MA10TR  VDD VSS VPW VNW QN   GN R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.3u L=0.06u
MNA1022 QN M VSS VPW NCH W=2.32u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.18u L=0.06u
MNA2 M R VSS VPW NCH W=0.3u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.58u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.23u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.7u L=0.06u
MPA1024 QN M VDD VNW PCH W=2.8u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.7u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.58u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNRPQNX4MA10TR

****
.SUBCKT LATNRQX0P5MA10TR  VDD VSS VPW VNW Q   GN RN D
MN0 NIN D NET031 VPW NCH W=0.31u L=0.06u
MN1 NET031 RN VSS VPW NCH W=0.31u L=0.06u
MN2 NM GN NET23 VPW NCH W=0.2u L=0.06u
MN3 NET23 M NET20 VPW NCH W=0.2u L=0.06u
MN4 NET20 RN VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.265u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.15u L=0.06u
MP0 NIN D VDD VNW PCH W=0.3u L=0.06u
MP1 NM RN VDD VNW PCH W=0.5u L=0.06u
MP2 NET33 M VDD VNW PCH W=0.15u L=0.06u
MP3 NM NCLK_ NET33 VNW PCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.35u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.15u L=0.06u
.ENDS	LATNRQX0P5MA10TR

****
.SUBCKT LATNRQX1MA10TR  VDD VSS VPW VNW Q   GN RN D
MN0 NIN D NET031 VPW NCH W=0.51u L=0.06u
MN1 NET031 RN VSS VPW NCH W=0.51u L=0.06u
MN2 NM GN NET23 VPW NCH W=0.2u L=0.06u
MN3 NET23 M NET20 VPW NCH W=0.2u L=0.06u
MN4 NET20 RN VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.53u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.28u L=0.06u
MP0 NIN D VDD VNW PCH W=0.5u L=0.06u
MP1 NM RN VDD VNW PCH W=0.5u L=0.06u
MP2 NET33 M VDD VNW PCH W=0.15u L=0.06u
MP3 NM NCLK_ NET33 VNW PCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.7u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.28u L=0.06u
.ENDS	LATNRQX1MA10TR

****
.SUBCKT LATNRQX2MA10TR  VDD VSS VPW VNW Q   GN RN D
MN0 NIN D NET031 VPW NCH W=0.58u L=0.06u
MN1 NET031 RN VSS VPW NCH W=0.58u L=0.06u
MN2 NM GN NET23 VPW NCH W=0.2u L=0.06u
MN3 NET23 M NET20 VPW NCH W=0.2u L=0.06u
MN4 NET20 RN VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=1.06u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.4u L=0.06u
MP0 NIN D VDD VNW PCH W=0.6u L=0.06u
MP1 NM RN VDD VNW PCH W=0.5u L=0.06u
MP2 NET33 M VDD VNW PCH W=0.15u L=0.06u
MP3 NM NCLK_ NET33 VNW PCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=1.4u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.4u L=0.06u
.ENDS	LATNRQX2MA10TR

****
.SUBCKT LATNRQX3MA10TR  VDD VSS VPW VNW Q   GN RN D
MN0 NIN D NET031 VPW NCH W=0.58u L=0.06u
MN1 NET031 RN VSS VPW NCH W=0.58u L=0.06u
MN2 NM GN NET23 VPW NCH W=0.2u L=0.06u
MN3 NET23 M NET20 VPW NCH W=0.2u L=0.06u
MN4 NET20 RN VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK_ GN VSS VPW NCH W=0.18u L=0.06u
MNA1017 Q NM VSS VPW NCH W=1.59u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.58u L=0.06u
MP0 NIN D VDD VNW PCH W=0.6u L=0.06u
MP1 NM RN VDD VNW PCH W=0.5u L=0.06u
MP2 NET33 M VDD VNW PCH W=0.15u L=0.06u
MP3 NM NCLK_ NET33 VNW PCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK_ GN VDD VNW PCH W=0.23u L=0.06u
MPA1019 Q NM VDD VNW PCH W=2.1u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.58u L=0.06u
.ENDS	LATNRQX3MA10TR

****
.SUBCKT LATNSPQX0P5MA10TR  VDD VSS VPW VNW Q   GN D S
MN0 NIN D VSS VPW NCH W=0.15u L=0.06u
MN2 NM GN NET23 VPW NCH W=0.15u L=0.06u
MN3 NET23 M VSS VPW NCH W=0.15u L=0.06u
MN5 NM S VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.29u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.15u L=0.06u
MP0 NIN D NET045 VNW PCH W=0.45u L=0.06u
MP2 NET33 M NET043 VNW PCH W=0.2u L=0.06u
MP3 NM NCLK_ NET33 VNW PCH W=0.2u L=0.06u
MP4 NET045 S VDD VNW PCH W=0.45u L=0.06u
MP5 NET043 S VDD VNW PCH W=0.2u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.35u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.15u L=0.06u
.ENDS	LATNSPQX0P5MA10TR

****
.SUBCKT LATNSPQX1MA10TR  VDD VSS VPW VNW Q   GN D S
MN0 NIN D VSS VPW NCH W=0.28u L=0.06u
MN2 NM GN NET23 VPW NCH W=0.15u L=0.06u
MN3 NET23 M VSS VPW NCH W=0.15u L=0.06u
MN5 NM S VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.58u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.28u L=0.06u
MP0 NIN D NET045 VNW PCH W=0.7u L=0.06u
MP2 NET33 M NET043 VNW PCH W=0.2u L=0.06u
MP3 NM NCLK_ NET33 VNW PCH W=0.2u L=0.06u
MP4 NET045 S VDD VNW PCH W=0.7u L=0.06u
MP5 NET043 S VDD VNW PCH W=0.2u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.7u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.28u L=0.06u
.ENDS	LATNSPQX1MA10TR

****
.SUBCKT LATNSPQX2MA10TR  VDD VSS VPW VNW Q   GN D S
MN0 NIN D VSS VPW NCH W=0.3u L=0.06u
MN2 NM GN NET23 VPW NCH W=0.15u L=0.06u
MN3 NET23 M VSS VPW NCH W=0.15u L=0.06u
MN5 NM S VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=1.16u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.4u L=0.06u
MP0 NIN D NET045 VNW PCH W=0.7u L=0.06u
MP2 NET33 M NET043 VNW PCH W=0.2u L=0.06u
MP3 NM NCLK_ NET33 VNW PCH W=0.2u L=0.06u
MP4 NET045 S VDD VNW PCH W=0.7u L=0.06u
MP5 NET043 S VDD VNW PCH W=0.2u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=1.4u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.4u L=0.06u
.ENDS	LATNSPQX2MA10TR

****

****
.SUBCKT LATNSQNX0P5MA10TR  VDD VSS VPW VNW QN   GN D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.3u L=0.06u
MNA1022 QN M VSS VPW NCH W=0.27u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.3u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.15u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.25u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.25u L=0.06u
MPA1024 QN M VDD VNW PCH W=0.35u L=0.06u
MPA2 M SN VDD VNW PCH W=0.25u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.15u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNSQNX0P5MA10TR

****
.SUBCKT LATNSQNX1MA10TR  VDD VSS VPW VNW QN   GN D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.32u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.4u L=0.06u
MNA1022 QN M VSS VPW NCH W=0.53u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.4u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.28u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.48u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.35u L=0.06u
MPA1024 QN M VDD VNW PCH W=0.7u L=0.06u
MPA2 M SN VDD VNW PCH W=0.35u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.28u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNSQNX1MA10TR

****
.SUBCKT LATNSQNX2MA10TR  VDD VSS VPW VNW QN   GN D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.58u L=0.06u
MNA1022 QN M VSS VPW NCH W=1.06u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.58u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.4u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.5u L=0.06u
MPA1024 QN M VDD VNW PCH W=1.4u L=0.06u
MPA2 M SN VDD VNW PCH W=0.5u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.4u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNSQNX2MA10TR

****
.SUBCKT LATNSQNX3MA10TR  VDD VSS VPW VNW QN   GN D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.45u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.58u L=0.06u
MNA1022 QN M VSS VPW NCH W=1.59u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.58u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.45u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.5u L=0.06u
MPA1024 QN M VDD VNW PCH W=2.1u L=0.06u
MPA2 M SN VDD VNW PCH W=0.5u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.45u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNSQNX3MA10TR

****
.SUBCKT LATNSQNX4MA10TR  VDD VSS VPW VNW QN   GN D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.58u L=0.06u
MNA1022 QN M VSS VPW NCH W=2.12u L=0.06u
MNA108 NCLK_ GN VSS VPW NCH W=0.18u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.58u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.58u L=0.06u
MNOE04 NM GN N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK_ GN VDD VNW PCH W=0.23u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.5u L=0.06u
MPA1024 QN M VDD VNW PCH W=2.8u L=0.06u
MPA2 M SN VDD VNW PCH W=0.5u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.58u L=0.06u
MPOEN06 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATNSQNX4MA10TR

****
.SUBCKT LATQNX0P5MA10TR  VDD VSS VPW VNW QN   G D
MNA1 M NM VSS VPW NCH W=0.21u L=0.06u
MNA1012 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.15u L=0.06u
MNA1020 QN M VSS VPW NCH W=0.27u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM G NIN VPW NCH W=0.15u L=0.06u
MNOE08 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.25u L=0.06u
MPA1014 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.25u L=0.06u
MPA1022 QN M VDD VNW PCH W=0.35u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.15u L=0.06u
MPOEN010 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATQNX0P5MA10TR

****
.SUBCKT LATQNX1MA10TR  VDD VSS VPW VNW QN   G D
MNA1 M NM VSS VPW NCH W=0.27u L=0.06u
MNA1012 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.32u L=0.06u
MNA1020 QN M VSS VPW NCH W=0.53u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM G NIN VPW NCH W=0.28u L=0.06u
MNOE08 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.35u L=0.06u
MPA1014 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.48u L=0.06u
MPA1022 QN M VDD VNW PCH W=0.7u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.28u L=0.06u
MPOEN010 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATQNX1MA10TR

****
.SUBCKT LATQNX2MA10TR  VDD VSS VPW VNW QN   G D
MNA1 M NM VSS VPW NCH W=0.51u L=0.06u
MNA1012 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA1020 QN M VSS VPW NCH W=1.06u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM G NIN VPW NCH W=0.4u L=0.06u
MNOE08 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.61u L=0.06u
MPA1014 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.6u L=0.06u
MPA1022 QN M VDD VNW PCH W=1.4u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.4u L=0.06u
MPOEN010 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATQNX2MA10TR

****
.SUBCKT LATQNX3MA10TR  VDD VSS VPW VNW QN   G D
MNA1 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1012 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.45u L=0.06u
MNA1020 QN M VSS VPW NCH W=1.59u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM G NIN VPW NCH W=0.45u L=0.06u
MNOE08 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1014 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1022 QN M VDD VNW PCH W=2.1u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.45u L=0.06u
MPOEN010 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATQNX3MA10TR

****
.SUBCKT LATQNX4MA10TR  VDD VSS VPW VNW QN   G D
MNA1 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1012 NCLK G VSS VPW NCH W=0.18u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA1020 QN M VSS VPW NCH W=2.12u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM G NIN VPW NCH W=0.58u L=0.06u
MNOE08 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1014 NCLK G VDD VNW PCH W=0.23u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1022 QN M VDD VNW PCH W=2.8u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.58u L=0.06u
MPOEN010 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATQNX4MA10TR

****
.SUBCKT LATQX0P5MA10TR  VDD VSS VPW VNW Q   G D
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.15u L=0.06u
MNA1020 Q NM VSS VPW NCH W=0.29u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM G NIN VPW NCH W=0.15u L=0.06u
MNOE08 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.25u L=0.06u
MPA1022 Q NM VDD VNW PCH W=0.35u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.15u L=0.06u
MPOEN010 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATQX0P5MA10TR

****
.SUBCKT LATQX1MA10TR  VDD VSS VPW VNW Q   G D
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.32u L=0.06u
MNA1020 Q NM VSS VPW NCH W=0.58u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM G NIN VPW NCH W=0.28u L=0.06u
MNOE08 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.48u L=0.06u
MPA1022 Q NM VDD VNW PCH W=0.7u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.28u L=0.06u
MPOEN010 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATQX1MA10TR

****
.SUBCKT LATQX2MA10TR  VDD VSS VPW VNW Q   G D
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.47u L=0.06u
MNA1020 Q NM VSS VPW NCH W=1.16u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM G NIN VPW NCH W=0.4u L=0.06u
MNOE08 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1022 Q NM VDD VNW PCH W=1.4u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.4u L=0.06u
MPOEN010 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATQX2MA10TR

****
.SUBCKT LATQX3MA10TR  VDD VSS VPW VNW Q   G D
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK G VSS VPW NCH W=0.18u L=0.06u
MNA1016 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA1020 Q NM VSS VPW NCH W=1.74u L=0.06u
MNA104 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM G NIN VPW NCH W=0.58u L=0.06u
MNOE08 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK G VDD VNW PCH W=0.23u L=0.06u
MPA1018 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1022 Q NM VDD VNW PCH W=2.1u L=0.06u
MPA106 P1 M VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.58u L=0.06u
MPOEN010 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATQX3MA10TR

****
.SUBCKT LATRPQNX0P5MA10TR  VDD VSS VPW VNW QN   G R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.21u L=0.06u
MNA1022 QN M VSS VPW NCH W=0.27u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.21u L=0.06u
MNOE NM G NIN VPW NCH W=0.15u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.25u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.44u L=0.06u
MPA1024 QN M VDD VNW PCH W=0.35u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.44u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.15u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATRPQNX0P5MA10TR

****
.SUBCKT LATRPQNX1MA10TR  VDD VSS VPW VNW QN   G R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.32u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.37u L=0.06u
MNA1022 QN M VSS VPW NCH W=0.58u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.37u L=0.06u
MNOE NM G NIN VPW NCH W=0.28u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.48u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.65u L=0.06u
MPA1024 QN M VDD VNW PCH W=0.7u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.65u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.28u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATRPQNX1MA10TR

****
.SUBCKT LATRPQNX2MA10TR  VDD VSS VPW VNW QN   G R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.5u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.38u L=0.06u
MNA1022 QN M VSS VPW NCH W=1.16u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.38u L=0.06u
MNOE NM G NIN VPW NCH W=0.4u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.6u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.7u L=0.06u
MPA1024 QN M VDD VNW PCH W=1.4u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.7u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.4u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATRPQNX2MA10TR

****
.SUBCKT LATRPQNX3MA10TR  VDD VSS VPW VNW QN   G R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.45u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.3u L=0.06u
MNA1022 QN M VSS VPW NCH W=1.74u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.3u L=0.06u
MNOE NM G NIN VPW NCH W=0.45u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.7u L=0.06u
MPA1024 QN M VDD VNW PCH W=2.1u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.7u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.45u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATRPQNX3MA10TR

****
.SUBCKT LATRPQNX4MA10TR  VDD VSS VPW VNW QN   G R D
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.3u L=0.06u
MNA1022 QN M VSS VPW NCH W=2.32u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.18u L=0.06u
MNA2 M R VSS VPW NCH W=0.3u L=0.06u
MNOE NM G NIN VPW NCH W=0.58u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.23u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM P1_6 VNW PCH W=0.7u L=0.06u
MPA1024 QN M VDD VNW PCH W=2.8u L=0.06u
MPA2 P1_6 R VDD VNW PCH W=0.7u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.58u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATRPQNX4MA10TR

****
.SUBCKT LATRQX0P5MA10TR  VDD VSS VPW VNW Q   G RN D
MN0 NIN D NET27 VPW NCH W=0.31u L=0.06u
MN1 NET27 RN VSS VPW NCH W=0.31u L=0.06u
MN2 NM NCLK NET23 VPW NCH W=0.2u L=0.06u
MN3 NET23 M NET20 VPW NCH W=0.2u L=0.06u
MN4 NET20 RN VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.265u L=0.06u
MNOE NM G NIN VPW NCH W=0.15u L=0.06u
MP0 NIN D VDD VNW PCH W=0.3u L=0.06u
MP1 NM RN VDD VNW PCH W=0.3u L=0.06u
MP2 NET33 M VDD VNW PCH W=0.15u L=0.06u
MP3 NM G NET33 VNW PCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.35u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.15u L=0.06u
.ENDS	LATRQX0P5MA10TR

****
.SUBCKT LATRQX1MA10TR  VDD VSS VPW VNW Q   G RN D
MN0 NIN D NET27 VPW NCH W=0.51u L=0.06u
MN1 NET27 RN VSS VPW NCH W=0.51u L=0.06u
MN2 NM NCLK NET23 VPW NCH W=0.2u L=0.06u
MN3 NET23 M NET20 VPW NCH W=0.2u L=0.06u
MN4 NET20 RN VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.53u L=0.06u
MNOE NM G NIN VPW NCH W=0.28u L=0.06u
MP0 NIN D VDD VNW PCH W=0.5u L=0.06u
MP1 NM RN VDD VNW PCH W=0.3u L=0.06u
MP2 NET33 M VDD VNW PCH W=0.15u L=0.06u
MP3 NM G NET33 VNW PCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.7u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.28u L=0.06u
.ENDS	LATRQX1MA10TR

****
.SUBCKT LATRQX2MA10TR  VDD VSS VPW VNW Q   G RN D
MN0 NIN D NET27 VPW NCH W=0.58u L=0.06u
MN1 NET27 RN VSS VPW NCH W=0.58u L=0.06u
MN2 NM NCLK NET23 VPW NCH W=0.2u L=0.06u
MN3 NET23 M NET20 VPW NCH W=0.2u L=0.06u
MN4 NET20 RN VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=1.06u L=0.06u
MNOE NM G NIN VPW NCH W=0.4u L=0.06u
MP0 NIN D VDD VNW PCH W=0.6u L=0.06u
MP1 NM RN VDD VNW PCH W=0.3u L=0.06u
MP2 NET33 M VDD VNW PCH W=0.15u L=0.06u
MP3 NM G NET33 VNW PCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=1.4u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.4u L=0.06u
.ENDS	LATRQX2MA10TR

****
.SUBCKT LATRQX3MA10TR  VDD VSS VPW VNW Q   G RN D
MN0 NIN D NET27 VPW NCH W=0.58u L=0.06u
MN1 NET27 RN VSS VPW NCH W=0.58u L=0.06u
MN2 NM NCLK NET23 VPW NCH W=0.2u L=0.06u
MN3 NET23 M NET20 VPW NCH W=0.2u L=0.06u
MN4 NET20 RN VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK G VSS VPW NCH W=0.18u L=0.06u
MNA1017 Q NM VSS VPW NCH W=1.59u L=0.06u
MNOE NM G NIN VPW NCH W=0.58u L=0.06u
MP0 NIN D VDD VNW PCH W=0.6u L=0.06u
MP1 NM RN VDD VNW PCH W=0.3u L=0.06u
MP2 NET33 M VDD VNW PCH W=0.15u L=0.06u
MP3 NM G NET33 VNW PCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK G VDD VNW PCH W=0.23u L=0.06u
MPA1019 Q NM VDD VNW PCH W=2.1u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.58u L=0.06u
.ENDS	LATRQX3MA10TR

****
.SUBCKT LATSPQX0P5MA10TR  VDD VSS VPW VNW Q   G D S
MN0 NIN D VSS VPW NCH W=0.15u L=0.06u
MN2 NM NCLK NET23 VPW NCH W=0.15u L=0.06u
MN3 NET23 M VSS VPW NCH W=0.15u L=0.06u
MN5 NM S VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.29u L=0.06u
MNOE NM G NIN VPW NCH W=0.15u L=0.06u
MP0 NIN D NET048 VNW PCH W=0.45u L=0.06u
MP2 NET33 M NET043 VNW PCH W=0.2u L=0.06u
MP3 NM G NET33 VNW PCH W=0.2u L=0.06u
MP4 NET048 S VDD VNW PCH W=0.45u L=0.06u
MP5 NET043 S VDD VNW PCH W=0.2u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.35u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.15u L=0.06u
.ENDS	LATSPQX0P5MA10TR

****
.SUBCKT LATSPQX1MA10TR  VDD VSS VPW VNW Q   G D S
MN0 NIN D VSS VPW NCH W=0.28u L=0.06u
MN2 NM NCLK NET23 VPW NCH W=0.15u L=0.06u
MN3 NET23 M VSS VPW NCH W=0.15u L=0.06u
MN5 NM S VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.58u L=0.06u
MNOE NM G NIN VPW NCH W=0.28u L=0.06u
MP0 NIN D NET048 VNW PCH W=0.7u L=0.06u
MP2 NET33 M NET043 VNW PCH W=0.2u L=0.06u
MP3 NM G NET33 VNW PCH W=0.2u L=0.06u
MP4 NET048 S VDD VNW PCH W=0.7u L=0.06u
MP5 NET043 S VDD VNW PCH W=0.2u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.7u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.28u L=0.06u
.ENDS	LATSPQX1MA10TR

****
.SUBCKT LATSPQX2MA10TR  VDD VSS VPW VNW Q   G D S
MN0 NIN D VSS VPW NCH W=0.3u L=0.06u
MN2 NM NCLK NET23 VPW NCH W=0.15u L=0.06u
MN3 NET23 M VSS VPW NCH W=0.15u L=0.06u
MN5 NM S VSS VPW NCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1013 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=1.16u L=0.06u
MNOE NM G NIN VPW NCH W=0.4u L=0.06u
MP0 NIN D NET048 VNW PCH W=0.7u L=0.06u
MP2 NET33 M NET043 VNW PCH W=0.2u L=0.06u
MP3 NM G NET33 VNW PCH W=0.2u L=0.06u
MP4 NET048 S VDD VNW PCH W=0.7u L=0.06u
MP5 NET043 S VDD VNW PCH W=0.2u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MPA1015 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1019 Q NM VDD VNW PCH W=1.4u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.4u L=0.06u
.ENDS	LATSPQX2MA10TR

****

****
.SUBCKT LATSQNX0P5MA10TR  VDD VSS VPW VNW QN   G D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.3u L=0.06u
MNA1022 QN M VSS VPW NCH W=0.27u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.3u L=0.06u
MNOE NM G NIN VPW NCH W=0.15u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.25u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.25u L=0.06u
MPA1024 QN M VDD VNW PCH W=0.35u L=0.06u
MPA2 M SN VDD VNW PCH W=0.25u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.15u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATSQNX0P5MA10TR

****
.SUBCKT LATSQNX1MA10TR  VDD VSS VPW VNW QN   G D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.32u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.4u L=0.06u
MNA1022 QN M VSS VPW NCH W=0.53u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.4u L=0.06u
MNOE NM G NIN VPW NCH W=0.28u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.48u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.35u L=0.06u
MPA1024 QN M VDD VNW PCH W=0.7u L=0.06u
MPA2 M SN VDD VNW PCH W=0.35u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.28u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATSQNX1MA10TR

****
.SUBCKT LATSQNX2MA10TR  VDD VSS VPW VNW QN   G D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.4u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.58u L=0.06u
MNA1022 QN M VSS VPW NCH W=1.06u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.58u L=0.06u
MNOE NM G NIN VPW NCH W=0.4u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.5u L=0.06u
MPA1024 QN M VDD VNW PCH W=1.4u L=0.06u
MPA2 M SN VDD VNW PCH W=0.5u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.4u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATSQNX2MA10TR

****
.SUBCKT LATSQNX3MA10TR  VDD VSS VPW VNW QN   G D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.45u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.58u L=0.06u
MNA1022 QN M VSS VPW NCH W=1.59u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.58u L=0.06u
MNOE NM G NIN VPW NCH W=0.45u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.2u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.5u L=0.06u
MPA1024 QN M VDD VNW PCH W=2.1u L=0.06u
MPA2 M SN VDD VNW PCH W=0.5u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.45u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATSQNX3MA10TR

****
.SUBCKT LATSQNX4MA10TR  VDD VSS VPW VNW QN   G D SN
MNA1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NIN D VSS VPW NCH W=0.58u L=0.06u
MNA1016 M NM N1_6 VPW NCH W=0.58u L=0.06u
MNA1022 QN M VSS VPW NCH W=2.12u L=0.06u
MNA108 NCLK G VSS VPW NCH W=0.18u L=0.06u
MNA2 N1_6 SN VSS VPW NCH W=0.58u L=0.06u
MNOE NM G NIN VPW NCH W=0.58u L=0.06u
MNOE04 NM NCLK N1 VPW NCH W=0.15u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1010 NCLK G VDD VNW PCH W=0.23u L=0.06u
MPA1014 NIN D VDD VNW PCH W=0.7u L=0.06u
MPA1019 M NM VDD VNW PCH W=0.5u L=0.06u
MPA1024 QN M VDD VNW PCH W=2.8u L=0.06u
MPA2 M SN VDD VNW PCH W=0.5u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.58u L=0.06u
MPOEN06 NM G P1 VNW PCH W=0.15u L=0.06u
.ENDS	LATSQNX4MA10TR

****
.SUBCKT M2DFFQNX0P5MA10TR  VDD VSS VPW VNW QN   CK D0 D1 S0
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1016 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1020 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1024 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1028 N1_12 NS VSS VPW NCH W=0.15u L=0.06u
MNA1036 QN S VSS VPW NCH W=0.28u L=0.06u
MNA1052 NET155 D1 VSS VPW NCH W=0.3u L=0.06u
MNA1056 NET151 D0 VSS VPW NCH W=0.3u L=0.06u
MNA108 NSEL S0 VSS VPW NCH W=0.21u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE012 S BCLK M VPW NCH W=0.15u L=0.06u
MNOE032 S NCLK N1_12 VPW NCH W=0.15u L=0.06u
MNOE040 NM NCLK NENMUX VPW NCH W=0.15u L=0.06u
MNOE044 NENMUX S0 NET155 VPW NCH W=0.3u L=0.06u
MNOE048 NENMUX NSEL NET151 VPW NCH W=0.3u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1010 NSEL S0 VDD VNW PCH W=0.28u L=0.06u
MPA1018 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1022 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1026 M NM VDD VNW PCH W=0.2u L=0.06u
MPA1030 P1_14 NS VDD VNW PCH W=0.15u L=0.06u
MPA1038 QN S VDD VNW PCH W=0.37u L=0.06u
MPA104 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1054 NET155 D1 VDD VNW PCH W=0.3u L=0.06u
MPA1058 NET151 D0 VDD VNW PCH W=0.3u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN014 S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN034 S BCLK P1_14 VNW PCH W=0.15u L=0.06u
MPOEN042 NM BCLK NENMUX VNW PCH W=0.15u L=0.06u
MPOEN046 NENMUX NSEL NET155 VNW PCH W=0.3u L=0.06u
MPOEN050 NENMUX S0 NET151 VNW PCH W=0.3u L=0.06u
.ENDS	M2DFFQNX0P5MA10TR

****
.SUBCKT M2DFFQNX1MA10TR  VDD VSS VPW VNW QN   CK D0 D1 S0
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.27u L=0.06u
MNA1016 QN S VSS VPW NCH W=0.53u L=0.06u
MNA102 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1024 NET81 D1 VSS VPW NCH W=0.32u L=0.06u
MNA1032 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1036 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 M NM VSS VPW NCH W=0.32u L=0.06u
MNA1048 NET77 D0 VSS VPW NCH W=0.32u L=0.06u
MNA1052 N1_12 NS VSS VPW NCH W=0.15u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE020 NENMUX S0 NET81 VPW NCH W=0.28u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.28u L=0.06u
MNOE044 NENMUX NSEL NET77 VPW NCH W=0.28u L=0.06u
MNOE056 S NCLK N1_12 VPW NCH W=0.15u L=0.06u
MNOE08 NM NCLK NENMUX VPW NCH W=0.28u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.36u L=0.06u
MPA1018 QN S VDD VNW PCH W=0.7u L=0.06u
MPA1026 NET81 D1 VDD VNW PCH W=0.48u L=0.06u
MPA1034 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1038 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA104 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1042 M NM VDD VNW PCH W=0.48u L=0.06u
MPA1050 NET77 D0 VDD VNW PCH W=0.48u L=0.06u
MPA1054 P1_14 NS VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 NM BCLK NENMUX VNW PCH W=0.28u L=0.06u
MPOEN022 NENMUX NSEL NET81 VNW PCH W=0.28u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN046 NENMUX S0 NET77 VNW PCH W=0.28u L=0.06u
MPOEN058 S BCLK P1_14 VNW PCH W=0.15u L=0.06u
.ENDS	M2DFFQNX1MA10TR

****
.SUBCKT M2DFFQNX2MA10TR  VDD VSS VPW VNW QN   CK D0 D1 S0
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.26u L=0.06u
MNA102 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1020 NIN1 D1 VSS VPW NCH W=0.4u L=0.06u
MNA1028 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1032 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1036 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1040 N1_12 NS VSS VPW NCH W=0.15u L=0.06u
MNA1048 QN S VSS VPW NCH W=1.06u L=0.06u
MNA1056 NIN0 D0 VSS VPW NCH W=0.4u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE016 NENMUX S0 NIN1 VPW NCH W=0.4u L=0.06u
MNOE024 S BCLK M VPW NCH W=0.4u L=0.06u
MNOE044 S NCLK N1_12 VPW NCH W=0.15u L=0.06u
MNOE052 NENMUX NSEL NIN0 VPW NCH W=0.4u L=0.06u
MNOE08 NM NCLK NENMUX VPW NCH W=0.4u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.34u L=0.06u
MPA1022 NIN1 D1 VDD VNW PCH W=0.45u L=0.06u
MPA1030 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1034 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1038 M NM VDD VNW PCH W=0.6u L=0.06u
MPA104 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1042 P1_14 NS VDD VNW PCH W=0.15u L=0.06u
MPA1050 QN S VDD VNW PCH W=1.4u L=0.06u
MPA1058 NIN0 D0 VDD VNW PCH W=0.45u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 NM BCLK NENMUX VNW PCH W=0.4u L=0.06u
MPOEN018 NENMUX NSEL NIN1 VNW PCH W=0.4u L=0.06u
MPOEN026 S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN046 S BCLK P1_14 VNW PCH W=0.15u L=0.06u
MPOEN054 NENMUX S0 NIN0 VNW PCH W=0.4u L=0.06u
.ENDS	M2DFFQNX2MA10TR

****
.SUBCKT M2DFFQNX3MA10TR  VDD VSS VPW VNW QN   CK D0 D1 S0
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.28u L=0.06u
MNA102 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1020 NIN1 D1 VSS VPW NCH W=0.5u L=0.06u
MNA1028 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1032 N1_12 NS VSS VPW NCH W=0.15u L=0.06u
MNA1040 QN S VSS VPW NCH W=1.68u L=0.06u
MNA1048 NIN0 D0 VSS VPW NCH W=0.5u L=0.06u
MNA1052 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1056 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE016 NENMUX S0 NIN1 VPW NCH W=0.45u L=0.06u
MNOE024 S BCLK M VPW NCH W=0.58u L=0.06u
MNOE036 S NCLK N1_12 VPW NCH W=0.15u L=0.06u
MNOE044 NENMUX NSEL NIN0 VPW NCH W=0.45u L=0.06u
MNOE08 NM NCLK NENMUX VPW NCH W=0.45u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.37u L=0.06u
MPA1022 NIN1 D1 VDD VNW PCH W=0.6u L=0.06u
MPA1030 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1034 P1_14 NS VDD VNW PCH W=0.15u L=0.06u
MPA104 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1042 QN S VDD VNW PCH W=2.1u L=0.06u
MPA1050 NIN0 D0 VDD VNW PCH W=0.6u L=0.06u
MPA1054 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1058 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 NM BCLK NENMUX VNW PCH W=0.45u L=0.06u
MPOEN018 NENMUX NSEL NIN1 VNW PCH W=0.45u L=0.06u
MPOEN026 S NCLK M VNW PCH W=0.58u L=0.06u
MPOEN038 S BCLK P1_14 VNW PCH W=0.15u L=0.06u
MPOEN046 NENMUX S0 NIN0 VNW PCH W=0.45u L=0.06u
.ENDS	M2DFFQNX3MA10TR

****
.SUBCKT M2DFFQX0P5MA10TR  VDD VSS VPW VNW Q   CK D0 D1 S0
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1024 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1028 NM M VSS VPW NCH W=0.15u L=0.06u
MNA1032 N1_13 S VSS VPW NCH W=0.15u L=0.06u
MNA1040 NET144 NENMUX VSS VPW NCH W=0.15u L=0.06u
MNA1044 Q NS VSS VPW NCH W=0.28u L=0.06u
MNA1056 NET0132 D1 VSS VPW NCH W=0.2u L=0.06u
MNA1060 NET0128 D0 VSS VPW NCH W=0.2u L=0.06u
MNOE M BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE016 NS BCLK NM VPW NCH W=0.15u L=0.06u
MNOE036 NS NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE048 NENMUX S0 NET0132 VPW NCH W=0.2u L=0.06u
MNOE052 NENMUX NSEL NET0128 VPW NCH W=0.2u L=0.06u
MNOE08 M NCLK NET144 VPW NCH W=0.15u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.2u L=0.06u
MPA1022 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1026 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1030 NM M VDD VNW PCH W=0.2u L=0.06u
MPA1034 P1_15 S VDD VNW PCH W=0.15u L=0.06u
MPA104 P1 NM VDD VNW PCH W=0.15u L=0.06u
MPA1042 NET144 NENMUX VDD VNW PCH W=0.15u L=0.06u
MPA1046 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA1058 NET0132 D1 VDD VNW PCH W=0.4u L=0.06u
MPA1062 NET0128 D0 VDD VNW PCH W=0.4u L=0.06u
MPOEN M NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 M BCLK NET144 VNW PCH W=0.15u L=0.06u
MPOEN018 NS NCLK NM VNW PCH W=0.15u L=0.06u
MPOEN038 NS BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN050 NENMUX NSEL NET0132 VNW PCH W=0.2u L=0.06u
MPOEN054 NENMUX S0 NET0128 VNW PCH W=0.2u L=0.06u
.ENDS	M2DFFQX0P5MA10TR

****
.SUBCKT M2DFFQX1MA10TR  VDD VSS VPW VNW Q   CK D0 D1 S0
MNA1 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1010 N1 NM VSS VPW NCH W=0.15u L=0.06u
MNA102 NM M VSS VPW NCH W=0.32u L=0.06u
MNA1024 N1_13 S VSS VPW NCH W=0.15u L=0.06u
MNA1032 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA1036 NET112 NENMUX VSS VPW NCH W=0.28u L=0.06u
MNA1048 NET80 D1 VSS VPW NCH W=0.24u L=0.06u
MNA1052 NET84 D0 VSS VPW NCH W=0.24u L=0.06u
MNA1056 S NS VSS VPW NCH W=0.15u L=0.06u
MNA106 NSEL S0 VSS VPW NCH W=0.26u L=0.06u
MNA1060 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNOE M BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE016 NENMUX S0 NET80 VPW NCH W=0.2u L=0.06u
MNOE020 M NCLK NET112 VPW NCH W=0.28u L=0.06u
MNOE028 NS NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE040 NS BCLK NM VPW NCH W=0.28u L=0.06u
MNOE044 NENMUX NSEL NET84 VPW NCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1012 P1 NM VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_15 S VDD VNW PCH W=0.15u L=0.06u
MPA1034 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA1038 NET112 NENMUX VDD VNW PCH W=0.28u L=0.06u
MPA104 NM M VDD VNW PCH W=0.48u L=0.06u
MPA1050 NET80 D1 VDD VNW PCH W=0.36u L=0.06u
MPA1054 NET84 D0 VDD VNW PCH W=0.36u L=0.06u
MPA1058 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1062 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA108 NSEL S0 VDD VNW PCH W=0.34u L=0.06u
MPOEN M NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN018 NENMUX NSEL NET80 VNW PCH W=0.3u L=0.06u
MPOEN022 M BCLK NET112 VNW PCH W=0.28u L=0.06u
MPOEN030 NS BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN042 NS NCLK NM VNW PCH W=0.28u L=0.06u
MPOEN046 NENMUX S0 NET84 VNW PCH W=0.3u L=0.06u
.ENDS	M2DFFQX1MA10TR

****
.SUBCKT M2DFFQX2MA10TR  VDD VSS VPW VNW Q   CK D0 D1 S0
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.26u L=0.06u
MNA102 N1 NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NET0135 D1 VSS VPW NCH W=0.3u L=0.06u
MNA1028 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1032 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1036 NM M VSS VPW NCH W=0.4u L=0.06u
MNA1040 N1_13 S VSS VPW NCH W=0.15u L=0.06u
MNA1048 NET144 NENMUX VSS VPW NCH W=0.4u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA1060 NET0139 D0 VSS VPW NCH W=0.3u L=0.06u
MNOE M BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE016 NENMUX S0 NET0135 VPW NCH W=0.3u L=0.06u
MNOE024 NS BCLK NM VPW NCH W=0.4u L=0.06u
MNOE044 NS NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE056 NENMUX NSEL NET0139 VPW NCH W=0.3u L=0.06u
MNOE08 M NCLK NET144 VPW NCH W=0.4u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.34u L=0.06u
MPA1022 NET0135 D1 VDD VNW PCH W=0.6u L=0.06u
MPA1030 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1034 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1038 NM M VDD VNW PCH W=0.6u L=0.06u
MPA104 P1 NM VDD VNW PCH W=0.15u L=0.06u
MPA1042 P1_15 S VDD VNW PCH W=0.15u L=0.06u
MPA1050 NET144 NENMUX VDD VNW PCH W=0.4u L=0.06u
MPA1054 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA1062 NET0139 D0 VDD VNW PCH W=0.6u L=0.06u
MPOEN M NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 M BCLK NET144 VNW PCH W=0.4u L=0.06u
MPOEN018 NENMUX NSEL NET0135 VNW PCH W=0.4u L=0.06u
MPOEN026 NS NCLK NM VNW PCH W=0.4u L=0.06u
MPOEN046 NS BCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN058 NENMUX S0 NET0139 VNW PCH W=0.4u L=0.06u
.ENDS	M2DFFQX2MA10TR

****
.SUBCKT M2DFFQX3MA10TR  VDD VSS VPW VNW Q   CK D0 D1 S0
MNA1 NSEL S0 VSS VPW NCH W=0.26u L=0.06u
MNA1012 NM M VSS VPW NCH W=0.58u L=0.06u
MNA102 N1 NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NET0135 D1 VSS VPW NCH W=0.3u L=0.06u
MNA1028 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1032 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1036 NET144 NENMUX VSS VPW NCH W=0.45u L=0.06u
MNA1044 NET0139 D0 VSS VPW NCH W=0.3u L=0.06u
MNA1048 N1_13 S VSS VPW NCH W=0.15u L=0.06u
MNA1056 Q NS VSS VPW NCH W=1.68u L=0.06u
MNA1060 S NS VSS VPW NCH W=0.15u L=0.06u
MNOE M BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE016 NENMUX S0 NET0135 VPW NCH W=0.3u L=0.06u
MNOE024 M NCLK NET144 VPW NCH W=0.45u L=0.06u
MNOE040 NENMUX NSEL NET0139 VPW NCH W=0.3u L=0.06u
MNOE052 NS NCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE08 NS BCLK NM VPW NCH W=0.58u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.34u L=0.06u
MPA1014 NM M VDD VNW PCH W=0.7u L=0.06u
MPA1022 NET0135 D1 VDD VNW PCH W=0.6u L=0.06u
MPA1030 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1034 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1038 NET144 NENMUX VDD VNW PCH W=0.45u L=0.06u
MPA104 P1 NM VDD VNW PCH W=0.15u L=0.06u
MPA1046 NET0139 D0 VDD VNW PCH W=0.6u L=0.06u
MPA1050 P1_15 S VDD VNW PCH W=0.15u L=0.06u
MPA1058 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1062 S NS VDD VNW PCH W=0.15u L=0.06u
MPOEN M NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN010 NS NCLK NM VNW PCH W=0.58u L=0.06u
MPOEN018 NENMUX NSEL NET0135 VNW PCH W=0.4u L=0.06u
MPOEN026 M BCLK NET144 VNW PCH W=0.45u L=0.06u
MPOEN042 NENMUX S0 NET0139 VNW PCH W=0.4u L=0.06u
MPOEN054 NS BCLK P1_15 VNW PCH W=0.15u L=0.06u
.ENDS	M2DFFQX3MA10TR

****
.SUBCKT M2DFFQX4MA10TR  VDD VSS VPW VNW Q   CK D0 D1 S0
MNA1 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1010 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1020 NSEL S0 VSS VPW NCH W=0.26u L=0.06u
MNA1028 NET0135 D1 VSS VPW NCH W=0.58u L=0.06u
MNA1036 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1040 N1_12 NS VSS VPW NCH W=0.15u L=0.06u
MNA1052 NET0139 D0 VSS VPW NCH W=0.58u L=0.06u
MNA1056 Q NS VSS VPW NCH W=2.12u L=0.06u
MNA106 NS S VSS VPW NCH W=0.7u L=0.06u
MNOE NM BCLK N1 VPW NCH W=0.15u L=0.06u
MNOE016 NM NCLK NENMUX VPW NCH W=0.45u L=0.06u
MNOE024 NENMUX S0 NET0135 VPW NCH W=0.4u L=0.06u
MNOE032 S BCLK M VPW NCH W=0.58u L=0.06u
MNOE044 S NCLK N1_12 VPW NCH W=0.15u L=0.06u
MNOE048 NENMUX NSEL NET0139 VPW NCH W=0.4u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1012 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1022 NSEL S0 VDD VNW PCH W=0.34u L=0.06u
MPA1030 NET0135 D1 VDD VNW PCH W=0.7u L=0.06u
MPA1038 M NM VDD VNW PCH W=0.7u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPA1042 P1_14 NS VDD VNW PCH W=0.15u L=0.06u
MPA1054 NET0139 D0 VDD VNW PCH W=0.7u L=0.06u
MPA1058 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA108 NS S VDD VNW PCH W=1u L=0.06u
MPOEN NM NCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN018 NM BCLK NENMUX VNW PCH W=0.45u L=0.06u
MPOEN026 NENMUX NSEL NET0135 VNW PCH W=0.4u L=0.06u
MPOEN034 S NCLK M VNW PCH W=0.58u L=0.06u
MPOEN046 S BCLK P1_14 VNW PCH W=0.15u L=0.06u
MPOEN050 NENMUX S0 NET0139 VNW PCH W=0.4u L=0.06u
.ENDS	M2DFFQX4MA10TR

****
.SUBCKT M2SDFFQNX0P5MA10TR  VDD VSS VPW VNW QN   CK D0 D1 SE S0 SI
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 S VSS VPW NCH W=0.15u L=0.06u
MNA1020 NSEL S0 VSS VPW NCH W=0.15u L=0.06u
MNA1028 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1032 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1036 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 NM M VSS VPW NCH W=0.15u L=0.06u
MNA1044 NET147 NSEMUX VSS VPW NCH W=0.15u L=0.06u
MNA1048 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA1068 NET155 D1 VSS VPW NCH W=0.2u L=0.06u
MNA1072 NET151 D0 VSS VPW NCH W=0.2u L=0.06u
MNA1076 QN S VSS VPW NCH W=0.31u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NS NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET147 VPW NCH W=0.15u L=0.06u
MNOE024 NS BCLK NM VPW NCH W=0.15u L=0.06u
MNOE052 NSEMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE056 NSEMUX NSE NENMUX VPW NCH W=0.2u L=0.06u
MNOE060 NENMUX S0 NET155 VPW NCH W=0.2u L=0.06u
MNOE064 NENMUX NSEL NET151 VPW NCH W=0.2u L=0.06u
MPA1 S NS VDD VNW PCH W=0.3u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NSEL S0 VDD VNW PCH W=0.2u L=0.06u
MPA1030 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1034 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1038 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA104 P1 S VDD VNW PCH W=0.15u L=0.06u
MPA1042 NM M VDD VNW PCH W=0.22u L=0.06u
MPA1046 NET147 NSEMUX VDD VNW PCH W=0.15u L=0.06u
MPA1050 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1070 NET155 D1 VDD VNW PCH W=0.4u L=0.06u
MPA1074 NET151 D0 VDD VNW PCH W=0.4u L=0.06u
MPA1078 QN S VDD VNW PCH W=0.37u L=0.06u
MPOEN NS BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET147 VNW PCH W=0.15u L=0.06u
MPOEN026 NS NCLK NM VNW PCH W=0.15u L=0.06u
MPOEN054 NSEMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN058 NSEMUX SE NENMUX VNW PCH W=0.25u L=0.06u
MPOEN062 NENMUX NSEL NET155 VNW PCH W=0.25u L=0.06u
MPOEN066 NENMUX S0 NET151 VNW PCH W=0.25u L=0.06u
.ENDS	M2SDFFQNX0P5MA10TR

****
.SUBCKT M2SDFFQNX1MA10TR  VDD VSS VPW VNW QN   CK D0 D1 SE S0 SI
MNA1 S NS VSS VPW NCH W=0.2u L=0.06u
MNA102 N1 S VSS VPW NCH W=0.15u L=0.06u
MNA1020 NSEL S0 VSS VPW NCH W=0.26u L=0.06u
MNA1028 NET104 D1 VSS VPW NCH W=0.2u L=0.06u
MNA1036 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1048 NM M VSS VPW NCH W=0.28u L=0.06u
MNA1052 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET96 NSEMUX VSS VPW NCH W=0.32u L=0.06u
MNA1072 NET100 D0 VSS VPW NCH W=0.2u L=0.06u
MNA1076 QN S VSS VPW NCH W=0.58u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NS NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET96 VPW NCH W=0.28u L=0.06u
MNOE024 NENMUX S0 NET104 VPW NCH W=0.2u L=0.06u
MNOE032 NS BCLK NM VPW NCH W=0.28u L=0.06u
MNOE056 NSEMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE060 NSEMUX NSE NENMUX VPW NCH W=0.2u L=0.06u
MNOE068 NENMUX NSEL NET100 VPW NCH W=0.2u L=0.06u
MPA1 S NS VDD VNW PCH W=0.4u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NSEL S0 VDD VNW PCH W=0.34u L=0.06u
MPA1030 NET104 D1 VDD VNW PCH W=0.4u L=0.06u
MPA1038 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA104 P1 S VDD VNW PCH W=0.15u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1050 NM M VDD VNW PCH W=0.52u L=0.06u
MPA1054 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1066 NET96 NSEMUX VDD VNW PCH W=0.32u L=0.06u
MPA1074 NET100 D0 VDD VNW PCH W=0.4u L=0.06u
MPA1078 QN S VDD VNW PCH W=0.7u L=0.06u
MPOEN NS BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET96 VNW PCH W=0.28u L=0.06u
MPOEN026 NENMUX NSEL NET104 VNW PCH W=0.3u L=0.06u
MPOEN034 NS NCLK NM VNW PCH W=0.28u L=0.06u
MPOEN058 NSEMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN062 NSEMUX SE NENMUX VNW PCH W=0.3u L=0.06u
MPOEN070 NENMUX S0 NET100 VNW PCH W=0.3u L=0.06u
.ENDS	M2SDFFQNX1MA10TR

****
.SUBCKT M2SDFFQNX2MA10TR  VDD VSS VPW VNW QN   CK D0 D1 SE S0 SI
MNA1 S NS VSS VPW NCH W=0.46u L=0.06u
MNA102 N1 S VSS VPW NCH W=0.15u L=0.06u
MNA1020 NSEL S0 VSS VPW NCH W=0.25u L=0.06u
MNA1028 NET104 D1 VSS VPW NCH W=0.3u L=0.06u
MNA1036 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1048 NM M VSS VPW NCH W=0.4u L=0.06u
MNA1052 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET96 NSEMUX VSS VPW NCH W=0.4u L=0.06u
MNA1072 NET100 D0 VSS VPW NCH W=0.3u L=0.06u
MNA1076 QN S VSS VPW NCH W=1.16u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NS NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET96 VPW NCH W=0.4u L=0.06u
MNOE024 NENMUX S0 NET104 VPW NCH W=0.3u L=0.06u
MNOE032 NS BCLK NM VPW NCH W=0.4u L=0.06u
MNOE056 NSEMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE060 NSEMUX NSE NENMUX VPW NCH W=0.3u L=0.06u
MNOE068 NENMUX NSEL NET100 VPW NCH W=0.3u L=0.06u
MPA1 S NS VDD VNW PCH W=0.7u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NSEL S0 VDD VNW PCH W=0.32u L=0.06u
MPA1030 NET104 D1 VDD VNW PCH W=0.6u L=0.06u
MPA1038 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA104 P1 S VDD VNW PCH W=0.15u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1050 NM M VDD VNW PCH W=0.65u L=0.06u
MPA1054 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1066 NET96 NSEMUX VDD VNW PCH W=0.4u L=0.06u
MPA1074 NET100 D0 VDD VNW PCH W=0.6u L=0.06u
MPA1078 QN S VDD VNW PCH W=1.4u L=0.06u
MPOEN NS BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET96 VNW PCH W=0.4u L=0.06u
MPOEN026 NENMUX NSEL NET104 VNW PCH W=0.45u L=0.06u
MPOEN034 NS NCLK NM VNW PCH W=0.4u L=0.06u
MPOEN058 NSEMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN062 NSEMUX SE NENMUX VNW PCH W=0.45u L=0.06u
MPOEN070 NENMUX S0 NET100 VNW PCH W=0.45u L=0.06u
.ENDS	M2SDFFQNX2MA10TR

****
.SUBCKT M2SDFFQNX3MA10TR  VDD VSS VPW VNW QN   CK D0 D1 SE S0 SI
MNA1 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1012 N1 S VSS VPW NCH W=0.15u L=0.06u
MNA1020 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNA1028 NSEL S0 VSS VPW NCH W=0.25u L=0.06u
MNA1036 NET104 D1 VSS VPW NCH W=0.3u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1044 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1048 NM M VSS VPW NCH W=0.51u L=0.06u
MNA1052 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA1064 NET96 NSEMUX VSS VPW NCH W=0.45u L=0.06u
MNA1072 NET100 D0 VSS VPW NCH W=0.3u L=0.06u
MNA1076 QN S VSS VPW NCH W=1.74u L=0.06u
MNA108 S NS VSS VPW NCH W=0.47u L=0.06u
MNOE NS BCLK NM VPW NCH W=0.45u L=0.06u
MNOE016 NS NCLK N1 VPW NCH W=0.15u L=0.06u
MNOE024 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE032 NENMUX S0 NET104 VPW NCH W=0.3u L=0.06u
MNOE040 M NCLK NET96 VPW NCH W=0.45u L=0.06u
MNOE056 NSEMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE060 NSEMUX NSE NENMUX VPW NCH W=0.3u L=0.06u
MNOE068 NENMUX NSEL NET100 VPW NCH W=0.3u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1010 S NS VDD VNW PCH W=0.7u L=0.06u
MPA1014 P1 S VDD VNW PCH W=0.15u L=0.06u
MPA1022 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1030 NSEL S0 VDD VNW PCH W=0.32u L=0.06u
MPA1038 NET104 D1 VDD VNW PCH W=0.6u L=0.06u
MPA1046 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1050 NM M VDD VNW PCH W=0.77u L=0.06u
MPA1054 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA1066 NET96 NSEMUX VDD VNW PCH W=0.45u L=0.06u
MPA1074 NET100 D0 VDD VNW PCH W=0.6u L=0.06u
MPA1078 QN S VDD VNW PCH W=2.1u L=0.06u
MPOEN NS NCLK NM VNW PCH W=0.45u L=0.06u
MPOEN018 NS BCLK P1 VNW PCH W=0.15u L=0.06u
MPOEN026 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN034 NENMUX NSEL NET104 VNW PCH W=0.45u L=0.06u
MPOEN042 M BCLK NET96 VNW PCH W=0.45u L=0.06u
MPOEN058 NSEMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN062 NSEMUX SE NENMUX VNW PCH W=0.45u L=0.06u
MPOEN070 NENMUX S0 NET100 VNW PCH W=0.45u L=0.06u
.ENDS	M2SDFFQNX3MA10TR

****
.SUBCKT M2SDFFQX0P5MA10TR  VDD VSS VPW VNW Q   CK D0 D1 SE S0 SI
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NSEL S0 VSS VPW NCH W=0.15u L=0.06u
MNA1028 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1032 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1036 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1040 NM M VSS VPW NCH W=0.15u L=0.06u
MNA1044 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1052 NET144 NSEMUX VSS VPW NCH W=0.15u L=0.06u
MNA1056 Q NS VSS VPW NCH W=0.28u L=0.06u
MNA1072 NET0132 D1 VSS VPW NCH W=0.2u L=0.06u
MNA1076 NET0128 D0 VSS VPW NCH W=0.2u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.15u L=0.06u
MNOE024 NS BCLK NM VPW NCH W=0.15u L=0.06u
MNOE048 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE060 NSEMUX NSE NENMUX VPW NCH W=0.2u L=0.06u
MNOE064 NENMUX S0 NET0132 VPW NCH W=0.2u L=0.06u
MNOE068 NENMUX NSEL NET0128 VPW NCH W=0.2u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NSEL S0 VDD VNW PCH W=0.2u L=0.06u
MPA1030 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1034 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1038 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NM M VDD VNW PCH W=0.2u L=0.06u
MPA1046 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1054 NET144 NSEMUX VDD VNW PCH W=0.15u L=0.06u
MPA1058 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA1074 NET0132 D1 VDD VNW PCH W=0.4u L=0.06u
MPA1078 NET0128 D0 VDD VNW PCH W=0.4u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.15u L=0.06u
MPOEN026 NS NCLK NM VNW PCH W=0.15u L=0.06u
MPOEN050 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN062 NSEMUX SE NENMUX VNW PCH W=0.3u L=0.06u
MPOEN066 NENMUX NSEL NET0132 VNW PCH W=0.25u L=0.06u
MPOEN070 NENMUX S0 NET0128 VNW PCH W=0.25u L=0.06u
.ENDS	M2SDFFQX0P5MA10TR

****
.SUBCKT M2SDFFQX1MA10TR  VDD VSS VPW VNW Q   CK D0 D1 SE S0 SI
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NSEL S0 VSS VPW NCH W=0.27u L=0.06u
MNA1028 NET0135 D1 VSS VPW NCH W=0.22u L=0.06u
MNA1036 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1048 NM M VSS VPW NCH W=0.32u L=0.06u
MNA1052 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1060 NET144 NSEMUX VSS VPW NCH W=0.28u L=0.06u
MNA1064 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA1076 NET0139 D0 VSS VPW NCH W=0.22u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.28u L=0.06u
MNOE024 NENMUX S0 NET0135 VPW NCH W=0.22u L=0.06u
MNOE032 NS BCLK NM VPW NCH W=0.28u L=0.06u
MNOE056 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE068 NSEMUX NSE NENMUX VPW NCH W=0.22u L=0.06u
MNOE072 NENMUX NSEL NET0139 VPW NCH W=0.22u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NSEL S0 VDD VNW PCH W=0.36u L=0.06u
MPA1030 NET0135 D1 VDD VNW PCH W=0.44u L=0.06u
MPA1038 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1050 NM M VDD VNW PCH W=0.5u L=0.06u
MPA1054 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1062 NET144 NSEMUX VDD VNW PCH W=0.28u L=0.06u
MPA1066 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA1078 NET0139 D0 VDD VNW PCH W=0.44u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.28u L=0.06u
MPOEN026 NENMUX NSEL NET0135 VNW PCH W=0.33u L=0.06u
MPOEN034 NS NCLK NM VNW PCH W=0.28u L=0.06u
MPOEN058 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN070 NSEMUX SE NENMUX VNW PCH W=0.33u L=0.06u
MPOEN074 NENMUX S0 NET0139 VNW PCH W=0.33u L=0.06u
.ENDS	M2SDFFQX1MA10TR

****
.SUBCKT M2SDFFQX2MA10TR  VDD VSS VPW VNW Q   CK D0 D1 SE S0 SI
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NSEL S0 VSS VPW NCH W=0.25u L=0.06u
MNA1028 NET0135 D1 VSS VPW NCH W=0.3u L=0.06u
MNA1036 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1048 NM M VSS VPW NCH W=0.4u L=0.06u
MNA1052 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1060 NET144 NSEMUX VSS VPW NCH W=0.4u L=0.06u
MNA1064 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA1076 NET0139 D0 VSS VPW NCH W=0.3u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.4u L=0.06u
MNOE024 NENMUX S0 NET0135 VPW NCH W=0.3u L=0.06u
MNOE032 NS BCLK NM VPW NCH W=0.4u L=0.06u
MNOE056 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE068 NSEMUX NSE NENMUX VPW NCH W=0.3u L=0.06u
MNOE072 NENMUX NSEL NET0139 VPW NCH W=0.3u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NSEL S0 VDD VNW PCH W=0.32u L=0.06u
MPA1030 NET0135 D1 VDD VNW PCH W=0.6u L=0.06u
MPA1038 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1050 NM M VDD VNW PCH W=0.6u L=0.06u
MPA1054 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1062 NET144 NSEMUX VDD VNW PCH W=0.4u L=0.06u
MPA1066 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA1078 NET0139 D0 VDD VNW PCH W=0.6u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.4u L=0.06u
MPOEN026 NENMUX NSEL NET0135 VNW PCH W=0.45u L=0.06u
MPOEN034 NS NCLK NM VNW PCH W=0.4u L=0.06u
MPOEN058 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN070 NSEMUX SE NENMUX VNW PCH W=0.45u L=0.06u
MPOEN074 NENMUX S0 NET0139 VNW PCH W=0.45u L=0.06u
.ENDS	M2SDFFQX2MA10TR

****
.SUBCKT M2SDFFQX3MA10TR  VDD VSS VPW VNW Q   CK D0 D1 SE S0 SI
MNA1 S NS VSS VPW NCH W=0.15u L=0.06u
MNA102 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1020 NSEL S0 VSS VPW NCH W=0.25u L=0.06u
MNA1028 NET0135 D1 VSS VPW NCH W=0.3u L=0.06u
MNA1036 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1048 NM M VSS VPW NCH W=0.5u L=0.06u
MNA1052 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA1060 NET144 NSEMUX VSS VPW NCH W=0.45u L=0.06u
MNA1064 Q NS VSS VPW NCH W=1.59u L=0.06u
MNA1076 NET0139 D0 VSS VPW NCH W=0.3u L=0.06u
MNA108 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE012 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE016 M NCLK NET144 VPW NCH W=0.45u L=0.06u
MNOE024 NENMUX S0 NET0135 VPW NCH W=0.3u L=0.06u
MNOE032 NS BCLK NM VPW NCH W=0.45u L=0.06u
MNOE056 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE068 NSEMUX NSE NENMUX VPW NCH W=0.3u L=0.06u
MNOE072 NENMUX NSEL NET0139 VPW NCH W=0.3u L=0.06u
MPA1 S NS VDD VNW PCH W=0.15u L=0.06u
MPA1010 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1022 NSEL S0 VDD VNW PCH W=0.32u L=0.06u
MPA1030 NET0135 D1 VDD VNW PCH W=0.6u L=0.06u
MPA1038 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA104 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1050 NM M VDD VNW PCH W=0.7u L=0.06u
MPA1054 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1062 NET144 NSEMUX VDD VNW PCH W=0.45u L=0.06u
MPA1066 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1078 NET0139 D0 VDD VNW PCH W=0.6u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN014 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN018 M BCLK NET144 VNW PCH W=0.45u L=0.06u
MPOEN026 NENMUX NSEL NET0135 VNW PCH W=0.45u L=0.06u
MPOEN034 NS NCLK NM VNW PCH W=0.45u L=0.06u
MPOEN058 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN070 NSEMUX SE NENMUX VNW PCH W=0.45u L=0.06u
MPOEN074 NENMUX S0 NET0139 VNW PCH W=0.45u L=0.06u
.ENDS	M2SDFFQX3MA10TR

****
.SUBCKT M2SDFFQX4MA10TR  VDD VSS VPW VNW Q   CK D0 D1 SE S0 SI
MNA1 NCLK CK VSS VPW NCH W=0.29u L=0.06u
MNA1010 N1 SI VSS VPW NCH W=0.15u L=0.06u
MNA1016 N1_15 NM VSS VPW NCH W=0.15u L=0.06u
MNA102 BCLK NCLK VSS VPW NCH W=0.26u L=0.06u
MNA1028 NSEL S0 VSS VPW NCH W=0.25u L=0.06u
MNA1036 NET0135 D1 VSS VPW NCH W=0.3u L=0.06u
MNA1044 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1048 NM M VSS VPW NCH W=0.58u L=0.06u
MNA1052 N1_19 S VSS VPW NCH W=0.15u L=0.06u
MNA106 S NS VSS VPW NCH W=0.15u L=0.06u
MNA1060 NET144 NSEMUX VSS VPW NCH W=0.45u L=0.06u
MNA1072 NET0139 D0 VSS VPW NCH W=0.3u L=0.06u
MNA1076 Q NS VSS VPW NCH W=2.12u L=0.06u
MNOE NSEMUX SE N1 VPW NCH W=0.15u L=0.06u
MNOE020 M BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE024 M NCLK NET144 VPW NCH W=0.45u L=0.06u
MNOE032 NENMUX S0 NET0135 VPW NCH W=0.3u L=0.06u
MNOE040 NS BCLK NM VPW NCH W=0.58u L=0.06u
MNOE056 NS NCLK N1_19 VPW NCH W=0.15u L=0.06u
MNOE064 NSEMUX NSE NENMUX VPW NCH W=0.3u L=0.06u
MNOE068 NENMUX NSEL NET0139 VPW NCH W=0.3u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.36u L=0.06u
MPA1012 P1 SI VDD VNW PCH W=0.2u L=0.06u
MPA1018 P1_17 NM VDD VNW PCH W=0.15u L=0.06u
MPA1030 NSEL S0 VDD VNW PCH W=0.32u L=0.06u
MPA1038 NET0135 D1 VDD VNW PCH W=0.6u L=0.06u
MPA104 BCLK NCLK VDD VNW PCH W=0.52u L=0.06u
MPA1046 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1050 NM M VDD VNW PCH W=0.7u L=0.06u
MPA1054 P1_21 S VDD VNW PCH W=0.15u L=0.06u
MPA1062 NET144 NSEMUX VDD VNW PCH W=0.45u L=0.06u
MPA1074 NET0139 D0 VDD VNW PCH W=0.6u L=0.06u
MPA1078 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA108 S NS VDD VNW PCH W=0.15u L=0.06u
MPOEN NSEMUX NSE P1 VNW PCH W=0.2u L=0.06u
MPOEN022 M NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN026 M BCLK NET144 VNW PCH W=0.45u L=0.06u
MPOEN034 NENMUX NSEL NET0135 VNW PCH W=0.45u L=0.06u
MPOEN042 NS NCLK NM VNW PCH W=0.58u L=0.06u
MPOEN058 NS BCLK P1_21 VNW PCH W=0.15u L=0.06u
MPOEN066 NSEMUX SE NENMUX VNW PCH W=0.45u L=0.06u
MPOEN070 NENMUX S0 NET0139 VNW PCH W=0.45u L=0.06u
.ENDS	M2SDFFQX4MA10TR

****
.SUBCKT MX2X0P5BA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 NSEL S0 VSS VPW NCH W=0.245u L=0.06u
MNA1016 INT0 A N1_6 VPW NCH W=0.15u L=0.06u
MNA102 Y INT0 N1 VPW NCH W=0.29u L=0.06u
MNA108 INT1 B N1_4 VPW NCH W=0.15u L=0.06u
MNA2 N1 INT1 VSS VPW NCH W=0.29u L=0.06u
MNA2010 N1_4 S0 VSS VPW NCH W=0.15u L=0.06u
MNA2018 N1_6 NSEL VSS VPW NCH W=0.15u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.325u L=0.06u
MPA1012 INT1 B VDD VNW PCH W=0.185u L=0.06u
MPA1020 INT0 A VDD VNW PCH W=0.185u L=0.06u
MPA105 Y INT0 VDD VNW PCH W=0.35u L=0.06u
MPA2 Y INT1 VDD VNW PCH W=0.35u L=0.06u
MPA2014 INT1 S0 VDD VNW PCH W=0.185u L=0.06u
MPA2022 INT0 NSEL VDD VNW PCH W=0.185u L=0.06u
.ENDS	MX2X0P5BA10TR

****
.SUBCKT MX2X0P5MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 NSEL S0 VSS VPW NCH W=0.27u L=0.06u
MNA1010 INT A N1A VPW NCH W=0.255u L=0.06u
MNA102 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA2 N1A NSEL VSS VPW NCH W=0.255u L=0.06u
MNB1 INT B N1B VPW NCH W=0.255u L=0.06u
MNB2 N1B S0 VSS VPW NCH W=0.255u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.36u L=0.06u
MPA1013 INT A P1 VNW PCH W=0.385u L=0.06u
MPA104 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA2 INT NSEL P1 VNW PCH W=0.385u L=0.06u
MPB1 P1 B VDD VNW PCH W=0.385u L=0.06u
MPB2 P1 S0 VDD VNW PCH W=0.385u L=0.06u
.ENDS	MX2X0P5MA10TR

****
.SUBCKT MX2X0P7BA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 NSEL S0 VSS VPW NCH W=0.265u L=0.06u
MNA1016 INT0 A N1_6 VPW NCH W=0.185u L=0.06u
MNA102 Y INT0 N1 VPW NCH W=0.405u L=0.06u
MNA108 INT1 B N1_4 VPW NCH W=0.185u L=0.06u
MNA2 N1 INT1 VSS VPW NCH W=0.405u L=0.06u
MNA2010 N1_4 S0 VSS VPW NCH W=0.185u L=0.06u
MNA2018 N1_6 NSEL VSS VPW NCH W=0.185u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.35u L=0.06u
MPA1012 INT1 B VDD VNW PCH W=0.23u L=0.06u
MPA1020 INT0 A VDD VNW PCH W=0.23u L=0.06u
MPA105 Y INT0 VDD VNW PCH W=0.49u L=0.06u
MPA2 Y INT1 VDD VNW PCH W=0.49u L=0.06u
MPA2014 INT1 S0 VDD VNW PCH W=0.23u L=0.06u
MPA2022 INT0 NSEL VDD VNW PCH W=0.23u L=0.06u
.ENDS	MX2X0P7BA10TR

****
.SUBCKT MX2X0P7MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 NSEL S0 VSS VPW NCH W=0.3u L=0.06u
MNA1010 INT A N1A VPW NCH W=0.315u L=0.06u
MNA102 Y INT VSS VPW NCH W=0.37u L=0.06u
MNA2 N1A NSEL VSS VPW NCH W=0.315u L=0.06u
MNB1 INT B N1B VPW NCH W=0.315u L=0.06u
MNB2 N1B S0 VSS VPW NCH W=0.315u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.4u L=0.06u
MPA1013 INT A P1 VNW PCH W=0.47u L=0.06u
MPA104 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA2 INT NSEL P1 VNW PCH W=0.47u L=0.06u
MPB1 P1 B VDD VNW PCH W=0.47u L=0.06u
MPB2 P1 S0 VDD VNW PCH W=0.47u L=0.06u
.ENDS	MX2X0P7MA10TR

****
.SUBCKT MX2X1BA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 NSEL S0 VSS VPW NCH W=0.29u L=0.06u
MNA1016 INT0 A N1_6 VPW NCH W=0.245u L=0.06u
MNA102 Y INT0 N1 VPW NCH W=0.58u L=0.06u
MNA108 INT1 B N1_4 VPW NCH W=0.245u L=0.06u
MNA2 N1 INT1 VSS VPW NCH W=0.58u L=0.06u
MNA2010 N1_4 S0 VSS VPW NCH W=0.245u L=0.06u
MNA2018 N1_6 NSEL VSS VPW NCH W=0.245u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.385u L=0.06u
MPA1012 INT1 B VDD VNW PCH W=0.3u L=0.06u
MPA1020 INT0 A VDD VNW PCH W=0.3u L=0.06u
MPA105 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MPA2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MPA2014 INT1 S0 VDD VNW PCH W=0.3u L=0.06u
MPA2022 INT0 NSEL VDD VNW PCH W=0.3u L=0.06u
.ENDS	MX2X1BA10TR

****
.SUBCKT MX2X1MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 NSEL S0 VSS VPW NCH W=0.31u L=0.06u
MNA1010 INT A N1A VPW NCH W=0.4u L=0.06u
MNA102 Y INT VSS VPW NCH W=0.53u L=0.06u
MNA2 N1A NSEL VSS VPW NCH W=0.4u L=0.06u
MNB1 INT B N1B VPW NCH W=0.4u L=0.06u
MNB2 N1B S0 VSS VPW NCH W=0.4u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.46u L=0.06u
MPA1013 INT A P1 VNW PCH W=0.6u L=0.06u
MPA104 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA2 INT NSEL P1 VNW PCH W=0.6u L=0.06u
MPB1 P1 B VDD VNW PCH W=0.6u L=0.06u
MPB2 P1 S0 VDD VNW PCH W=0.6u L=0.06u
.ENDS	MX2X1MA10TR

****

****

****

****

****

****
.SUBCKT MX2X3MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 NSEL S0 VSS VPW NCH W=0.92u L=0.06u
MNA1010 INT A N1A VPW NCH W=1.08u L=0.06u
MNA102 Y INT VSS VPW NCH W=1.59u L=0.06u
MNA2 N1A NSEL VSS VPW NCH W=1.08u L=0.06u
MNB1 INT B N1B VPW NCH W=1.08u L=0.06u
MNB2 N1B S0 VSS VPW NCH W=1.08u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=1.22u L=0.06u
MPA1013 INT A P1 VNW PCH W=1.635u L=0.06u
MPA104 Y INT VDD VNW PCH W=2.1u L=0.06u
MPA2 INT NSEL P1 VNW PCH W=1.635u L=0.06u
MPB1 P1 B VDD VNW PCH W=1.635u L=0.06u
MPB2 P1 S0 VDD VNW PCH W=1.635u L=0.06u
.ENDS	MX2X3MA10TR

****

****
.SUBCKT MX2X4MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 NSEL S0 VSS VPW NCH W=1.06u L=0.06u
MNA1010 INT A N1A VPW NCH W=1.395u L=0.06u
MNA102 Y INT VSS VPW NCH W=2.12u L=0.06u
MNA2 N1A NSEL VSS VPW NCH W=1.395u L=0.06u
MNB1 INT B N1B VPW NCH W=1.395u L=0.06u
MNB2 N1B S0 VSS VPW NCH W=1.395u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=1.4u L=0.06u
MPA1013 INT A P1 VNW PCH W=2.1u L=0.06u
MPA104 Y INT VDD VNW PCH W=2.8u L=0.06u
MPA2 INT NSEL P1 VNW PCH W=2.1u L=0.06u
MPB1 P1 B VDD VNW PCH W=2.1u L=0.06u
MPB2 P1 S0 VDD VNW PCH W=2.1u L=0.06u
.ENDS	MX2X4MA10TR

****

****
.SUBCKT MX2X6MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 NSEL S0 VSS VPW NCH W=1.59u L=0.06u
MNA1010 INT A N1A VPW NCH W=2.15u L=0.06u
MNA102 Y INT VSS VPW NCH W=3.18u L=0.06u
MNA2 N1A NSEL VSS VPW NCH W=2.15u L=0.06u
MNB1 INT B N1B VPW NCH W=2.15u L=0.06u
MNB2 N1B S0 VSS VPW NCH W=2.15u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=2.1u L=0.06u
MPA1013 INT A P1 VNW PCH W=3.25u L=0.06u
MPA104 Y INT VDD VNW PCH W=4.2u L=0.06u
MPA2 INT NSEL P1 VNW PCH W=3.25u L=0.06u
MPB1 P1 B VDD VNW PCH W=3.25u L=0.06u
MPB2 P1 S0 VDD VNW PCH W=3.25u L=0.06u
.ENDS	MX2X6MA10TR

****

****
.SUBCKT MXIT2X0P5MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 INT0 A VSS VPW NCH W=0.235u L=0.06u
MNA1012 INT1 B VSS VPW NCH W=0.235u L=0.06u
MNA108 NSEL S0 VSS VPW NCH W=0.275u L=0.06u
MNOE Y NSEL INT0 VPW NCH W=0.235u L=0.06u
MNOE02 Y S0 INT1 VPW NCH W=0.235u L=0.06u
MPA1 INT0 A VDD VNW PCH W=0.35u L=0.06u
MPA1010 NSEL S0 VDD VNW PCH W=0.365u L=0.06u
MPA1014 INT1 B VDD VNW PCH W=0.35u L=0.06u
MPOEN Y S0 INT0 VNW PCH W=0.235u L=0.06u
MPOEN04 Y NSEL INT1 VNW PCH W=0.235u L=0.06u
.ENDS	MXIT2X0P5MA10TR

****
.SUBCKT MXIT2X0P7MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 INT0 A VSS VPW NCH W=0.33u L=0.06u
MNA1012 INT1 B VSS VPW NCH W=0.33u L=0.06u
MNA108 NSEL S0 VSS VPW NCH W=0.31u L=0.06u
MNOE Y NSEL INT0 VPW NCH W=0.33u L=0.06u
MNOE02 Y S0 INT1 VPW NCH W=0.33u L=0.06u
MPA1 INT0 A VDD VNW PCH W=0.49u L=0.06u
MPA1010 NSEL S0 VDD VNW PCH W=0.42u L=0.06u
MPA1014 INT1 B VDD VNW PCH W=0.49u L=0.06u
MPOEN Y S0 INT0 VNW PCH W=0.33u L=0.06u
MPOEN04 Y NSEL INT1 VNW PCH W=0.33u L=0.06u
.ENDS	MXIT2X0P7MA10TR

****
.SUBCKT MXIT2X1MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 INT0 A VSS VPW NCH W=0.47u L=0.06u
MNA1012 INT1 B VSS VPW NCH W=0.47u L=0.06u
MNA108 NSEL S0 VSS VPW NCH W=0.35u L=0.06u
MNOE Y NSEL INT0 VPW NCH W=0.47u L=0.06u
MNOE02 Y S0 INT1 VPW NCH W=0.47u L=0.06u
MPA1 INT0 A VDD VNW PCH W=0.7u L=0.06u
MPA1010 NSEL S0 VDD VNW PCH W=0.47u L=0.06u
MPA1014 INT1 B VDD VNW PCH W=0.7u L=0.06u
MPOEN Y S0 INT0 VNW PCH W=0.47u L=0.06u
MPOEN04 Y NSEL INT1 VNW PCH W=0.47u L=0.06u
.ENDS	MXIT2X1MA10TR

****
.SUBCKT MXIT2X1P4MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 INT0 A VSS VPW NCH W=0.66u L=0.06u
MNA1012 INT1 B VSS VPW NCH W=0.66u L=0.06u
MNA108 NSEL S0 VSS VPW NCH W=0.5u L=0.06u
MNOE Y NSEL INT0 VPW NCH W=0.66u L=0.06u
MNOE02 Y S0 INT1 VPW NCH W=0.66u L=0.06u
MPA1 INT0 A VDD VNW PCH W=0.98u L=0.06u
MPA1010 NSEL S0 VDD VNW PCH W=0.66u L=0.06u
MPA1014 INT1 B VDD VNW PCH W=0.98u L=0.06u
MPOEN Y S0 INT0 VNW PCH W=0.66u L=0.06u
MPOEN04 Y NSEL INT1 VNW PCH W=0.66u L=0.06u
.ENDS	MXIT2X1P4MA10TR

****
.SUBCKT MXIT2X2MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 INT0 A VSS VPW NCH W=0.94u L=0.06u
MNA1012 INT1 B VSS VPW NCH W=0.94u L=0.06u
MNA108 NSEL S0 VSS VPW NCH W=0.7u L=0.06u
MNOE Y NSEL INT0 VPW NCH W=0.94u L=0.06u
MNOE02 Y S0 INT1 VPW NCH W=0.94u L=0.06u
MPA1 INT0 A VDD VNW PCH W=1.4u L=0.06u
MPA1010 NSEL S0 VDD VNW PCH W=0.92u L=0.06u
MPA1014 INT1 B VDD VNW PCH W=1.4u L=0.06u
MPOEN Y S0 INT0 VNW PCH W=0.94u L=0.06u
MPOEN04 Y NSEL INT1 VNW PCH W=0.94u L=0.06u
.ENDS	MXIT2X2MA10TR

****
.SUBCKT MXIT2X3MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 INT0 A VSS VPW NCH W=1.41u L=0.06u
MNA1012 INT1 B VSS VPW NCH W=1.41u L=0.06u
MNA108 NSEL S0 VSS VPW NCH W=0.94u L=0.06u
MNOE Y NSEL INT0 VPW NCH W=1.41u L=0.06u
MNOE02 Y S0 INT1 VPW NCH W=1.41u L=0.06u
MPA1 INT0 A VDD VNW PCH W=2.1u L=0.06u
MPA1010 NSEL S0 VDD VNW PCH W=1.25u L=0.06u
MPA1014 INT1 B VDD VNW PCH W=2.1u L=0.06u
MPOEN Y S0 INT0 VNW PCH W=1.41u L=0.06u
MPOEN04 Y NSEL INT1 VNW PCH W=1.41u L=0.06u
.ENDS	MXIT2X3MA10TR

****
.SUBCKT MXIT2X4MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 INT0 A VSS VPW NCH W=1.88u L=0.06u
MNA1012 INT1 B VSS VPW NCH W=1.88u L=0.06u
MNA108 NSEL S0 VSS VPW NCH W=1.23u L=0.06u
MNOE Y NSEL INT0 VPW NCH W=1.88u L=0.06u
MNOE02 Y S0 INT1 VPW NCH W=1.88u L=0.06u
MPA1 INT0 A VDD VNW PCH W=2.8u L=0.06u
MPA1010 NSEL S0 VDD VNW PCH W=1.65u L=0.06u
MPA1014 INT1 B VDD VNW PCH W=2.8u L=0.06u
MPOEN Y S0 INT0 VNW PCH W=1.88u L=0.06u
MPOEN04 Y NSEL INT1 VNW PCH W=1.88u L=0.06u
.ENDS	MXIT2X4MA10TR

****
.SUBCKT MXIT4X0P5MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=0.29u L=0.06u
MNA1012 NIN0 A VSS VPW NCH W=0.155u L=0.06u
MNA1024 NIN2 C VSS VPW NCH W=0.155u L=0.06u
MNA1028 NIN3 D VSS VPW NCH W=0.155u L=0.06u
MNA1032 NSEL1 S1 VSS VPW NCH W=0.2u L=0.06u
MNA1036 NSEL0 S0 VSS VPW NCH W=0.335u L=0.06u
MNA104 BIN01 NIN01 VSS VPW NCH W=0.155u L=0.06u
MNA1044 NIN1 B VSS VPW NCH W=0.155u L=0.06u
MNA1052 BIN23 NIN23 VSS VPW NCH W=0.155u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.155u L=0.06u
MNOE016 NIN23 NSEL0 NIN2 VPW NCH W=0.155u L=0.06u
MNOE020 NIN23 S0 NIN3 VPW NCH W=0.155u L=0.06u
MNOE040 NOUT NSEL1 BIN01 VPW NCH W=0.155u L=0.06u
MNOE048 NOUT S1 BIN23 VPW NCH W=0.155u L=0.06u
MNOE08 NIN01 S0 NIN1 VPW NCH W=0.155u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.35u L=0.06u
MPA1014 NIN0 A VDD VNW PCH W=0.26u L=0.06u
MPA1026 NIN2 C VDD VNW PCH W=0.26u L=0.06u
MPA1030 NIN3 D VDD VNW PCH W=0.26u L=0.06u
MPA1034 NSEL1 S1 VDD VNW PCH W=0.255u L=0.06u
MPA1038 NSEL0 S0 VDD VNW PCH W=0.425u L=0.06u
MPA1046 NIN1 B VDD VNW PCH W=0.26u L=0.06u
MPA1054 BIN23 NIN23 VDD VNW PCH W=0.19u L=0.06u
MPA106 BIN01 NIN01 VDD VNW PCH W=0.19u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.155u L=0.06u
MPOEN010 NIN01 NSEL0 NIN1 VNW PCH W=0.155u L=0.06u
MPOEN018 NIN23 S0 NIN2 VNW PCH W=0.155u L=0.06u
MPOEN022 NIN23 NSEL0 NIN3 VNW PCH W=0.155u L=0.06u
MPOEN042 NOUT S1 BIN01 VNW PCH W=0.155u L=0.06u
MPOEN050 NOUT NSEL1 BIN23 VNW PCH W=0.155u L=0.06u
.ENDS	MXIT4X0P5MA10TR

****
.SUBCKT MXIT4X0P7MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=0.41u L=0.06u
MNA1012 NIN0 A VSS VPW NCH W=0.195u L=0.06u
MNA1024 NIN2 C VSS VPW NCH W=0.195u L=0.06u
MNA1028 NIN3 D VSS VPW NCH W=0.195u L=0.06u
MNA1032 NSEL1 S1 VSS VPW NCH W=0.22u L=0.06u
MNA1036 NSEL0 S0 VSS VPW NCH W=0.37u L=0.06u
MNA104 BIN01 NIN01 VSS VPW NCH W=0.195u L=0.06u
MNA1044 NIN1 B VSS VPW NCH W=0.195u L=0.06u
MNA1052 BIN23 NIN23 VSS VPW NCH W=0.195u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.195u L=0.06u
MNOE016 NIN23 NSEL0 NIN2 VPW NCH W=0.195u L=0.06u
MNOE020 NIN23 S0 NIN3 VPW NCH W=0.195u L=0.06u
MNOE040 NOUT NSEL1 BIN01 VPW NCH W=0.195u L=0.06u
MNOE048 NOUT S1 BIN23 VPW NCH W=0.195u L=0.06u
MNOE08 NIN01 S0 NIN1 VPW NCH W=0.195u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.49u L=0.06u
MPA1014 NIN0 A VDD VNW PCH W=0.33u L=0.06u
MPA1026 NIN2 C VDD VNW PCH W=0.33u L=0.06u
MPA1030 NIN3 D VDD VNW PCH W=0.33u L=0.06u
MPA1034 NSEL1 S1 VDD VNW PCH W=0.275u L=0.06u
MPA1038 NSEL0 S0 VDD VNW PCH W=0.47u L=0.06u
MPA1046 NIN1 B VDD VNW PCH W=0.33u L=0.06u
MPA1054 BIN23 NIN23 VDD VNW PCH W=0.235u L=0.06u
MPA106 BIN01 NIN01 VDD VNW PCH W=0.235u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.195u L=0.06u
MPOEN010 NIN01 NSEL0 NIN1 VNW PCH W=0.195u L=0.06u
MPOEN018 NIN23 S0 NIN2 VNW PCH W=0.195u L=0.06u
MPOEN022 NIN23 NSEL0 NIN3 VNW PCH W=0.195u L=0.06u
MPOEN042 NOUT S1 BIN01 VNW PCH W=0.195u L=0.06u
MPOEN050 NOUT NSEL1 BIN23 VNW PCH W=0.195u L=0.06u
.ENDS	MXIT4X0P7MA10TR

****
.SUBCKT MXIT4X1MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=0.58u L=0.06u
MNA1012 NIN0 A VSS VPW NCH W=0.25u L=0.06u
MNA1024 NIN2 C VSS VPW NCH W=0.25u L=0.06u
MNA1028 NIN3 D VSS VPW NCH W=0.25u L=0.06u
MNA1032 NSEL1 S1 VSS VPW NCH W=0.26u L=0.06u
MNA1036 NSEL0 S0 VSS VPW NCH W=0.42u L=0.06u
MNA104 BIN01 NIN01 VSS VPW NCH W=0.25u L=0.06u
MNA1044 NIN1 B VSS VPW NCH W=0.25u L=0.06u
MNA1052 BIN23 NIN23 VSS VPW NCH W=0.25u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.25u L=0.06u
MNOE016 NIN23 NSEL0 NIN2 VPW NCH W=0.25u L=0.06u
MNOE020 NIN23 S0 NIN3 VPW NCH W=0.25u L=0.06u
MNOE040 NOUT NSEL1 BIN01 VPW NCH W=0.25u L=0.06u
MNOE048 NOUT S1 BIN23 VPW NCH W=0.25u L=0.06u
MNOE08 NIN01 S0 NIN1 VPW NCH W=0.25u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.7u L=0.06u
MPA1014 NIN0 A VDD VNW PCH W=0.42u L=0.06u
MPA1026 NIN2 C VDD VNW PCH W=0.42u L=0.06u
MPA1030 NIN3 D VDD VNW PCH W=0.42u L=0.06u
MPA1034 NSEL1 S1 VDD VNW PCH W=0.33u L=0.06u
MPA1038 NSEL0 S0 VDD VNW PCH W=0.53u L=0.06u
MPA1046 NIN1 B VDD VNW PCH W=0.42u L=0.06u
MPA1054 BIN23 NIN23 VDD VNW PCH W=0.3u L=0.06u
MPA106 BIN01 NIN01 VDD VNW PCH W=0.3u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.25u L=0.06u
MPOEN010 NIN01 NSEL0 NIN1 VNW PCH W=0.25u L=0.06u
MPOEN018 NIN23 S0 NIN2 VNW PCH W=0.25u L=0.06u
MPOEN022 NIN23 NSEL0 NIN3 VNW PCH W=0.25u L=0.06u
MPOEN042 NOUT S1 BIN01 VNW PCH W=0.25u L=0.06u
MPOEN050 NOUT NSEL1 BIN23 VNW PCH W=0.25u L=0.06u
.ENDS	MXIT4X1MA10TR

****
.SUBCKT MXIT4X1P4MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=0.81u L=0.06u
MNA1012 NIN0 A VSS VPW NCH W=0.32u L=0.06u
MNA1024 NIN2 C VSS VPW NCH W=0.32u L=0.06u
MNA1028 NIN3 D VSS VPW NCH W=0.32u L=0.06u
MNA1032 NSEL1 S1 VSS VPW NCH W=0.315u L=0.06u
MNA1036 NSEL0 S0 VSS VPW NCH W=0.5u L=0.06u
MNA104 BIN01 NIN01 VSS VPW NCH W=0.32u L=0.06u
MNA1044 NIN1 B VSS VPW NCH W=0.32u L=0.06u
MNA1052 BIN23 NIN23 VSS VPW NCH W=0.32u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.32u L=0.06u
MNOE016 NIN23 NSEL0 NIN2 VPW NCH W=0.32u L=0.06u
MNOE020 NIN23 S0 NIN3 VPW NCH W=0.32u L=0.06u
MNOE040 NOUT NSEL1 BIN01 VPW NCH W=0.32u L=0.06u
MNOE048 NOUT S1 BIN23 VPW NCH W=0.32u L=0.06u
MNOE08 NIN01 S0 NIN1 VPW NCH W=0.32u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.98u L=0.06u
MPA1014 NIN0 A VDD VNW PCH W=0.535u L=0.06u
MPA1026 NIN2 C VDD VNW PCH W=0.535u L=0.06u
MPA1030 NIN3 D VDD VNW PCH W=0.535u L=0.06u
MPA1034 NSEL1 S1 VDD VNW PCH W=0.405u L=0.06u
MPA1038 NSEL0 S0 VDD VNW PCH W=0.64u L=0.06u
MPA1046 NIN1 B VDD VNW PCH W=0.535u L=0.06u
MPA1054 BIN23 NIN23 VDD VNW PCH W=0.38u L=0.06u
MPA106 BIN01 NIN01 VDD VNW PCH W=0.38u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.32u L=0.06u
MPOEN010 NIN01 NSEL0 NIN1 VNW PCH W=0.32u L=0.06u
MPOEN018 NIN23 S0 NIN2 VNW PCH W=0.32u L=0.06u
MPOEN022 NIN23 NSEL0 NIN3 VNW PCH W=0.32u L=0.06u
MPOEN042 NOUT S1 BIN01 VNW PCH W=0.32u L=0.06u
MPOEN050 NOUT NSEL1 BIN23 VNW PCH W=0.32u L=0.06u
.ENDS	MXIT4X1P4MA10TR

****
.SUBCKT MXIT4X2MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=1.16u L=0.06u
MNA1012 NIN0 A VSS VPW NCH W=0.36u L=0.06u
MNA1024 NIN2 C VSS VPW NCH W=0.36u L=0.06u
MNA1028 NIN3 D VSS VPW NCH W=0.36u L=0.06u
MNA1032 NSEL1 S1 VSS VPW NCH W=0.365u L=0.06u
MNA1036 NSEL0 S0 VSS VPW NCH W=0.54u L=0.06u
MNA104 BIN01 NIN01 VSS VPW NCH W=0.36u L=0.06u
MNA1044 NIN1 B VSS VPW NCH W=0.36u L=0.06u
MNA1052 BIN23 NIN23 VSS VPW NCH W=0.36u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.36u L=0.06u
MNOE016 NIN23 NSEL0 NIN2 VPW NCH W=0.36u L=0.06u
MNOE020 NIN23 S0 NIN3 VPW NCH W=0.36u L=0.06u
MNOE040 NOUT NSEL1 BIN01 VPW NCH W=0.36u L=0.06u
MNOE048 NOUT S1 BIN23 VPW NCH W=0.36u L=0.06u
MNOE08 NIN01 S0 NIN1 VPW NCH W=0.36u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=1.4u L=0.06u
MPA1014 NIN0 A VDD VNW PCH W=0.61u L=0.06u
MPA1026 NIN2 C VDD VNW PCH W=0.61u L=0.06u
MPA1030 NIN3 D VDD VNW PCH W=0.61u L=0.06u
MPA1034 NSEL1 S1 VDD VNW PCH W=0.465u L=0.06u
MPA1038 NSEL0 S0 VDD VNW PCH W=0.68u L=0.06u
MPA1046 NIN1 B VDD VNW PCH W=0.61u L=0.06u
MPA1054 BIN23 NIN23 VDD VNW PCH W=0.43u L=0.06u
MPA106 BIN01 NIN01 VDD VNW PCH W=0.43u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.36u L=0.06u
MPOEN010 NIN01 NSEL0 NIN1 VNW PCH W=0.36u L=0.06u
MPOEN018 NIN23 S0 NIN2 VNW PCH W=0.36u L=0.06u
MPOEN022 NIN23 NSEL0 NIN3 VNW PCH W=0.36u L=0.06u
MPOEN042 NOUT S1 BIN01 VNW PCH W=0.36u L=0.06u
MPOEN050 NOUT NSEL1 BIN23 VNW PCH W=0.36u L=0.06u
.ENDS	MXIT4X2MA10TR

****
.SUBCKT MXIT4X3MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=1.74u L=0.06u
MNA1012 NIN0 A VSS VPW NCH W=0.42u L=0.06u
MNA1024 NIN2 C VSS VPW NCH W=0.42u L=0.06u
MNA1028 NIN3 D VSS VPW NCH W=0.42u L=0.06u
MNA1032 NSEL1 S1 VSS VPW NCH W=0.47u L=0.06u
MNA1036 NSEL0 S0 VSS VPW NCH W=0.65u L=0.06u
MNA104 BIN01 NIN01 VSS VPW NCH W=0.42u L=0.06u
MNA1044 NIN1 B VSS VPW NCH W=0.42u L=0.06u
MNA1052 BIN23 NIN23 VSS VPW NCH W=0.42u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.42u L=0.06u
MNOE016 NIN23 NSEL0 NIN2 VPW NCH W=0.42u L=0.06u
MNOE020 NIN23 S0 NIN3 VPW NCH W=0.42u L=0.06u
MNOE040 NOUT NSEL1 BIN01 VPW NCH W=0.42u L=0.06u
MNOE048 NOUT S1 BIN23 VPW NCH W=0.42u L=0.06u
MNOE08 NIN01 S0 NIN1 VPW NCH W=0.42u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=2.1u L=0.06u
MPA1014 NIN0 A VDD VNW PCH W=0.7u L=0.06u
MPA1026 NIN2 C VDD VNW PCH W=0.7u L=0.06u
MPA1030 NIN3 D VDD VNW PCH W=0.7u L=0.06u
MPA1034 NSEL1 S1 VDD VNW PCH W=0.595u L=0.06u
MPA1038 NSEL0 S0 VDD VNW PCH W=0.94u L=0.06u
MPA1046 NIN1 B VDD VNW PCH W=0.7u L=0.06u
MPA1054 BIN23 NIN23 VDD VNW PCH W=0.505u L=0.06u
MPA106 BIN01 NIN01 VDD VNW PCH W=0.505u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.42u L=0.06u
MPOEN010 NIN01 NSEL0 NIN1 VNW PCH W=0.42u L=0.06u
MPOEN018 NIN23 S0 NIN2 VNW PCH W=0.42u L=0.06u
MPOEN022 NIN23 NSEL0 NIN3 VNW PCH W=0.42u L=0.06u
MPOEN042 NOUT S1 BIN01 VNW PCH W=0.42u L=0.06u
MPOEN050 NOUT NSEL1 BIN23 VNW PCH W=0.42u L=0.06u
.ENDS	MXIT4X3MA10TR

****
.SUBCKT MXT2X0P5MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 Y NOUT VSS VPW NCH W=0.29u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.21u L=0.06u
MNA1016 INT1 B VSS VPW NCH W=0.2u L=0.06u
MNA108 INT0 A VSS VPW NCH W=0.2u L=0.06u
MNOE NOUT NSEL INT0 VPW NCH W=0.2u L=0.06u
MNOE04 NOUT S0 INT1 VPW NCH W=0.2u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.35u L=0.06u
MPA1010 INT0 A VDD VNW PCH W=0.29u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.31u L=0.06u
MPA1018 INT1 B VDD VNW PCH W=0.29u L=0.06u
MPOEN NOUT S0 INT0 VNW PCH W=0.2u L=0.06u
MPOEN06 NOUT NSEL INT1 VNW PCH W=0.2u L=0.06u
.ENDS	MXT2X0P5MA10TR

****
.SUBCKT MXT2X0P7MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 Y NOUT VSS VPW NCH W=0.405u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.235u L=0.06u
MNA1016 INT1 B VSS VPW NCH W=0.25u L=0.06u
MNA108 INT0 A VSS VPW NCH W=0.25u L=0.06u
MNOE NOUT NSEL INT0 VPW NCH W=0.25u L=0.06u
MNOE04 NOUT S0 INT1 VPW NCH W=0.25u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.49u L=0.06u
MPA1010 INT0 A VDD VNW PCH W=0.35u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.35u L=0.06u
MPA1018 INT1 B VDD VNW PCH W=0.35u L=0.06u
MPOEN NOUT S0 INT0 VNW PCH W=0.25u L=0.06u
MPOEN06 NOUT NSEL INT1 VNW PCH W=0.25u L=0.06u
.ENDS	MXT2X0P7MA10TR

****
.SUBCKT MXT2X1MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 Y NOUT VSS VPW NCH W=0.58u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.26u L=0.06u
MNA1016 INT1 B VSS VPW NCH W=0.32u L=0.06u
MNA108 INT0 A VSS VPW NCH W=0.32u L=0.06u
MNOE NOUT NSEL INT0 VPW NCH W=0.32u L=0.06u
MNOE04 NOUT S0 INT1 VPW NCH W=0.32u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.7u L=0.06u
MPA1010 INT0 A VDD VNW PCH W=0.45u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.4u L=0.06u
MPA1018 INT1 B VDD VNW PCH W=0.45u L=0.06u
MPOEN NOUT S0 INT0 VNW PCH W=0.32u L=0.06u
MPOEN06 NOUT NSEL INT1 VNW PCH W=0.32u L=0.06u
.ENDS	MXT2X1MA10TR

****
.SUBCKT MXT2X1P4MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 Y NOUT VSS VPW NCH W=0.81u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.28u L=0.06u
MNA1016 INT1 B VSS VPW NCH W=0.36u L=0.06u
MNA108 INT0 A VSS VPW NCH W=0.36u L=0.06u
MNOE NOUT NSEL INT0 VPW NCH W=0.36u L=0.06u
MNOE04 NOUT S0 INT1 VPW NCH W=0.36u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.98u L=0.06u
MPA1010 INT0 A VDD VNW PCH W=0.51u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.38u L=0.06u
MPA1018 INT1 B VDD VNW PCH W=0.51u L=0.06u
MPOEN NOUT S0 INT0 VNW PCH W=0.36u L=0.06u
MPOEN06 NOUT NSEL INT1 VNW PCH W=0.36u L=0.06u
.ENDS	MXT2X1P4MA10TR

****
.SUBCKT MXT2X2MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 Y NOUT VSS VPW NCH W=1.16u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.35u L=0.06u
MNA1016 INT1 B VSS VPW NCH W=0.47u L=0.06u
MNA108 INT0 A VSS VPW NCH W=0.47u L=0.06u
MNOE NOUT NSEL INT0 VPW NCH W=0.47u L=0.06u
MNOE04 NOUT S0 INT1 VPW NCH W=0.47u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=1.4u L=0.06u
MPA1010 INT0 A VDD VNW PCH W=0.7u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.47u L=0.06u
MPA1018 INT1 B VDD VNW PCH W=0.7u L=0.06u
MPOEN NOUT S0 INT0 VNW PCH W=0.47u L=0.06u
MPOEN06 NOUT NSEL INT1 VNW PCH W=0.47u L=0.06u
.ENDS	MXT2X2MA10TR

****
.SUBCKT MXT2X3MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 Y NOUT VSS VPW NCH W=1.74u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.5u L=0.06u
MNA1016 INT1 B VSS VPW NCH W=0.74u L=0.06u
MNA108 INT0 A VSS VPW NCH W=0.74u L=0.06u
MNOE NOUT NSEL INT0 VPW NCH W=0.74u L=0.06u
MNOE04 NOUT S0 INT1 VPW NCH W=0.74u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=2.1u L=0.06u
MPA1010 INT0 A VDD VNW PCH W=1.04u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.74u L=0.06u
MPA1018 INT1 B VDD VNW PCH W=1.04u L=0.06u
MPOEN NOUT S0 INT0 VNW PCH W=0.74u L=0.06u
MPOEN06 NOUT NSEL INT1 VNW PCH W=0.74u L=0.06u
.ENDS	MXT2X3MA10TR

****
.SUBCKT MXT2X4MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 Y NOUT VSS VPW NCH W=2.32u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.64u L=0.06u
MNA1016 INT1 B VSS VPW NCH W=0.94u L=0.06u
MNA108 INT0 A VSS VPW NCH W=0.94u L=0.06u
MNOE NOUT NSEL INT0 VPW NCH W=0.94u L=0.06u
MNOE04 NOUT S0 INT1 VPW NCH W=0.94u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=2.8u L=0.06u
MPA1010 INT0 A VDD VNW PCH W=1.32u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=0.95u L=0.06u
MPA1018 INT1 B VDD VNW PCH W=1.32u L=0.06u
MPOEN NOUT S0 INT0 VNW PCH W=0.94u L=0.06u
MPOEN06 NOUT NSEL INT1 VNW PCH W=0.94u L=0.06u
.ENDS	MXT2X4MA10TR

****
.SUBCKT MXT2X6MA10TR  VDD VSS VPW VNW Y   A B S0
MNA1 Y NOUT VSS VPW NCH W=3.48u L=0.06u
MNA1012 NSEL S0 VSS VPW NCH W=0.92u L=0.06u
MNA1016 INT1 B VSS VPW NCH W=1.41u L=0.06u
MNA108 INT0 A VSS VPW NCH W=1.41u L=0.06u
MNOE NOUT NSEL INT0 VPW NCH W=1.41u L=0.06u
MNOE04 NOUT S0 INT1 VPW NCH W=1.41u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=4.2u L=0.06u
MPA1010 INT0 A VDD VNW PCH W=2.01u L=0.06u
MPA1014 NSEL S0 VDD VNW PCH W=1.38u L=0.06u
MPA1018 INT1 B VDD VNW PCH W=2.01u L=0.06u
MPOEN NOUT S0 INT0 VNW PCH W=1.41u L=0.06u
MPOEN06 NOUT NSEL INT1 VNW PCH W=1.41u L=0.06u
.ENDS	MXT2X6MA10TR

****
.SUBCKT MXT4X0P5MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=0.29u L=0.06u
MNA1020 NIN2 C VSS VPW NCH W=0.2u L=0.06u
MNA1024 NIN3 D VSS VPW NCH W=0.2u L=0.06u
MNA1028 NSEL1 S1 VSS VPW NCH W=0.205u L=0.06u
MNA1032 NSEL0 S0 VSS VPW NCH W=0.35u L=0.06u
MNA1040 NIN1 B VSS VPW NCH W=0.2u L=0.06u
MNA108 NIN0 A VSS VPW NCH W=0.2u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.2u L=0.06u
MNOE012 NIN23 NSEL0 NIN2 VPW NCH W=0.2u L=0.06u
MNOE016 NIN23 S0 NIN3 VPW NCH W=0.2u L=0.06u
MNOE036 NOUT NSEL1 NIN01 VPW NCH W=0.2u L=0.06u
MNOE04 NIN01 S0 NIN1 VPW NCH W=0.2u L=0.06u
MNOE044 NOUT S1 NIN23 VPW NCH W=0.2u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.35u L=0.06u
MPA1010 NIN0 A VDD VNW PCH W=0.335u L=0.06u
MPA1022 NIN2 C VDD VNW PCH W=0.335u L=0.06u
MPA1026 NIN3 D VDD VNW PCH W=0.335u L=0.06u
MPA1030 NSEL1 S1 VDD VNW PCH W=0.295u L=0.06u
MPA1034 NSEL0 S0 VDD VNW PCH W=0.5u L=0.06u
MPA1042 NIN1 B VDD VNW PCH W=0.335u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.2u L=0.06u
MPOEN014 NIN23 S0 NIN2 VNW PCH W=0.2u L=0.06u
MPOEN018 NIN23 NSEL0 NIN3 VNW PCH W=0.2u L=0.06u
MPOEN038 NOUT S1 NIN01 VNW PCH W=0.2u L=0.06u
MPOEN046 NOUT NSEL1 NIN23 VNW PCH W=0.2u L=0.06u
MPOEN06 NIN01 NSEL0 NIN1 VNW PCH W=0.2u L=0.06u
.ENDS	MXT4X0P5MA10TR

****
.SUBCKT MXT4X0P7MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=0.41u L=0.06u
MNA1020 NIN2 C VSS VPW NCH W=0.26u L=0.06u
MNA1024 NIN3 D VSS VPW NCH W=0.26u L=0.06u
MNA1028 NSEL1 S1 VSS VPW NCH W=0.235u L=0.06u
MNA1032 NSEL0 S0 VSS VPW NCH W=0.395u L=0.06u
MNA1040 NIN1 B VSS VPW NCH W=0.26u L=0.06u
MNA108 NIN0 A VSS VPW NCH W=0.26u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.26u L=0.06u
MNOE012 NIN23 NSEL0 NIN2 VPW NCH W=0.26u L=0.06u
MNOE016 NIN23 S0 NIN3 VPW NCH W=0.26u L=0.06u
MNOE036 NOUT NSEL1 NIN01 VPW NCH W=0.26u L=0.06u
MNOE04 NIN01 S0 NIN1 VPW NCH W=0.26u L=0.06u
MNOE044 NOUT S1 NIN23 VPW NCH W=0.26u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.49u L=0.06u
MPA1010 NIN0 A VDD VNW PCH W=0.435u L=0.06u
MPA1022 NIN2 C VDD VNW PCH W=0.435u L=0.06u
MPA1026 NIN3 D VDD VNW PCH W=0.435u L=0.06u
MPA1030 NSEL1 S1 VDD VNW PCH W=0.345u L=0.06u
MPA1034 NSEL0 S0 VDD VNW PCH W=0.575u L=0.06u
MPA1042 NIN1 B VDD VNW PCH W=0.435u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.26u L=0.06u
MPOEN014 NIN23 S0 NIN2 VNW PCH W=0.26u L=0.06u
MPOEN018 NIN23 NSEL0 NIN3 VNW PCH W=0.26u L=0.06u
MPOEN038 NOUT S1 NIN01 VNW PCH W=0.26u L=0.06u
MPOEN046 NOUT NSEL1 NIN23 VNW PCH W=0.26u L=0.06u
MPOEN06 NIN01 NSEL0 NIN1 VNW PCH W=0.26u L=0.06u
.ENDS	MXT4X0P7MA10TR

****
.SUBCKT MXT4X1MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=0.58u L=0.06u
MNA1020 NIN2 C VSS VPW NCH W=0.32u L=0.06u
MNA1024 NIN3 D VSS VPW NCH W=0.32u L=0.06u
MNA1028 NSEL1 S1 VSS VPW NCH W=0.26u L=0.06u
MNA1032 NSEL0 S0 VSS VPW NCH W=0.455u L=0.06u
MNA1040 NIN1 B VSS VPW NCH W=0.32u L=0.06u
MNA108 NIN0 A VSS VPW NCH W=0.32u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.32u L=0.06u
MNOE012 NIN23 NSEL0 NIN2 VPW NCH W=0.32u L=0.06u
MNOE016 NIN23 S0 NIN3 VPW NCH W=0.32u L=0.06u
MNOE036 NOUT NSEL1 NIN01 VPW NCH W=0.32u L=0.06u
MNOE04 NIN01 S0 NIN1 VPW NCH W=0.32u L=0.06u
MNOE044 NOUT S1 NIN23 VPW NCH W=0.32u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.7u L=0.06u
MPA1010 NIN0 A VDD VNW PCH W=0.535u L=0.06u
MPA1022 NIN2 C VDD VNW PCH W=0.535u L=0.06u
MPA1026 NIN3 D VDD VNW PCH W=0.535u L=0.06u
MPA1030 NSEL1 S1 VDD VNW PCH W=0.36u L=0.06u
MPA1034 NSEL0 S0 VDD VNW PCH W=0.635u L=0.06u
MPA1042 NIN1 B VDD VNW PCH W=0.535u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.32u L=0.06u
MPOEN014 NIN23 S0 NIN2 VNW PCH W=0.32u L=0.06u
MPOEN018 NIN23 NSEL0 NIN3 VNW PCH W=0.32u L=0.06u
MPOEN038 NOUT S1 NIN01 VNW PCH W=0.32u L=0.06u
MPOEN046 NOUT NSEL1 NIN23 VNW PCH W=0.32u L=0.06u
MPOEN06 NIN01 NSEL0 NIN1 VNW PCH W=0.32u L=0.06u
.ENDS	MXT4X1MA10TR

****
.SUBCKT MXT4X1P4MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=0.81u L=0.06u
MNA1020 NIN2 C VSS VPW NCH W=0.37u L=0.06u
MNA1024 NIN3 D VSS VPW NCH W=0.37u L=0.06u
MNA1028 NSEL1 S1 VSS VPW NCH W=0.34u L=0.06u
MNA1032 NSEL0 S0 VSS VPW NCH W=0.58u L=0.06u
MNA1040 NIN1 B VSS VPW NCH W=0.37u L=0.06u
MNA108 NIN0 A VSS VPW NCH W=0.37u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.37u L=0.06u
MNOE012 NIN23 NSEL0 NIN2 VPW NCH W=0.37u L=0.06u
MNOE016 NIN23 S0 NIN3 VPW NCH W=0.37u L=0.06u
MNOE036 NOUT NSEL1 NIN01 VPW NCH W=0.37u L=0.06u
MNOE04 NIN01 S0 NIN1 VPW NCH W=0.37u L=0.06u
MNOE044 NOUT S1 NIN23 VPW NCH W=0.37u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=0.98u L=0.06u
MPA1010 NIN0 A VDD VNW PCH W=0.55u L=0.06u
MPA1022 NIN2 C VDD VNW PCH W=0.55u L=0.06u
MPA1026 NIN3 D VDD VNW PCH W=0.55u L=0.06u
MPA1030 NSEL1 S1 VDD VNW PCH W=0.48u L=0.06u
MPA1034 NSEL0 S0 VDD VNW PCH W=0.7u L=0.06u
MPA1042 NIN1 B VDD VNW PCH W=0.55u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.37u L=0.06u
MPOEN014 NIN23 S0 NIN2 VNW PCH W=0.37u L=0.06u
MPOEN018 NIN23 NSEL0 NIN3 VNW PCH W=0.37u L=0.06u
MPOEN038 NOUT S1 NIN01 VNW PCH W=0.37u L=0.06u
MPOEN046 NOUT NSEL1 NIN23 VNW PCH W=0.37u L=0.06u
MPOEN06 NIN01 NSEL0 NIN1 VNW PCH W=0.37u L=0.06u
.ENDS	MXT4X1P4MA10TR

****
.SUBCKT MXT4X2MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=1.16u L=0.06u
MNA1020 NIN2 C VSS VPW NCH W=0.42u L=0.06u
MNA1024 NIN3 D VSS VPW NCH W=0.42u L=0.06u
MNA1028 NSEL1 S1 VSS VPW NCH W=0.385u L=0.06u
MNA1032 NSEL0 S0 VSS VPW NCH W=0.52u L=0.06u
MNA1040 NIN1 B VSS VPW NCH W=0.42u L=0.06u
MNA108 NIN0 A VSS VPW NCH W=0.42u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.42u L=0.06u
MNOE012 NIN23 NSEL0 NIN2 VPW NCH W=0.42u L=0.06u
MNOE016 NIN23 S0 NIN3 VPW NCH W=0.42u L=0.06u
MNOE036 NOUT NSEL1 NIN01 VPW NCH W=0.42u L=0.06u
MNOE04 NIN01 S0 NIN1 VPW NCH W=0.42u L=0.06u
MNOE044 NOUT S1 NIN23 VPW NCH W=0.42u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=1.4u L=0.06u
MPA1010 NIN0 A VDD VNW PCH W=0.7u L=0.06u
MPA1022 NIN2 C VDD VNW PCH W=0.7u L=0.06u
MPA1026 NIN3 D VDD VNW PCH W=0.7u L=0.06u
MPA1030 NSEL1 S1 VDD VNW PCH W=0.535u L=0.06u
MPA1034 NSEL0 S0 VDD VNW PCH W=0.7u L=0.06u
MPA1042 NIN1 B VDD VNW PCH W=0.7u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.42u L=0.06u
MPOEN014 NIN23 S0 NIN2 VNW PCH W=0.42u L=0.06u
MPOEN018 NIN23 NSEL0 NIN3 VNW PCH W=0.42u L=0.06u
MPOEN038 NOUT S1 NIN01 VNW PCH W=0.42u L=0.06u
MPOEN046 NOUT NSEL1 NIN23 VNW PCH W=0.42u L=0.06u
MPOEN06 NIN01 NSEL0 NIN1 VNW PCH W=0.42u L=0.06u
.ENDS	MXT4X2MA10TR

****
.SUBCKT MXT4X3MA10TR  VDD VSS VPW VNW Y   A B C D S0 S1
MNA1 Y NOUT VSS VPW NCH W=1.74u L=0.06u
MNA1020 NIN2 C VSS VPW NCH W=0.82u L=0.06u
MNA1024 NIN3 D VSS VPW NCH W=0.82u L=0.06u
MNA1028 NSEL1 S1 VSS VPW NCH W=0.64u L=0.06u
MNA1032 NSEL0 S0 VSS VPW NCH W=1.08u L=0.06u
MNA1040 NIN1 B VSS VPW NCH W=0.82u L=0.06u
MNA108 NIN0 A VSS VPW NCH W=0.82u L=0.06u
MNOE NIN01 NSEL0 NIN0 VPW NCH W=0.82u L=0.06u
MNOE012 NIN23 NSEL0 NIN2 VPW NCH W=0.82u L=0.06u
MNOE016 NIN23 S0 NIN3 VPW NCH W=0.82u L=0.06u
MNOE036 NOUT NSEL1 NIN01 VPW NCH W=0.82u L=0.06u
MNOE04 NIN01 S0 NIN1 VPW NCH W=0.82u L=0.06u
MNOE044 NOUT S1 NIN23 VPW NCH W=0.82u L=0.06u
MPA1 Y NOUT VDD VNW PCH W=2.1u L=0.06u
MPA1010 NIN0 A VDD VNW PCH W=1.38u L=0.06u
MPA1022 NIN2 C VDD VNW PCH W=1.38u L=0.06u
MPA1026 NIN3 D VDD VNW PCH W=1.38u L=0.06u
MPA1030 NSEL1 S1 VDD VNW PCH W=0.88u L=0.06u
MPA1034 NSEL0 S0 VDD VNW PCH W=1.47u L=0.06u
MPA1042 NIN1 B VDD VNW PCH W=1.38u L=0.06u
MPOEN NIN01 S0 NIN0 VNW PCH W=0.82u L=0.06u
MPOEN014 NIN23 S0 NIN2 VNW PCH W=0.82u L=0.06u
MPOEN018 NIN23 NSEL0 NIN3 VNW PCH W=0.82u L=0.06u
MPOEN038 NOUT S1 NIN01 VNW PCH W=0.82u L=0.06u
MPOEN046 NOUT NSEL1 NIN23 VNW PCH W=0.82u L=0.06u
MPOEN06 NIN01 NSEL0 NIN1 VNW PCH W=0.82u L=0.06u
.ENDS	MXT4X3MA10TR

****
.SUBCKT NAND2BX0P5MA10TR  VDD VSS VPW VNW Y   AN B
MNA1 Y NET24 N1 VPW NCH W=0.29u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.29u L=0.06u
MPA1 Y NET24 VDD VNW PCH W=0.24u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.2u L=0.06u
MPA2 Y B VDD VNW PCH W=0.24u L=0.06u
.ENDS	NAND2BX0P5MA10TR

****
.SUBCKT NAND2BX0P7MA10TR  VDD VSS VPW VNW Y   AN B
MNA1 Y NET24 N1 VPW NCH W=0.41u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.41u L=0.06u
MPA1 Y NET24 VDD VNW PCH W=0.34u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.2u L=0.06u
MPA2 Y B VDD VNW PCH W=0.34u L=0.06u
.ENDS	NAND2BX0P7MA10TR

****
.SUBCKT NAND2BX1MA10TR  VDD VSS VPW VNW Y   AN B
MNA1 Y NET24 N1 VPW NCH W=0.58u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.58u L=0.06u
MPA1 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.2u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS	NAND2BX1MA10TR

****

****

****

****

****

****

****
.SUBCKT NAND2X0P5AA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A N1 VPW NCH W=0.29u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.29u L=0.06u
MPA1 Y A VDD VNW PCH W=0.295u L=0.06u
MPA2 Y B VDD VNW PCH W=0.295u L=0.06u
.ENDS	NAND2X0P5AA10TR

****
.SUBCKT NAND2X0P5BA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A N1 VPW NCH W=0.29u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.29u L=0.06u
MPA1 Y A VDD VNW PCH W=0.35u L=0.06u
MPA2 Y B VDD VNW PCH W=0.35u L=0.06u
.ENDS	NAND2X0P5BA10TR

****
.SUBCKT NAND2X0P5MA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A N1 VPW NCH W=0.29u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.29u L=0.06u
MPA1 Y A VDD VNW PCH W=0.24u L=0.06u
MPA2 Y B VDD VNW PCH W=0.24u L=0.06u
.ENDS	NAND2X0P5MA10TR

****
.SUBCKT NAND2X0P7AA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A N1 VPW NCH W=0.405u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.405u L=0.06u
MPA1 Y A VDD VNW PCH W=0.415u L=0.06u
MPA2 Y B VDD VNW PCH W=0.415u L=0.06u
.ENDS	NAND2X0P7AA10TR

****
.SUBCKT NAND2X0P7BA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A N1 VPW NCH W=0.405u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.405u L=0.06u
MPA1 Y A VDD VNW PCH W=0.49u L=0.06u
MPA2 Y B VDD VNW PCH W=0.49u L=0.06u
.ENDS	NAND2X0P7BA10TR

****
.SUBCKT NAND2X0P7MA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A N1 VPW NCH W=0.41u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.34u L=0.06u
MPA2 Y B VDD VNW PCH W=0.34u L=0.06u
.ENDS	NAND2X0P7MA10TR

****
.SUBCKT NAND2X1AA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A N1 VPW NCH W=0.58u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.59u L=0.06u
MPA2 Y B VDD VNW PCH W=0.59u L=0.06u
.ENDS	NAND2X1AA10TR

****
.SUBCKT NAND2X1BA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A N1 VPW NCH W=0.58u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.7u L=0.06u
MPA2 Y B VDD VNW PCH W=0.7u L=0.06u
.ENDS	NAND2X1BA10TR

****
.SUBCKT NAND2X1MA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A N1 VPW NCH W=0.58u L=0.06u
MNA2 N1 B VSS VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS	NAND2X1MA10TR

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****

****
.SUBCKT NAND2XBX0P5MA10TR  VDD VSS VPW VNW Y   A BN
MNA1 Y A N1 VPW NCH W=0.29u L=0.06u
MNA104 NET24 BN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1 NET24 VSS VPW NCH W=0.29u L=0.06u
MPA1 Y A VDD VNW PCH W=0.24u L=0.06u
MPA106 NET24 BN VDD VNW PCH W=0.2u L=0.06u
MPA2 Y NET24 VDD VNW PCH W=0.24u L=0.06u
.ENDS	NAND2XBX0P5MA10TR

****
.SUBCKT NAND2XBX0P7MA10TR  VDD VSS VPW VNW Y   A BN
MNA1 Y A N1 VPW NCH W=0.41u L=0.06u
MNA104 NET24 BN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1 NET24 VSS VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.34u L=0.06u
MPA106 NET24 BN VDD VNW PCH W=0.2u L=0.06u
MPA2 Y NET24 VDD VNW PCH W=0.34u L=0.06u
.ENDS	NAND2XBX0P7MA10TR

****
.SUBCKT NAND2XBX1MA10TR  VDD VSS VPW VNW Y   A BN
MNA1 Y A N1 VPW NCH W=0.58u L=0.06u
MNA104 NET24 BN VSS VPW NCH W=0.15u L=0.06u
MNA2 N1 NET24 VSS VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MPA106 NET24 BN VDD VNW PCH W=0.2u L=0.06u
MPA2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
.ENDS	NAND2XBX1MA10TR

****

****

****

****

****

****

****
.SUBCKT NAND3BX0P5MA10TR  VDD VSS VPW VNW Y   AN B C
MNA1 NET14 AN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET14 N2 VPW NCH W=0.29u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.29u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.29u L=0.06u
MPA1 NET14 AN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y NET14 VDD VNW PCH W=0.18u L=0.06u
MPA2 Y B VDD VNW PCH W=0.18u L=0.06u
MPA3 Y C VDD VNW PCH W=0.18u L=0.06u
.ENDS	NAND3BX0P5MA10TR

****
.SUBCKT NAND3BX0P7MA10TR  VDD VSS VPW VNW Y   AN B C
MNA1 NET14 AN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET14 N2 VPW NCH W=0.41u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.41u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.41u L=0.06u
MPA1 NET14 AN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y NET14 VDD VNW PCH W=0.25u L=0.06u
MPA2 Y B VDD VNW PCH W=0.25u L=0.06u
MPA3 Y C VDD VNW PCH W=0.25u L=0.06u
.ENDS	NAND3BX0P7MA10TR

****
.SUBCKT NAND3BX1MA10TR  VDD VSS VPW VNW Y   AN B C
MNA1 NET14 AN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET14 N2 VPW NCH W=0.58u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.58u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.58u L=0.06u
MPA1 NET14 AN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y NET14 VDD VNW PCH W=0.36u L=0.06u
MPA2 Y B VDD VNW PCH W=0.36u L=0.06u
MPA3 Y C VDD VNW PCH W=0.36u L=0.06u
.ENDS	NAND3BX1MA10TR

****

****

****
.SUBCKT NAND3BX3MA10TR  VDD VSS VPW VNW Y   AN B C
MNA1 NET14 AN VSS VPW NCH W=0.385u L=0.06u
MNA102 Y NET14 N2 VPW NCH W=1.74u L=0.06u
MNA2 N2 B N1 VPW NCH W=1.74u L=0.06u
MNA3 N1 C VSS VPW NCH W=1.74u L=0.06u
MPA1 NET14 AN VDD VNW PCH W=0.51u L=0.06u
MPA105 Y NET14 VDD VNW PCH W=1.08u L=0.06u
MPA2 Y B VDD VNW PCH W=1.08u L=0.06u
MPA3 Y C VDD VNW PCH W=1.08u L=0.06u
.ENDS	NAND3BX3MA10TR

****
.SUBCKT NAND3BX4MA10TR  VDD VSS VPW VNW Y   AN B C
MNA1 NET14 AN VSS VPW NCH W=0.5u L=0.06u
MNA102 Y NET14 N2 VPW NCH W=2.32u L=0.06u
MNA2 N2 B N1 VPW NCH W=2.32u L=0.06u
MNA3 N1 C VSS VPW NCH W=2.32u L=0.06u
MPA1 NET14 AN VDD VNW PCH W=0.66u L=0.06u
MPA105 Y NET14 VDD VNW PCH W=1.44u L=0.06u
MPA2 Y B VDD VNW PCH W=1.44u L=0.06u
MPA3 Y C VDD VNW PCH W=1.44u L=0.06u
.ENDS	NAND3BX4MA10TR

****
.SUBCKT NAND3BX6MA10TR  VDD VSS VPW VNW Y   AN B C
MNA1 NET14 AN VSS VPW NCH W=0.75u L=0.06u
MNA102 Y NET14 N2 VPW NCH W=3.48u L=0.06u
MNA2 N2 B N1 VPW NCH W=3.48u L=0.06u
MNA3 N1 C VSS VPW NCH W=3.48u L=0.06u
MPA1 NET14 AN VDD VNW PCH W=0.99u L=0.06u
MPA105 Y NET14 VDD VNW PCH W=2.16u L=0.06u
MPA2 Y B VDD VNW PCH W=2.16u L=0.06u
MPA3 Y C VDD VNW PCH W=2.16u L=0.06u
.ENDS	NAND3BX6MA10TR

****
.SUBCKT NAND3X0P5AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=0.29u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.29u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.29u L=0.06u
MPA1 Y A VDD VNW PCH W=0.27u L=0.06u
MPA2 Y B VDD VNW PCH W=0.27u L=0.06u
MPA3 Y C VDD VNW PCH W=0.27u L=0.06u
.ENDS	NAND3X0P5AA10TR

****
.SUBCKT NAND3X0P5MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=0.29u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.29u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.29u L=0.06u
MPA1 Y A VDD VNW PCH W=0.18u L=0.06u
MPA2 Y B VDD VNW PCH W=0.18u L=0.06u
MPA3 Y C VDD VNW PCH W=0.18u L=0.06u
.ENDS	NAND3X0P5MA10TR

****
.SUBCKT NAND3X0P7AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=0.41u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.41u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.38u L=0.06u
MPA2 Y B VDD VNW PCH W=0.38u L=0.06u
MPA3 Y C VDD VNW PCH W=0.38u L=0.06u
.ENDS	NAND3X0P7AA10TR

****
.SUBCKT NAND3X0P7MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=0.41u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.41u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.25u L=0.06u
MPA2 Y B VDD VNW PCH W=0.25u L=0.06u
MPA3 Y C VDD VNW PCH W=0.25u L=0.06u
.ENDS	NAND3X0P7MA10TR

****
.SUBCKT NAND3X1AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=0.58u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.58u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.54u L=0.06u
MPA2 Y B VDD VNW PCH W=0.54u L=0.06u
MPA3 Y C VDD VNW PCH W=0.54u L=0.06u
.ENDS	NAND3X1AA10TR

****
.SUBCKT NAND3X1MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=0.58u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.58u L=0.06u
MNA3 N1 C VSS VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.36u L=0.06u
MPA2 Y B VDD VNW PCH W=0.36u L=0.06u
MPA3 Y C VDD VNW PCH W=0.36u L=0.06u
.ENDS	NAND3X1MA10TR

****

****

****

****

****
.SUBCKT NAND3X3AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=1.74u L=0.06u
MNA2 N2 B N1 VPW NCH W=1.74u L=0.06u
MNA3 N1 C VSS VPW NCH W=1.74u L=0.06u
MPA1 Y A VDD VNW PCH W=1.62u L=0.06u
MPA2 Y B VDD VNW PCH W=1.62u L=0.06u
MPA3 Y C VDD VNW PCH W=1.62u L=0.06u
.ENDS	NAND3X3AA10TR

****

****
.SUBCKT NAND3X4AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=2.32u L=0.06u
MNA2 N2 B N1 VPW NCH W=2.32u L=0.06u
MNA3 N1 C VSS VPW NCH W=2.32u L=0.06u
MPA1 Y A VDD VNW PCH W=2.16u L=0.06u
MPA2 Y B VDD VNW PCH W=2.16u L=0.06u
MPA3 Y C VDD VNW PCH W=2.16u L=0.06u
.ENDS	NAND3X4AA10TR

****
.SUBCKT NAND3X4MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=2.32u L=0.06u
MNA2 N2 B N1 VPW NCH W=2.32u L=0.06u
MNA3 N1 C VSS VPW NCH W=2.32u L=0.06u
MPA1 Y A VDD VNW PCH W=1.44u L=0.06u
MPA2 Y B VDD VNW PCH W=1.44u L=0.06u
MPA3 Y C VDD VNW PCH W=1.44u L=0.06u
.ENDS	NAND3X4MA10TR

****
.SUBCKT NAND3X6AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=3.48u L=0.06u
MNA2 N2 B N1 VPW NCH W=3.48u L=0.06u
MNA3 N1 C VSS VPW NCH W=3.48u L=0.06u
MPA1 Y A VDD VNW PCH W=3.24u L=0.06u
MPA2 Y B VDD VNW PCH W=3.24u L=0.06u
MPA3 Y C VDD VNW PCH W=3.24u L=0.06u
.ENDS	NAND3X6AA10TR

****
.SUBCKT NAND3X6MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A N2 VPW NCH W=3.48u L=0.06u
MNA2 N2 B N1 VPW NCH W=3.48u L=0.06u
MNA3 N1 C VSS VPW NCH W=3.48u L=0.06u
MPA1 Y A VDD VNW PCH W=2.16u L=0.06u
MPA2 Y B VDD VNW PCH W=2.16u L=0.06u
MPA3 Y C VDD VNW PCH W=2.16u L=0.06u
.ENDS	NAND3X6MA10TR

****
.SUBCKT NAND3XXBX0P5MA10TR  VDD VSS VPW VNW Y   A B CN
MNA1 NET14 CN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y A N2 VPW NCH W=0.29u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.29u L=0.06u
MNA3 N1 NET14 VSS VPW NCH W=0.29u L=0.06u
MPA1 NET14 CN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y A VDD VNW PCH W=0.18u L=0.06u
MPA2 Y B VDD VNW PCH W=0.18u L=0.06u
MPA3 Y NET14 VDD VNW PCH W=0.18u L=0.06u
.ENDS	NAND3XXBX0P5MA10TR

****
.SUBCKT NAND3XXBX0P7MA10TR  VDD VSS VPW VNW Y   A B CN
MNA1 NET14 CN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y A N2 VPW NCH W=0.41u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.41u L=0.06u
MNA3 N1 NET14 VSS VPW NCH W=0.41u L=0.06u
MPA1 NET14 CN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y A VDD VNW PCH W=0.25u L=0.06u
MPA2 Y B VDD VNW PCH W=0.25u L=0.06u
MPA3 Y NET14 VDD VNW PCH W=0.25u L=0.06u
.ENDS	NAND3XXBX0P7MA10TR

****
.SUBCKT NAND3XXBX1MA10TR  VDD VSS VPW VNW Y   A B CN
MNA1 NET14 CN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y A N2 VPW NCH W=0.58u L=0.06u
MNA2 N2 B N1 VPW NCH W=0.58u L=0.06u
MNA3 N1 NET14 VSS VPW NCH W=0.58u L=0.06u
MPA1 NET14 CN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y A VDD VNW PCH W=0.36u L=0.06u
MPA2 Y B VDD VNW PCH W=0.36u L=0.06u
MPA3 Y NET14 VDD VNW PCH W=0.36u L=0.06u
.ENDS	NAND3XXBX1MA10TR

****

****

****
.SUBCKT NAND3XXBX3MA10TR  VDD VSS VPW VNW Y   A B CN
MNA1 NET14 CN VSS VPW NCH W=0.385u L=0.06u
MNA102 Y A N2 VPW NCH W=1.74u L=0.06u
MNA2 N2 B N1 VPW NCH W=1.74u L=0.06u
MNA3 N1 NET14 VSS VPW NCH W=1.74u L=0.06u
MPA1 NET14 CN VDD VNW PCH W=0.51u L=0.06u
MPA105 Y A VDD VNW PCH W=1.08u L=0.06u
MPA2 Y B VDD VNW PCH W=1.08u L=0.06u
MPA3 Y NET14 VDD VNW PCH W=1.08u L=0.06u
.ENDS	NAND3XXBX3MA10TR

****
.SUBCKT NAND3XXBX4MA10TR  VDD VSS VPW VNW Y   A B CN
MNA1 NET14 CN VSS VPW NCH W=0.5u L=0.06u
MNA102 Y A N2 VPW NCH W=2.32u L=0.06u
MNA2 N2 B N1 VPW NCH W=2.32u L=0.06u
MNA3 N1 NET14 VSS VPW NCH W=2.32u L=0.06u
MPA1 NET14 CN VDD VNW PCH W=0.66u L=0.06u
MPA105 Y A VDD VNW PCH W=1.44u L=0.06u
MPA2 Y B VDD VNW PCH W=1.44u L=0.06u
MPA3 Y NET14 VDD VNW PCH W=1.44u L=0.06u
.ENDS	NAND3XXBX4MA10TR

****
.SUBCKT NAND3XXBX6MA10TR  VDD VSS VPW VNW Y   A B CN
MNA1 NET14 CN VSS VPW NCH W=0.75u L=0.06u
MNA102 Y A N2 VPW NCH W=3.48u L=0.06u
MNA2 N2 B N1 VPW NCH W=3.48u L=0.06u
MNA3 N1 NET14 VSS VPW NCH W=3.48u L=0.06u
MPA1 NET14 CN VDD VNW PCH W=0.99u L=0.06u
MPA105 Y A VDD VNW PCH W=2.16u L=0.06u
MPA2 Y B VDD VNW PCH W=2.16u L=0.06u
MPA3 Y NET14 VDD VNW PCH W=2.16u L=0.06u
.ENDS	NAND3XXBX6MA10TR

****
.SUBCKT NAND4BX0P5MA10TR  VDD VSS VPW VNW Y   AN B C D
MNA1 NET32 AN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET32 N3 VPW NCH W=0.31u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.31u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.31u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.31u L=0.06u
MPA1 NET32 AN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y NET32 VDD VNW PCH W=0.15u L=0.06u
MPA2 Y B VDD VNW PCH W=0.15u L=0.06u
MPA3 Y C VDD VNW PCH W=0.15u L=0.06u
MPA4 Y D VDD VNW PCH W=0.15u L=0.06u
.ENDS	NAND4BX0P5MA10TR

****
.SUBCKT NAND4BX0P7MA10TR  VDD VSS VPW VNW Y   AN B C D
MNA1 NET32 AN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET32 N3 VPW NCH W=0.41u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.41u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.41u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.41u L=0.06u
MPA1 NET32 AN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y NET32 VDD VNW PCH W=0.2u L=0.06u
MPA2 Y B VDD VNW PCH W=0.2u L=0.06u
MPA3 Y C VDD VNW PCH W=0.2u L=0.06u
MPA4 Y D VDD VNW PCH W=0.2u L=0.06u
.ENDS	NAND4BX0P7MA10TR

****
.SUBCKT NAND4BX1MA10TR  VDD VSS VPW VNW Y   AN B C D
MNA1 NET32 AN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y NET32 N3 VPW NCH W=0.58u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.58u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.58u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.58u L=0.06u
MPA1 NET32 AN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y NET32 VDD VNW PCH W=0.285u L=0.06u
MPA2 Y B VDD VNW PCH W=0.285u L=0.06u
MPA3 Y C VDD VNW PCH W=0.285u L=0.06u
MPA4 Y D VDD VNW PCH W=0.285u L=0.06u
.ENDS	NAND4BX1MA10TR

****

****

****
.SUBCKT NAND4BX3MA10TR  VDD VSS VPW VNW Y   AN B C D
MNA1 NET32 AN VSS VPW NCH W=0.395u L=0.06u
MNA102 Y NET32 N3 VPW NCH W=1.74u L=0.06u
MNA2 N3 B N2 VPW NCH W=1.74u L=0.06u
MNA3 N2 C N1 VPW NCH W=1.74u L=0.06u
MNA4 N1 D VSS VPW NCH W=1.74u L=0.06u
MPA1 NET32 AN VDD VNW PCH W=0.52u L=0.06u
MPA105 Y NET32 VDD VNW PCH W=0.855u L=0.06u
MPA2 Y B VDD VNW PCH W=0.855u L=0.06u
MPA3 Y C VDD VNW PCH W=0.855u L=0.06u
MPA4 Y D VDD VNW PCH W=0.855u L=0.06u
.ENDS	NAND4BX3MA10TR

****
.SUBCKT NAND4BX4MA10TR  VDD VSS VPW VNW Y   AN B C D
MNA1 NET32 AN VSS VPW NCH W=0.515u L=0.06u
MNA102 Y NET32 N3 VPW NCH W=2.32u L=0.06u
MNA2 N3 B N2 VPW NCH W=2.32u L=0.06u
MNA3 N2 C N1 VPW NCH W=2.32u L=0.06u
MNA4 N1 D VSS VPW NCH W=2.32u L=0.06u
MPA1 NET32 AN VDD VNW PCH W=0.68u L=0.06u
MPA105 Y NET32 VDD VNW PCH W=1.14u L=0.06u
MPA2 Y B VDD VNW PCH W=1.14u L=0.06u
MPA3 Y C VDD VNW PCH W=1.14u L=0.06u
MPA4 Y D VDD VNW PCH W=1.14u L=0.06u
.ENDS	NAND4BX4MA10TR

****
.SUBCKT NAND4X0P5AA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=0.29u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.29u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.29u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.29u L=0.06u
MPA1 Y A VDD VNW PCH W=0.24u L=0.06u
MPA2 Y B VDD VNW PCH W=0.24u L=0.06u
MPA3 Y C VDD VNW PCH W=0.24u L=0.06u
MPA4 Y D VDD VNW PCH W=0.24u L=0.06u
.ENDS	NAND4X0P5AA10TR

****
.SUBCKT NAND4X0P5MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=0.31u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.31u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.31u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.31u L=0.06u
MPA1 Y A VDD VNW PCH W=0.15u L=0.06u
MPA2 Y B VDD VNW PCH W=0.15u L=0.06u
MPA3 Y C VDD VNW PCH W=0.15u L=0.06u
MPA4 Y D VDD VNW PCH W=0.15u L=0.06u
.ENDS	NAND4X0P5MA10TR

****
.SUBCKT NAND4X0P7AA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=0.41u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.41u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.41u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.34u L=0.06u
MPA2 Y B VDD VNW PCH W=0.34u L=0.06u
MPA3 Y C VDD VNW PCH W=0.34u L=0.06u
MPA4 Y D VDD VNW PCH W=0.34u L=0.06u
.ENDS	NAND4X0P7AA10TR

****
.SUBCKT NAND4X0P7MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=0.41u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.41u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.41u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.2u L=0.06u
MPA2 Y B VDD VNW PCH W=0.2u L=0.06u
MPA3 Y C VDD VNW PCH W=0.2u L=0.06u
MPA4 Y D VDD VNW PCH W=0.2u L=0.06u
.ENDS	NAND4X0P7MA10TR

****
.SUBCKT NAND4X1AA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=0.58u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.58u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.58u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
MPA3 Y C VDD VNW PCH W=0.48u L=0.06u
MPA4 Y D VDD VNW PCH W=0.48u L=0.06u
.ENDS	NAND4X1AA10TR

****
.SUBCKT NAND4X1MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=0.58u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.58u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.58u L=0.06u
MNA4 N1 D VSS VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.285u L=0.06u
MPA2 Y B VDD VNW PCH W=0.285u L=0.06u
MPA3 Y C VDD VNW PCH W=0.285u L=0.06u
MPA4 Y D VDD VNW PCH W=0.285u L=0.06u
.ENDS	NAND4X1MA10TR

****

****

****

****

****
.SUBCKT NAND4X3AA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=1.74u L=0.06u
MNA2 N3 B N2 VPW NCH W=1.74u L=0.06u
MNA3 N2 C N1 VPW NCH W=1.74u L=0.06u
MNA4 N1 D VSS VPW NCH W=1.74u L=0.06u
MPA1 Y A VDD VNW PCH W=1.44u L=0.06u
MPA2 Y B VDD VNW PCH W=1.44u L=0.06u
MPA3 Y C VDD VNW PCH W=1.44u L=0.06u
MPA4 Y D VDD VNW PCH W=1.44u L=0.06u
.ENDS	NAND4X3AA10TR

****
.SUBCKT NAND4X3MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=1.74u L=0.06u
MNA2 N3 B N2 VPW NCH W=1.74u L=0.06u
MNA3 N2 C N1 VPW NCH W=1.74u L=0.06u
MNA4 N1 D VSS VPW NCH W=1.74u L=0.06u
MPA1 Y A VDD VNW PCH W=0.855u L=0.06u
MPA2 Y B VDD VNW PCH W=0.855u L=0.06u
MPA3 Y C VDD VNW PCH W=0.855u L=0.06u
MPA4 Y D VDD VNW PCH W=0.855u L=0.06u
.ENDS	NAND4X3MA10TR

****
.SUBCKT NAND4X4AA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=2.32u L=0.06u
MNA2 N3 B N2 VPW NCH W=2.32u L=0.06u
MNA3 N2 C N1 VPW NCH W=2.32u L=0.06u
MNA4 N1 D VSS VPW NCH W=2.32u L=0.06u
MPA1 Y A VDD VNW PCH W=1.92u L=0.06u
MPA2 Y B VDD VNW PCH W=1.92u L=0.06u
MPA3 Y C VDD VNW PCH W=1.92u L=0.06u
MPA4 Y D VDD VNW PCH W=1.92u L=0.06u
.ENDS	NAND4X4AA10TR

****
.SUBCKT NAND4X4MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 Y A N3 VPW NCH W=2.32u L=0.06u
MNA2 N3 B N2 VPW NCH W=2.32u L=0.06u
MNA3 N2 C N1 VPW NCH W=2.32u L=0.06u
MNA4 N1 D VSS VPW NCH W=2.32u L=0.06u
MPA1 Y A VDD VNW PCH W=1.14u L=0.06u
MPA2 Y B VDD VNW PCH W=1.14u L=0.06u
MPA3 Y C VDD VNW PCH W=1.14u L=0.06u
MPA4 Y D VDD VNW PCH W=1.14u L=0.06u
.ENDS	NAND4X4MA10TR

****
.SUBCKT NAND4XXXBX0P5MA10TR  VDD VSS VPW VNW Y   A B C DN
MNA1 NET32 DN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y A N3 VPW NCH W=0.31u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.31u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.31u L=0.06u
MNA4 N1 NET32 VSS VPW NCH W=0.31u L=0.06u
MPA1 NET32 DN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y A VDD VNW PCH W=0.15u L=0.06u
MPA2 Y B VDD VNW PCH W=0.15u L=0.06u
MPA3 Y C VDD VNW PCH W=0.15u L=0.06u
MPA4 Y NET32 VDD VNW PCH W=0.15u L=0.06u
.ENDS	NAND4XXXBX0P5MA10TR

****
.SUBCKT NAND4XXXBX0P7MA10TR  VDD VSS VPW VNW Y   A B C DN
MNA1 NET32 DN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y A N3 VPW NCH W=0.41u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.41u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.41u L=0.06u
MNA4 N1 NET32 VSS VPW NCH W=0.41u L=0.06u
MPA1 NET32 DN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y A VDD VNW PCH W=0.2u L=0.06u
MPA2 Y B VDD VNW PCH W=0.2u L=0.06u
MPA3 Y C VDD VNW PCH W=0.2u L=0.06u
MPA4 Y NET32 VDD VNW PCH W=0.2u L=0.06u
.ENDS	NAND4XXXBX0P7MA10TR

****
.SUBCKT NAND4XXXBX1MA10TR  VDD VSS VPW VNW Y   A B C DN
MNA1 NET32 DN VSS VPW NCH W=0.15u L=0.06u
MNA102 Y A N3 VPW NCH W=0.58u L=0.06u
MNA2 N3 B N2 VPW NCH W=0.58u L=0.06u
MNA3 N2 C N1 VPW NCH W=0.58u L=0.06u
MNA4 N1 NET32 VSS VPW NCH W=0.58u L=0.06u
MPA1 NET32 DN VDD VNW PCH W=0.2u L=0.06u
MPA105 Y A VDD VNW PCH W=0.28u L=0.06u
MPA2 Y B VDD VNW PCH W=0.28u L=0.06u
MPA3 Y C VDD VNW PCH W=0.28u L=0.06u
MPA4 Y NET32 VDD VNW PCH W=0.28u L=0.06u
.ENDS	NAND4XXXBX1MA10TR

****

****

****
.SUBCKT NAND4XXXBX3MA10TR  VDD VSS VPW VNW Y   A B C DN
MNA1 NET32 DN VSS VPW NCH W=0.395u L=0.06u
MNA102 Y A N3 VPW NCH W=1.74u L=0.06u
MNA2 N3 B N2 VPW NCH W=1.74u L=0.06u
MNA3 N2 C N1 VPW NCH W=1.74u L=0.06u
MNA4 N1 NET32 VSS VPW NCH W=1.74u L=0.06u
MPA1 NET32 DN VDD VNW PCH W=0.52u L=0.06u
MPA105 Y A VDD VNW PCH W=0.855u L=0.06u
MPA2 Y B VDD VNW PCH W=0.855u L=0.06u
MPA3 Y C VDD VNW PCH W=0.855u L=0.06u
MPA4 Y NET32 VDD VNW PCH W=0.855u L=0.06u
.ENDS	NAND4XXXBX3MA10TR

****
.SUBCKT NAND4XXXBX4MA10TR  VDD VSS VPW VNW Y   A B C DN
MNA1 NET32 DN VSS VPW NCH W=0.515u L=0.06u
MNA102 Y A N3 VPW NCH W=2.32u L=0.06u
MNA2 N3 B N2 VPW NCH W=2.32u L=0.06u
MNA3 N2 C N1 VPW NCH W=2.32u L=0.06u
MNA4 N1 NET32 VSS VPW NCH W=2.32u L=0.06u
MPA1 NET32 DN VDD VNW PCH W=0.68u L=0.06u
MPA105 Y A VDD VNW PCH W=1.14u L=0.06u
MPA2 Y B VDD VNW PCH W=1.14u L=0.06u
MPA3 Y C VDD VNW PCH W=1.14u L=0.06u
MPA4 Y NET32 VDD VNW PCH W=1.14u L=0.06u
.ENDS	NAND4XXXBX4MA10TR

****
.SUBCKT NOR2BX0P5MA10TR  VDD VSS VPW VNW Y   AN B
MNA1 Y NET24 VSS VPW NCH W=0.15u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.15u L=0.06u
MNA2 Y B VSS VPW NCH W=0.15u L=0.06u
MPA1 Y NET24 P1 VNW PCH W=0.37u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.2u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.37u L=0.06u
.ENDS	NOR2BX0P5MA10TR

****
.SUBCKT NOR2BX0P7MA10TR  VDD VSS VPW VNW Y   AN B
MNA1 Y NET24 VSS VPW NCH W=0.2u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.15u L=0.06u
MNA2 Y B VSS VPW NCH W=0.2u L=0.06u
MPA1 Y NET24 P1 VNW PCH W=0.49u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.2u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.49u L=0.06u
.ENDS	NOR2BX0P7MA10TR

****
.SUBCKT NOR2BX1MA10TR  VDD VSS VPW VNW Y   AN B
MNA1 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.15u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1 Y NET24 P1 VNW PCH W=0.7u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.2u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.7u L=0.06u
.ENDS	NOR2BX1MA10TR

****

****

****

****

****

****

****
.SUBCKT NOR2X0P5AA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A VSS VPW NCH W=0.245u L=0.06u
MNA2 Y B VSS VPW NCH W=0.245u L=0.06u
MPA1 Y A P1 VNW PCH W=0.37u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.37u L=0.06u
.ENDS	NOR2X0P5AA10TR

****
.SUBCKT NOR2X0P5MA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A VSS VPW NCH W=0.15u L=0.06u
MNA2 Y B VSS VPW NCH W=0.15u L=0.06u
MPA1 Y A P1 VNW PCH W=0.37u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.37u L=0.06u
.ENDS	NOR2X0P5MA10TR

****
.SUBCKT NOR2X0P7AA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A VSS VPW NCH W=0.345u L=0.06u
MNA2 Y B VSS VPW NCH W=0.345u L=0.06u
MPA1 Y A P1 VNW PCH W=0.49u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.49u L=0.06u
.ENDS	NOR2X0P7AA10TR

****
.SUBCKT NOR2X0P7MA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A VSS VPW NCH W=0.2u L=0.06u
MNA2 Y B VSS VPW NCH W=0.2u L=0.06u
MPA1 Y A P1 VNW PCH W=0.49u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.49u L=0.06u
.ENDS	NOR2X0P7MA10TR

****
.SUBCKT NOR2X1AA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A VSS VPW NCH W=0.49u L=0.06u
MNA2 Y B VSS VPW NCH W=0.49u L=0.06u
MPA1 Y A P1 VNW PCH W=0.7u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.7u L=0.06u
.ENDS	NOR2X1AA10TR

****
.SUBCKT NOR2X1MA10TR  VDD VSS VPW VNW Y   A B
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A P1 VNW PCH W=0.7u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.7u L=0.06u
.ENDS	NOR2X1MA10TR

****

****

****

****

****

****

****

****

****

****

****

****

****
.SUBCKT NOR2XBX0P5MA10TR  VDD VSS VPW VNW Y   A BN
MNA1 Y A VSS VPW NCH W=0.15u L=0.06u
MNA104 NET014 BN VSS VPW NCH W=0.15u L=0.06u
MNA2 Y NET014 VSS VPW NCH W=0.15u L=0.06u
MPA1 Y A P1 VNW PCH W=0.37u L=0.06u
MPA106 NET014 BN VDD VNW PCH W=0.2u L=0.06u
MPA2 P1 NET014 VDD VNW PCH W=0.37u L=0.06u
.ENDS	NOR2XBX0P5MA10TR

****
.SUBCKT NOR2XBX0P7MA10TR  VDD VSS VPW VNW Y   A BN
MNA1 Y A VSS VPW NCH W=0.2u L=0.06u
MNA104 NET014 BN VSS VPW NCH W=0.15u L=0.06u
MNA2 Y NET014 VSS VPW NCH W=0.2u L=0.06u
MPA1 Y A P1 VNW PCH W=0.49u L=0.06u
MPA106 NET014 BN VDD VNW PCH W=0.2u L=0.06u
MPA2 P1 NET014 VDD VNW PCH W=0.49u L=0.06u
.ENDS	NOR2XBX0P7MA10TR

****
.SUBCKT NOR2XBX1MA10TR  VDD VSS VPW VNW Y   A BN
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MNA104 NET014 BN VSS VPW NCH W=0.15u L=0.06u
MNA2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A P1 VNW PCH W=0.7u L=0.06u
MPA106 NET014 BN VDD VNW PCH W=0.2u L=0.06u
MPA2 P1 NET014 VDD VNW PCH W=0.7u L=0.06u
.ENDS	NOR2XBX1MA10TR

****

****

****

****

****

****

****
.SUBCKT NOR3X0P5AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A VSS VPW NCH W=0.19u L=0.06u
MNA2 Y B VSS VPW NCH W=0.19u L=0.06u
MNA3 Y C VSS VPW NCH W=0.19u L=0.06u
MPA1 Y A P2 VNW PCH W=0.35u L=0.06u
MPA2 P2 B P1 VNW PCH W=0.35u L=0.06u
MPA3 P1 C VDD VNW PCH W=0.35u L=0.06u
.ENDS	NOR3X0P5AA10TR

****
.SUBCKT NOR3X0P5MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A VSS VPW NCH W=0.15u L=0.06u
MNA2 Y B VSS VPW NCH W=0.15u L=0.06u
MNA3 Y C VSS VPW NCH W=0.15u L=0.06u
MPA1 Y A P2 VNW PCH W=0.35u L=0.06u
MPA2 P2 B P1 VNW PCH W=0.35u L=0.06u
MPA3 P1 C VDD VNW PCH W=0.35u L=0.06u
.ENDS	NOR3X0P5MA10TR

****
.SUBCKT NOR3X0P7AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A VSS VPW NCH W=0.27u L=0.06u
MNA2 Y B VSS VPW NCH W=0.27u L=0.06u
MNA3 Y C VSS VPW NCH W=0.27u L=0.06u
MPA1 Y A P2 VNW PCH W=0.49u L=0.06u
MPA2 P2 B P1 VNW PCH W=0.49u L=0.06u
MPA3 P1 C VDD VNW PCH W=0.49u L=0.06u
.ENDS	NOR3X0P7AA10TR

****

****
.SUBCKT NOR3X1AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A VSS VPW NCH W=0.38u L=0.06u
MNA2 Y B VSS VPW NCH W=0.38u L=0.06u
MNA3 Y C VSS VPW NCH W=0.38u L=0.06u
MPA1 Y A P2 VNW PCH W=0.7u L=0.06u
MPA2 P2 B P1 VNW PCH W=0.7u L=0.06u
MPA3 P1 C VDD VNW PCH W=0.7u L=0.06u
.ENDS	NOR3X1AA10TR

****

****

****

****

****

****
.SUBCKT NOR3X3AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A VSS VPW NCH W=1.14u L=0.06u
MNA2 Y B VSS VPW NCH W=1.14u L=0.06u
MNA3 Y C VSS VPW NCH W=1.14u L=0.06u
MPA1 Y A P2 VNW PCH W=2.1u L=0.06u
MPA2 P2 B P1 VNW PCH W=2.1u L=0.06u
MPA3 P1 C VDD VNW PCH W=2.1u L=0.06u
.ENDS	NOR3X3AA10TR

****
.SUBCKT NOR3X3MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A VSS VPW NCH W=0.615u L=0.06u
MNA2 Y B VSS VPW NCH W=0.615u L=0.06u
MNA3 Y C VSS VPW NCH W=0.615u L=0.06u
MPA1 Y A P2 VNW PCH W=2.1u L=0.06u
MPA2 P2 B P1 VNW PCH W=2.1u L=0.06u
MPA3 P1 C VDD VNW PCH W=2.1u L=0.06u
.ENDS	NOR3X3MA10TR

****
.SUBCKT NOR3X4AA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A VSS VPW NCH W=1.52u L=0.06u
MNA2 Y B VSS VPW NCH W=1.52u L=0.06u
MNA3 Y C VSS VPW NCH W=1.52u L=0.06u
MPA1 Y A P2 VNW PCH W=2.8u L=0.06u
MPA2 P2 B P1 VNW PCH W=2.8u L=0.06u
MPA3 P1 C VDD VNW PCH W=2.8u L=0.06u
.ENDS	NOR3X4AA10TR

****
.SUBCKT NOR3X4MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y A VSS VPW NCH W=0.82u L=0.06u
MNA2 Y B VSS VPW NCH W=0.82u L=0.06u
MNA3 Y C VSS VPW NCH W=0.82u L=0.06u
MPA1 Y A P2 VNW PCH W=2.8u L=0.06u
MPA2 P2 B P1 VNW PCH W=2.8u L=0.06u
MPA3 P1 C VDD VNW PCH W=2.8u L=0.06u
.ENDS	NOR3X4MA10TR

****
.SUBCKT OA211X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 C0
MNA1 INT C0 N2 VPW NCH W=0.42u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.265u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.42u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.42u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.42u L=0.06u
MPA1 INT C0 VDD VNW PCH W=0.255u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.35u L=0.06u
MPB1 INT B0 VDD VNW PCH W=0.255u L=0.06u
MPC1 INT A0 P1 VNW PCH W=0.54u L=0.06u
MPC2 P1 A1 VDD VNW PCH W=0.54u L=0.06u
.ENDS	OA211X0P5MA10TR

****
.SUBCKT OA211X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 C0
MNA1 INT C0 N2 VPW NCH W=0.5u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.37u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.5u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.5u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.5u L=0.06u
MPA1 INT C0 VDD VNW PCH W=0.305u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.49u L=0.06u
MPB1 INT B0 VDD VNW PCH W=0.305u L=0.06u
MPC1 INT A0 P1 VNW PCH W=0.65u L=0.06u
MPC2 P1 A1 VDD VNW PCH W=0.65u L=0.06u
.ENDS	OA211X0P7MA10TR

****

****

****

****

****

****

****
.SUBCKT OA21X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA106 INT B0 N1 VPW NCH W=0.22u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.22u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.22u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA108 INT B0 VDD VNW PCH W=0.18u L=0.06u
MPB1 INT A0 P1 VNW PCH W=0.36u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.36u L=0.06u
.ENDS	OA21X0P5MA10TR

****
.SUBCKT OA21X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MNA106 INT B0 N1 VPW NCH W=0.27u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.27u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.27u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA108 INT B0 VDD VNW PCH W=0.225u L=0.06u
MPB1 INT A0 P1 VNW PCH W=0.45u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.45u L=0.06u
.ENDS	OA21X0P7MA10TR

****
.SUBCKT OA21X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MNA106 INT B0 N1 VPW NCH W=0.355u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.355u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.355u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA108 INT B0 VDD VNW PCH W=0.29u L=0.06u
MPB1 INT A0 P1 VNW PCH W=0.585u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.585u L=0.06u
.ENDS	OA21X1MA10TR

****

****

****

****

****
.SUBCKT OA21X6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=3.18u L=0.06u
MNA106 INT B0 N1 VPW NCH W=1.92u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=1.92u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.92u L=0.06u
MPA1 Y INT VDD VNW PCH W=4.2u L=0.06u
MPA108 INT B0 VDD VNW PCH W=1.575u L=0.06u
MPB1 INT A0 P1 VNW PCH W=3.175u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=3.175u L=0.06u
.ENDS	OA21X6MA10TR

****
.SUBCKT OA21X8MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y INT VSS VPW NCH W=4.24u L=0.06u
MNA106 INT B0 N1 VPW NCH W=2.55u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=2.55u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=2.55u L=0.06u
MPA1 Y INT VDD VNW PCH W=5.6u L=0.06u
MPA108 INT B0 VDD VNW PCH W=2.1u L=0.06u
MPB1 INT A0 P1 VNW PCH W=4.2u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=4.2u L=0.06u
.ENDS	OA21X8MA10TR

****
.SUBCKT OA22X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 INT B0 N1 VPW NCH W=0.245u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA2 INT B1 N1 VPW NCH W=0.245u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.245u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.245u L=0.06u
MPA1 INT B0 P1A VNW PCH W=0.365u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=0.365u L=0.06u
MPB1 INT A0 P1B VNW PCH W=0.365u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=0.365u L=0.06u
.ENDS	OA22X0P5MA10TR

****
.SUBCKT OA22X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 INT B0 N1 VPW NCH W=0.3u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.37u L=0.06u
MNA2 INT B1 N1 VPW NCH W=0.3u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.3u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.3u L=0.06u
MPA1 INT B0 P1A VNW PCH W=0.45u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=0.45u L=0.06u
MPB1 INT A0 P1B VNW PCH W=0.45u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=0.45u L=0.06u
.ENDS	OA22X0P7MA10TR

****
.SUBCKT OA22X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 INT B0 N1 VPW NCH W=0.39u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.53u L=0.06u
MNA2 INT B1 N1 VPW NCH W=0.39u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.39u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.39u L=0.06u
MPA1 INT B0 P1A VNW PCH W=0.58u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=0.58u L=0.06u
MPB1 INT A0 P1B VNW PCH W=0.58u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=0.58u L=0.06u
.ENDS	OA22X1MA10TR

****

****

****
.SUBCKT OA22X3MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 INT B0 N1 VPW NCH W=1.065u L=0.06u
MNA108 Y INT VSS VPW NCH W=1.59u L=0.06u
MNA2 INT B1 N1 VPW NCH W=1.065u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=1.065u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.065u L=0.06u
MPA1 INT B0 P1A VNW PCH W=1.59u L=0.06u
MPA1010 Y INT VDD VNW PCH W=2.1u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=1.59u L=0.06u
MPB1 INT A0 P1B VNW PCH W=1.59u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=1.59u L=0.06u
.ENDS	OA22X3MA10TR

****
.SUBCKT OA22X4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 INT B0 N1 VPW NCH W=1.41u L=0.06u
MNA108 Y INT VSS VPW NCH W=2.12u L=0.06u
MNA2 INT B1 N1 VPW NCH W=1.41u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=1.41u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.41u L=0.06u
MPA1 INT B0 P1A VNW PCH W=2.1u L=0.06u
MPA1010 Y INT VDD VNW PCH W=2.8u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=2.1u L=0.06u
MPB1 INT A0 P1B VNW PCH W=2.1u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=2.1u L=0.06u
.ENDS	OA22X4MA10TR

****
.SUBCKT OA22X6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 INT B0 N1 VPW NCH W=2.1u L=0.06u
MNA108 Y INT VSS VPW NCH W=3.18u L=0.06u
MNA2 INT B1 N1 VPW NCH W=2.1u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=2.1u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=2.1u L=0.06u
MPA1 INT B0 P1A VNW PCH W=3.125u L=0.06u
MPA1010 Y INT VDD VNW PCH W=4.2u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=3.125u L=0.06u
MPB1 INT A0 P1B VNW PCH W=3.125u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=3.125u L=0.06u
.ENDS	OA22X6MA10TR

****
.SUBCKT OA22X8MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 INT B0 N1 VPW NCH W=2.82u L=0.06u
MNA108 Y INT VSS VPW NCH W=4.24u L=0.06u
MNA2 INT B1 N1 VPW NCH W=2.82u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=2.82u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=2.82u L=0.06u
MPA1 INT B0 P1A VNW PCH W=4.2u L=0.06u
MPA1010 Y INT VDD VNW PCH W=5.6u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=4.2u L=0.06u
MPB1 INT A0 P1B VNW PCH W=4.2u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=4.2u L=0.06u
.ENDS	OA22X8MA10TR

****
.SUBCKT OAI211X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 C0
MNA1 Y C0 N2 VPW NCH W=0.29u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.29u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.29u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.29u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.18u L=0.06u
MPB1 Y B0 VDD VNW PCH W=0.18u L=0.06u
MPC1 Y A0 P1 VNW PCH W=0.335u L=0.06u
MPC2 P1 A1 VDD VNW PCH W=0.335u L=0.06u
.ENDS	OAI211X0P5MA10TR

****
.SUBCKT OAI211X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 C0
MNA1 Y C0 N2 VPW NCH W=0.41u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.41u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.41u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.41u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.25u L=0.06u
MPB1 Y B0 VDD VNW PCH W=0.25u L=0.06u
MPC1 Y A0 P1 VNW PCH W=0.47u L=0.06u
MPC2 P1 A1 VDD VNW PCH W=0.47u L=0.06u
.ENDS	OAI211X0P7MA10TR

****
.SUBCKT OAI211X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 C0
MNA1 Y C0 N2 VPW NCH W=0.58u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.36u L=0.06u
MPB1 Y B0 VDD VNW PCH W=0.36u L=0.06u
MPC1 Y A0 P1 VNW PCH W=0.665u L=0.06u
MPC2 P1 A1 VDD VNW PCH W=0.665u L=0.06u
.ENDS	OAI211X1MA10TR

****

****

****

****

****
.SUBCKT OAI21BX0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.15u L=0.06u
MNA106 Y NET28 N1 VPW NCH W=0.23u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.23u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.23u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.2u L=0.06u
MPA108 Y NET28 VDD VNW PCH W=0.19u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.35u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.35u L=0.06u
.ENDS	OAI21BX0P5MA10TR

****
.SUBCKT OAI21BX0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.15u L=0.06u
MNA106 Y NET28 N1 VPW NCH W=0.32u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.32u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.2u L=0.06u
MPA108 Y NET28 VDD VNW PCH W=0.265u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.49u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
.ENDS	OAI21BX0P7MA10TR

****
.SUBCKT OAI21BX1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.15u L=0.06u
MNA106 Y NET28 N1 VPW NCH W=0.455u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.2u L=0.06u
MPA108 Y NET28 VDD VNW PCH W=0.38u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.7u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
.ENDS	OAI21BX1MA10TR

****
.SUBCKT OAI21BX1P4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.185u L=0.06u
MNA106 Y NET28 N1 VPW NCH W=0.64u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.64u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.64u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.245u L=0.06u
MPA108 Y NET28 VDD VNW PCH W=0.53u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.98u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.98u L=0.06u
.ENDS	OAI21BX1P4MA10TR

****
.SUBCKT OAI21BX2MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.24u L=0.06u
MNA106 Y NET28 N1 VPW NCH W=0.91u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.91u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.91u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.315u L=0.06u
MPA108 Y NET28 VDD VNW PCH W=0.76u L=0.06u
MPB1 Y A0 P1 VNW PCH W=1.4u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=1.4u L=0.06u
.ENDS	OAI21BX2MA10TR

****
.SUBCKT OAI21BX3MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.365u L=0.06u
MNA106 Y NET28 N1 VPW NCH W=1.365u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=1.365u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.365u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.485u L=0.06u
MPA108 Y NET28 VDD VNW PCH W=1.14u L=0.06u
MPB1 Y A0 P1 VNW PCH W=2.1u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.1u L=0.06u
.ENDS	OAI21BX3MA10TR

****
.SUBCKT OAI21BX4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.48u L=0.06u
MNA106 Y NET28 N1 VPW NCH W=1.82u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=1.82u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.82u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.63u L=0.06u
MPA108 Y NET28 VDD VNW PCH W=1.52u L=0.06u
MPB1 Y A0 P1 VNW PCH W=2.8u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.8u L=0.06u
.ENDS	OAI21BX4MA10TR

****
.SUBCKT OAI21BX6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.72u L=0.06u
MNA106 Y NET28 N1 VPW NCH W=2.73u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=2.73u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=2.73u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.95u L=0.06u
MPA108 Y NET28 VDD VNW PCH W=2.28u L=0.06u
MPB1 Y A0 P1 VNW PCH W=4.2u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=4.2u L=0.06u
.ENDS	OAI21BX6MA10TR

****
.SUBCKT OAI21BX8MA10TR  VDD VSS VPW VNW Y   A0 A1 B0N
MNA1 NET28 B0N VSS VPW NCH W=0.96u L=0.06u
MNA106 Y NET28 N1 VPW NCH W=3.64u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=3.64u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=3.64u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=1.26u L=0.06u
MPA108 Y NET28 VDD VNW PCH W=3.04u L=0.06u
MPB1 Y A0 P1 VNW PCH W=5.6u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=5.6u L=0.06u
.ENDS	OAI21BX8MA10TR

****
.SUBCKT OAI21X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 N1 VPW NCH W=0.23u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.23u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.23u L=0.06u
MPA1 Y B0 VDD VNW PCH W=0.19u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.35u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.35u L=0.06u
.ENDS	OAI21X0P5MA10TR

****
.SUBCKT OAI21X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 N1 VPW NCH W=0.32u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.32u L=0.06u
MPA1 Y B0 VDD VNW PCH W=0.265u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.49u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
.ENDS	OAI21X0P7MA10TR

****
.SUBCKT OAI21X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 N1 VPW NCH W=0.455u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPA1 Y B0 VDD VNW PCH W=0.38u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.7u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
.ENDS	OAI21X1MA10TR

****

****

****

****
.SUBCKT OAI21X4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 N1 VPW NCH W=1.82u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=1.82u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.82u L=0.06u
MPA1 Y B0 VDD VNW PCH W=1.52u L=0.06u
MPB1 Y A0 P1 VNW PCH W=2.8u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=2.8u L=0.06u
.ENDS	OAI21X4MA10TR

****
.SUBCKT OAI21X6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 N1 VPW NCH W=2.73u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=2.73u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=2.73u L=0.06u
MPA1 Y B0 VDD VNW PCH W=2.28u L=0.06u
MPB1 Y A0 P1 VNW PCH W=4.2u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=4.2u L=0.06u
.ENDS	OAI21X6MA10TR

****
.SUBCKT OAI21X8MA10TR  VDD VSS VPW VNW Y   A0 A1 B0
MNA1 Y B0 N1 VPW NCH W=3.64u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=3.64u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=3.64u L=0.06u
MPA1 Y B0 VDD VNW PCH W=3.04u L=0.06u
MPB1 Y A0 P1 VNW PCH W=5.6u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=5.6u L=0.06u
.ENDS	OAI21X8MA10TR

****
.SUBCKT OAI221X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0
MNA1 Y C0 N2 VPW NCH W=0.29u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.29u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.29u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.29u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.29u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.18u L=0.06u
MPB1 Y B0 P1B VNW PCH W=0.335u L=0.06u
MPB2 P1B B1 VDD VNW PCH W=0.335u L=0.06u
MPC1 Y A0 P1C VNW PCH W=0.335u L=0.06u
MPC2 P1C A1 VDD VNW PCH W=0.335u L=0.06u
.ENDS	OAI221X0P5MA10TR

****
.SUBCKT OAI221X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0
MNA1 Y C0 N2 VPW NCH W=0.41u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.41u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.41u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.41u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.41u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.25u L=0.06u
MPB1 Y B0 P1B VNW PCH W=0.47u L=0.06u
MPB2 P1B B1 VDD VNW PCH W=0.47u L=0.06u
MPC1 Y A0 P1C VNW PCH W=0.47u L=0.06u
MPC2 P1C A1 VDD VNW PCH W=0.47u L=0.06u
.ENDS	OAI221X0P7MA10TR

****
.SUBCKT OAI221X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0
MNA1 Y C0 N2 VPW NCH W=0.58u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.36u L=0.06u
MPB1 Y B0 P1B VNW PCH W=0.665u L=0.06u
MPB2 P1B B1 VDD VNW PCH W=0.665u L=0.06u
MPC1 Y A0 P1C VNW PCH W=0.665u L=0.06u
MPC2 P1C A1 VDD VNW PCH W=0.665u L=0.06u
.ENDS	OAI221X1MA10TR

****

****

****

****

****
.SUBCKT OAI222X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0 C1
MNA1 Y C0 N2 VPW NCH W=0.29u L=0.06u
MNA2 Y C1 N2 VPW NCH W=0.29u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.29u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.29u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.29u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.29u L=0.06u
MPA1 Y C0 P1A VNW PCH W=0.335u L=0.06u
MPA2 P1A C1 VDD VNW PCH W=0.335u L=0.06u
MPB1 Y B0 P1B VNW PCH W=0.335u L=0.06u
MPB2 P1B B1 VDD VNW PCH W=0.335u L=0.06u
MPC1 Y A0 P1C VNW PCH W=0.335u L=0.06u
MPC2 P1C A1 VDD VNW PCH W=0.335u L=0.06u
.ENDS	OAI222X0P5MA10TR

****
.SUBCKT OAI222X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0 C1
MNA1 Y C0 N2 VPW NCH W=0.41u L=0.06u
MNA2 Y C1 N2 VPW NCH W=0.41u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.41u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.41u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.41u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.41u L=0.06u
MPA1 Y C0 P1A VNW PCH W=0.465u L=0.06u
MPA2 P1A C1 VDD VNW PCH W=0.465u L=0.06u
MPB1 Y B0 P1B VNW PCH W=0.465u L=0.06u
MPB2 P1B B1 VDD VNW PCH W=0.465u L=0.06u
MPC1 Y A0 P1C VNW PCH W=0.465u L=0.06u
MPC2 P1C A1 VDD VNW PCH W=0.465u L=0.06u
.ENDS	OAI222X0P7MA10TR

****
.SUBCKT OAI222X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1 C0 C1
MNA1 Y C0 N2 VPW NCH W=0.58u L=0.06u
MNA2 Y C1 N2 VPW NCH W=0.58u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPA1 Y C0 P1A VNW PCH W=0.665u L=0.06u
MPA2 P1A C1 VDD VNW PCH W=0.665u L=0.06u
MPB1 Y B0 P1B VNW PCH W=0.665u L=0.06u
MPB2 P1B B1 VDD VNW PCH W=0.665u L=0.06u
MPC1 Y A0 P1C VNW PCH W=0.665u L=0.06u
MPC2 P1C A1 VDD VNW PCH W=0.665u L=0.06u
.ENDS	OAI222X1MA10TR

****

****

****

****

****
.SUBCKT OAI22X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1 VPW NCH W=0.23u L=0.06u
MNA2 Y B1 N1 VPW NCH W=0.23u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.23u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.23u L=0.06u
MPA1 Y B0 P1A VNW PCH W=0.35u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=0.35u L=0.06u
MPB1 Y A0 P1B VNW PCH W=0.35u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=0.35u L=0.06u
.ENDS	OAI22X0P5MA10TR

****
.SUBCKT OAI22X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1 VPW NCH W=0.32u L=0.06u
MNA2 Y B1 N1 VPW NCH W=0.32u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.32u L=0.06u
MPA1 Y B0 P1A VNW PCH W=0.49u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=0.49u L=0.06u
MPB1 Y A0 P1B VNW PCH W=0.49u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=0.49u L=0.06u
.ENDS	OAI22X0P7MA10TR

****
.SUBCKT OAI22X1MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1 VPW NCH W=0.455u L=0.06u
MNA2 Y B1 N1 VPW NCH W=0.455u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPA1 Y B0 P1A VNW PCH W=0.7u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=0.7u L=0.06u
MPB1 Y A0 P1B VNW PCH W=0.7u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=0.7u L=0.06u
.ENDS	OAI22X1MA10TR

****

****

****
.SUBCKT OAI22X3MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1 VPW NCH W=1.365u L=0.06u
MNA2 Y B1 N1 VPW NCH W=1.365u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=1.365u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.365u L=0.06u
MPA1 Y B0 P1A VNW PCH W=2.1u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=2.1u L=0.06u
MPB1 Y A0 P1B VNW PCH W=2.1u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=2.1u L=0.06u
.ENDS	OAI22X3MA10TR

****
.SUBCKT OAI22X4MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1 VPW NCH W=1.82u L=0.06u
MNA2 Y B1 N1 VPW NCH W=1.82u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=1.82u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=1.82u L=0.06u
MPA1 Y B0 P1A VNW PCH W=2.8u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=2.8u L=0.06u
MPB1 Y A0 P1B VNW PCH W=2.8u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=2.8u L=0.06u
.ENDS	OAI22X4MA10TR

****
.SUBCKT OAI22X6MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1 VPW NCH W=2.73u L=0.06u
MNA2 Y B1 N1 VPW NCH W=2.73u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=2.73u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=2.73u L=0.06u
MPA1 Y B0 P1A VNW PCH W=4.2u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=4.2u L=0.06u
MPB1 Y A0 P1B VNW PCH W=4.2u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=4.2u L=0.06u
.ENDS	OAI22X6MA10TR

****
.SUBCKT OAI22X8MA10TR  VDD VSS VPW VNW Y   A0 A1 B0 B1
MNA1 Y B0 N1 VPW NCH W=3.64u L=0.06u
MNA2 Y B1 N1 VPW NCH W=3.64u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=3.64u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=3.64u L=0.06u
MPA1 Y B0 P1A VNW PCH W=5.6u L=0.06u
MPA2 P1A B1 VDD VNW PCH W=5.6u L=0.06u
MPB1 Y A0 P1B VNW PCH W=5.6u L=0.06u
MPB2 P1B A1 VDD VNW PCH W=5.6u L=0.06u
.ENDS	OAI22X8MA10TR

****
.SUBCKT OAI2XB1X0P5MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.15u L=0.06u
MNA106 Y B0 N1 VPW NCH W=0.23u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.23u L=0.06u
MNB2 N1 INT VSS VPW NCH W=0.23u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.2u L=0.06u
MPA108 Y B0 VDD VNW PCH W=0.19u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.35u L=0.06u
MPB2 P1 INT VDD VNW PCH W=0.35u L=0.06u
.ENDS	OAI2XB1X0P5MA10TR

****
.SUBCKT OAI2XB1X0P7MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.15u L=0.06u
MNA106 Y B0 N1 VPW NCH W=0.32u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MNB2 N1 INT VSS VPW NCH W=0.32u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.2u L=0.06u
MPA108 Y B0 VDD VNW PCH W=0.265u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.49u L=0.06u
MPB2 P1 INT VDD VNW PCH W=0.49u L=0.06u
.ENDS	OAI2XB1X0P7MA10TR

****
.SUBCKT OAI2XB1X1MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.155u L=0.06u
MNA106 Y B0 N1 VPW NCH W=0.455u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MNB2 N1 INT VSS VPW NCH W=0.455u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.205u L=0.06u
MPA108 Y B0 VDD VNW PCH W=0.38u L=0.06u
MPB1 Y A0 P1 VNW PCH W=0.7u L=0.06u
MPB2 P1 INT VDD VNW PCH W=0.7u L=0.06u
.ENDS	OAI2XB1X1MA10TR

****

****

****

****
.SUBCKT OAI2XB1X4MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.59u L=0.06u
MNA106 Y B0 N1 VPW NCH W=1.82u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=1.82u L=0.06u
MNB2 N1 INT VSS VPW NCH W=1.82u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.78u L=0.06u
MPA108 Y B0 VDD VNW PCH W=1.52u L=0.06u
MPB1 Y A0 P1 VNW PCH W=2.8u L=0.06u
MPB2 P1 INT VDD VNW PCH W=2.8u L=0.06u
.ENDS	OAI2XB1X4MA10TR

****
.SUBCKT OAI2XB1X6MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.89u L=0.06u
MNA106 Y B0 N1 VPW NCH W=2.73u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=2.73u L=0.06u
MNB2 N1 INT VSS VPW NCH W=2.73u L=0.06u
MPA1 INT A1N VDD VNW PCH W=1.18u L=0.06u
MPA108 Y B0 VDD VNW PCH W=2.28u L=0.06u
MPB1 Y A0 P1 VNW PCH W=4.2u L=0.06u
MPB2 P1 INT VDD VNW PCH W=4.2u L=0.06u
.ENDS	OAI2XB1X6MA10TR

****
.SUBCKT OAI2XB1X8MA10TR  VDD VSS VPW VNW Y   A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=1.185u L=0.06u
MNA106 Y B0 N1 VPW NCH W=3.64u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=3.64u L=0.06u
MNB2 N1 INT VSS VPW NCH W=3.64u L=0.06u
MPA1 INT A1N VDD VNW PCH W=1.56u L=0.06u
MPA108 Y B0 VDD VNW PCH W=3.04u L=0.06u
MPB1 Y A0 P1 VNW PCH W=5.6u L=0.06u
MPB2 P1 INT VDD VNW PCH W=5.6u L=0.06u
.ENDS	OAI2XB1X8MA10TR

****
.SUBCKT OR2X0P5MA10TR  VDD VSS VPW VNW Y   A B
MNA1 INT A VSS VPW NCH W=0.15u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA2 INT B VSS VPW NCH W=0.15u L=0.06u
MPA1 INT A P1 VNW PCH W=0.38u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.38u L=0.06u
.ENDS	OR2X0P5MA10TR

****
.SUBCKT OR2X0P7MA10TR  VDD VSS VPW VNW Y   A B
MNA1 INT A VSS VPW NCH W=0.16u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.37u L=0.06u
MNA2 INT B VSS VPW NCH W=0.16u L=0.06u
MPA1 INT A P1 VNW PCH W=0.405u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.49u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.405u L=0.06u
.ENDS	OR2X0P7MA10TR

****

****
.SUBCKT OR2X1MA10TR  VDD VSS VPW VNW Y   A B
MNA1 INT A VSS VPW NCH W=0.205u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MNA2 INT B VSS VPW NCH W=0.205u L=0.06u
MPA1 INT A P1 VNW PCH W=0.52u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.52u L=0.06u
.ENDS	OR2X1MA10TR

****

****

****

****

****

****

****
.SUBCKT OR3X0P5MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=0.265u L=0.06u
MNA102 INT A VSS VPW NCH W=0.215u L=0.06u
MNA2 INT B VSS VPW NCH W=0.215u L=0.06u
MNA3 INT C VSS VPW NCH W=0.215u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.35u L=0.06u
MPA106 INT A P2 VNW PCH W=0.655u L=0.06u
MPA2 P2 B P1 VNW PCH W=0.655u L=0.06u
MPA3 P1 C VDD VNW PCH W=0.655u L=0.06u
.ENDS	OR3X0P5MA10TR

****

****

****

****
.SUBCKT OR3X2MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=1.06u L=0.06u
MNA102 INT A VSS VPW NCH W=0.6u L=0.06u
MNA2 INT B VSS VPW NCH W=0.6u L=0.06u
MNA3 INT C VSS VPW NCH W=0.6u L=0.06u
MPA1 Y INT VDD VNW PCH W=1.4u L=0.06u
MPA106 INT A P2 VNW PCH W=1.86u L=0.06u
MPA2 P2 B P1 VNW PCH W=1.86u L=0.06u
MPA3 P1 C VDD VNW PCH W=1.86u L=0.06u
.ENDS	OR3X2MA10TR

****
.SUBCKT OR3X3MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=1.59u L=0.06u
MNA102 INT A VSS VPW NCH W=0.92u L=0.06u
MNA2 INT B VSS VPW NCH W=0.92u L=0.06u
MNA3 INT C VSS VPW NCH W=0.92u L=0.06u
MPA1 Y INT VDD VNW PCH W=2.1u L=0.06u
MPA106 INT A P2 VNW PCH W=2.8u L=0.06u
MPA2 P2 B P1 VNW PCH W=2.8u L=0.06u
MPA3 P1 C VDD VNW PCH W=2.8u L=0.06u
.ENDS	OR3X3MA10TR

****
.SUBCKT OR3X4MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=2.12u L=0.06u
MNA102 INT A VSS VPW NCH W=1.2u L=0.06u
MNA2 INT B VSS VPW NCH W=1.2u L=0.06u
MNA3 INT C VSS VPW NCH W=1.2u L=0.06u
MPA1 Y INT VDD VNW PCH W=2.8u L=0.06u
MPA106 INT A P2 VNW PCH W=3.72u L=0.06u
MPA2 P2 B P1 VNW PCH W=3.72u L=0.06u
MPA3 P1 C VDD VNW PCH W=3.72u L=0.06u
.ENDS	OR3X4MA10TR

****
.SUBCKT OR3X6MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=3.18u L=0.06u
MNA102 INT A VSS VPW NCH W=1.8u L=0.06u
MNA2 INT B VSS VPW NCH W=1.8u L=0.06u
MNA3 INT C VSS VPW NCH W=1.8u L=0.06u
MPA1 Y INT VDD VNW PCH W=4.2u L=0.06u
MPA106 INT A P2 VNW PCH W=5.56u L=0.06u
MPA2 P2 B P1 VNW PCH W=5.56u L=0.06u
MPA3 P1 C VDD VNW PCH W=5.56u L=0.06u
.ENDS	OR3X6MA10TR

****
.SUBCKT OR3X8MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 Y INT VSS VPW NCH W=4.24u L=0.06u
MNA102 INT A VSS VPW NCH W=2.42u L=0.06u
MNA2 INT B VSS VPW NCH W=2.42u L=0.06u
MNA3 INT C VSS VPW NCH W=2.42u L=0.06u
MPA1 Y INT VDD VNW PCH W=5.6u L=0.06u
MPA106 INT A P2 VNW PCH W=7.425u L=0.06u
MPA2 P2 B P1 VNW PCH W=7.425u L=0.06u
MPA3 P1 C VDD VNW PCH W=7.425u L=0.06u
.ENDS	OR3X8MA10TR

****
.SUBCKT OR4X0P5MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 INT1 A VSS VPW NCH W=0.15u L=0.06u
MNA1012 Y INT1 N1 VPW NCH W=0.29u L=0.06u
MNA104 INT2 C VSS VPW NCH W=0.15u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.15u L=0.06u
MNA2014 N1 INT2 VSS VPW NCH W=0.29u L=0.06u
MNA206 INT2 D VSS VPW NCH W=0.15u L=0.06u
MPA1 INT1 A P1 VNW PCH W=0.37u L=0.06u
MPA1016 Y INT1 VDD VNW PCH W=0.24u L=0.06u
MPA108 INT2 C P1_3 VNW PCH W=0.37u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.37u L=0.06u
MPA2010 P1_3 D VDD VNW PCH W=0.37u L=0.06u
MPA2018 Y INT2 VDD VNW PCH W=0.24u L=0.06u
.ENDS	OR4X0P5MA10TR

****
.SUBCKT OR4X0P7MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 INT1 A VSS VPW NCH W=0.15u L=0.06u
MNA1012 Y INT1 N1 VPW NCH W=0.41u L=0.06u
MNA104 INT2 C VSS VPW NCH W=0.15u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.15u L=0.06u
MNA2014 N1 INT2 VSS VPW NCH W=0.41u L=0.06u
MNA206 INT2 D VSS VPW NCH W=0.15u L=0.06u
MPA1 INT1 A P1 VNW PCH W=0.37u L=0.06u
MPA1016 Y INT1 VDD VNW PCH W=0.34u L=0.06u
MPA108 INT2 C P1_3 VNW PCH W=0.37u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.37u L=0.06u
MPA2010 P1_3 D VDD VNW PCH W=0.37u L=0.06u
MPA2018 Y INT2 VDD VNW PCH W=0.34u L=0.06u
.ENDS	OR4X0P7MA10TR

****
.SUBCKT OR4X1MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 INT1 A VSS VPW NCH W=0.18u L=0.06u
MNA1012 Y INT1 N1 VPW NCH W=0.58u L=0.06u
MNA104 INT2 C VSS VPW NCH W=0.18u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.18u L=0.06u
MNA2014 N1 INT2 VSS VPW NCH W=0.58u L=0.06u
MNA206 INT2 D VSS VPW NCH W=0.18u L=0.06u
MPA1 INT1 A P1 VNW PCH W=0.44u L=0.06u
MPA1016 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MPA108 INT2 C P1_3 VNW PCH W=0.44u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.44u L=0.06u
MPA2010 P1_3 D VDD VNW PCH W=0.44u L=0.06u
MPA2018 Y INT2 VDD VNW PCH W=0.48u L=0.06u
.ENDS	OR4X1MA10TR

****
.SUBCKT OR4X1P4MA10TR  VDD VSS VPW VNW Y   A B C D
MNA1 INT1 A VSS VPW NCH W=0.25u L=0.06u
MNA1012 Y INT1 N1 VPW NCH W=0.82u L=0.06u
MNA104 INT2 C VSS VPW NCH W=0.25u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.25u L=0.06u
MNA2014 N1 INT2 VSS VPW NCH W=0.82u L=0.06u
MNA206 INT2 D VSS VPW NCH W=0.25u L=0.06u
MPA1 INT1 A P1 VNW PCH W=0.615u L=0.06u
MPA1016 Y INT1 VDD VNW PCH W=0.68u L=0.06u
MPA108 INT2 C P1_3 VNW PCH W=0.615u L=0.06u
MPA2 P1 B VDD VNW PCH W=0.615u L=0.06u
MPA2010 P1_3 D VDD VNW PCH W=0.615u L=0.06u
MPA2018 Y INT2 VDD VNW PCH W=0.68u L=0.06u
.ENDS	OR4X1P4MA10TR

****

****

****

****

****

****
.SUBCKT OR6X0P5MA10TR  VDD VSS VPW VNW Y   A B C D E F
MNA1 INT1 A VSS VPW NCH W=0.15u L=0.06u
MNA1018 Y INT1 N1 VPW NCH W=0.29u L=0.06u
MNA106 INT2 D VSS VPW NCH W=0.15u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.15u L=0.06u
MNA2020 N1 INT2 VSS VPW NCH W=0.29u L=0.06u
MNA208 INT2 E VSS VPW NCH W=0.15u L=0.06u
MNA3 INT1 C VSS VPW NCH W=0.15u L=0.06u
MNA3010 INT2 F VSS VPW NCH W=0.15u L=0.06u
MPA1 INT1 A P2 VNW PCH W=0.51u L=0.06u
MPA1012 INT2 D P2_6 VNW PCH W=0.51u L=0.06u
MPA1022 Y INT1 VDD VNW PCH W=0.24u L=0.06u
MPA2 P2 B P1 VNW PCH W=0.51u L=0.06u
MPA2014 P2_6 E P1_4 VNW PCH W=0.51u L=0.06u
MPA2024 Y INT2 VDD VNW PCH W=0.24u L=0.06u
MPA3 P1 C VDD VNW PCH W=0.51u L=0.06u
MPA3016 P1_4 F VDD VNW PCH W=0.51u L=0.06u
.ENDS	OR6X0P5MA10TR

****
.SUBCKT OR6X0P7MA10TR  VDD VSS VPW VNW Y   A B C D E F
MNA1 INT1 A VSS VPW NCH W=0.16u L=0.06u
MNA1018 Y INT1 N1 VPW NCH W=0.41u L=0.06u
MNA106 INT2 D VSS VPW NCH W=0.16u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.16u L=0.06u
MNA2020 N1 INT2 VSS VPW NCH W=0.41u L=0.06u
MNA208 INT2 E VSS VPW NCH W=0.16u L=0.06u
MNA3 INT1 C VSS VPW NCH W=0.16u L=0.06u
MNA3010 INT2 F VSS VPW NCH W=0.16u L=0.06u
MPA1 INT1 A P2 VNW PCH W=0.545u L=0.06u
MPA1012 INT2 D P2_6 VNW PCH W=0.545u L=0.06u
MPA1022 Y INT1 VDD VNW PCH W=0.34u L=0.06u
MPA2 P2 B P1 VNW PCH W=0.545u L=0.06u
MPA2014 P2_6 E P1_4 VNW PCH W=0.545u L=0.06u
MPA2024 Y INT2 VDD VNW PCH W=0.34u L=0.06u
MPA3 P1 C VDD VNW PCH W=0.545u L=0.06u
MPA3016 P1_4 F VDD VNW PCH W=0.545u L=0.06u
.ENDS	OR6X0P7MA10TR

****
.SUBCKT OR6X1MA10TR  VDD VSS VPW VNW Y   A B C D E F
MNA1 INT1 A VSS VPW NCH W=0.205u L=0.06u
MNA1018 Y INT1 N1 VPW NCH W=0.58u L=0.06u
MNA106 INT2 D VSS VPW NCH W=0.205u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.205u L=0.06u
MNA2020 N1 INT2 VSS VPW NCH W=0.58u L=0.06u
MNA208 INT2 E VSS VPW NCH W=0.205u L=0.06u
MNA3 INT1 C VSS VPW NCH W=0.205u L=0.06u
MNA3010 INT2 F VSS VPW NCH W=0.205u L=0.06u
MPA1 INT1 A P2 VNW PCH W=0.7u L=0.06u
MPA1012 INT2 D P2_6 VNW PCH W=0.7u L=0.06u
MPA1022 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MPA2 P2 B P1 VNW PCH W=0.7u L=0.06u
MPA2014 P2_6 E P1_4 VNW PCH W=0.7u L=0.06u
MPA2024 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MPA3 P1 C VDD VNW PCH W=0.7u L=0.06u
MPA3016 P1_4 F VDD VNW PCH W=0.7u L=0.06u
.ENDS	OR6X1MA10TR

****

****

****
.SUBCKT OR6X3MA10TR  VDD VSS VPW VNW Y   A B C D E F
MNA1 INT1 A VSS VPW NCH W=0.6u L=0.06u
MNA1018 Y INT1 N1 VPW NCH W=1.74u L=0.06u
MNA106 INT2 D VSS VPW NCH W=0.6u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.6u L=0.06u
MNA2020 N1 INT2 VSS VPW NCH W=1.74u L=0.06u
MNA208 INT2 E VSS VPW NCH W=0.6u L=0.06u
MNA3 INT1 C VSS VPW NCH W=0.6u L=0.06u
MNA3010 INT2 F VSS VPW NCH W=0.6u L=0.06u
MPA1 INT1 A P2 VNW PCH W=2.025u L=0.06u
MPA1012 INT2 D P2_6 VNW PCH W=2.025u L=0.06u
MPA1022 Y INT1 VDD VNW PCH W=1.44u L=0.06u
MPA2 P2 B P1 VNW PCH W=2.025u L=0.06u
MPA2014 P2_6 E P1_4 VNW PCH W=2.025u L=0.06u
MPA2024 Y INT2 VDD VNW PCH W=1.44u L=0.06u
MPA3 P1 C VDD VNW PCH W=2.025u L=0.06u
MPA3016 P1_4 F VDD VNW PCH W=2.025u L=0.06u
.ENDS	OR6X3MA10TR

****
.SUBCKT OR6X4MA10TR  VDD VSS VPW VNW Y   A B C D E F
MNA1 INT1 A VSS VPW NCH W=0.76u L=0.06u
MNA1018 Y INT1 N1 VPW NCH W=2.32u L=0.06u
MNA106 INT2 D VSS VPW NCH W=0.76u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.76u L=0.06u
MNA2020 N1 INT2 VSS VPW NCH W=2.32u L=0.06u
MNA208 INT2 E VSS VPW NCH W=0.76u L=0.06u
MNA3 INT1 C VSS VPW NCH W=0.76u L=0.06u
MNA3010 INT2 F VSS VPW NCH W=0.76u L=0.06u
MPA1 INT1 A P2 VNW PCH W=2.64u L=0.06u
MPA1012 INT2 D P2_6 VNW PCH W=2.64u L=0.06u
MPA1022 Y INT1 VDD VNW PCH W=1.92u L=0.06u
MPA2 P2 B P1 VNW PCH W=2.64u L=0.06u
MPA2014 P2_6 E P1_4 VNW PCH W=2.64u L=0.06u
MPA2024 Y INT2 VDD VNW PCH W=1.92u L=0.06u
MPA3 P1 C VDD VNW PCH W=2.64u L=0.06u
MPA3016 P1_4 F VDD VNW PCH W=2.64u L=0.06u
.ENDS	OR6X4MA10TR

****
.SUBCKT OR6X6MA10TR  VDD VSS VPW VNW Y   A B C D E F
MNA1 INT1 A VSS VPW NCH W=1.17u L=0.06u
MNA1018 Y INT1 N1 VPW NCH W=3.48u L=0.06u
MNA106 INT2 D VSS VPW NCH W=1.17u L=0.06u
MNA2 INT1 B VSS VPW NCH W=1.17u L=0.06u
MNA2020 N1 INT2 VSS VPW NCH W=3.48u L=0.06u
MNA208 INT2 E VSS VPW NCH W=1.17u L=0.06u
MNA3 INT1 C VSS VPW NCH W=1.17u L=0.06u
MNA3010 INT2 F VSS VPW NCH W=1.17u L=0.06u
MPA1 INT1 A P2 VNW PCH W=3.96u L=0.06u
MPA1012 INT2 D P2_6 VNW PCH W=3.96u L=0.06u
MPA1022 Y INT1 VDD VNW PCH W=2.88u L=0.06u
MPA2 P2 B P1 VNW PCH W=3.96u L=0.06u
MPA2014 P2_6 E P1_4 VNW PCH W=3.96u L=0.06u
MPA2024 Y INT2 VDD VNW PCH W=2.88u L=0.06u
MPA3 P1 C VDD VNW PCH W=3.96u L=0.06u
MPA3016 P1_4 F VDD VNW PCH W=3.96u L=0.06u
.ENDS	OR6X6MA10TR

****
.SUBCKT POSTICGX0P5BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.15u L=0.06u
MN1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.265u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.18u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.265u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.18u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.3u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.35u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.19u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX0P5BA10TR

****
.SUBCKT POSTICGX0P6BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.15u L=0.06u
MN1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.265u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.215u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.265u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.18u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.3u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.42u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.19u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX0P6BA10TR

****
.SUBCKT POSTICGX0P7BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.15u L=0.06u
MN1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.265u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.255u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.265u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.18u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.3u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.49u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.19u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX0P7BA10TR

****
.SUBCKT POSTICGX0P8BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.155u L=0.06u
MN1 N1 M VSS VPW NCH W=0.155u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.265u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.29u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.265u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.185u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.3u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.56u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.19u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX0P8BA10TR

****

****

****

****
.SUBCKT POSTICGX1BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.18u L=0.06u
MN1 N1 M VSS VPW NCH W=0.18u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.265u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.36u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.265u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.22u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.3u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.19u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX1BA10TR

****
.SUBCKT POSTICGX1P2BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.235u L=0.06u
MN1 N1 M VSS VPW NCH W=0.235u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.28u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.28u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.29u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.3u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.2u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX1P2BA10TR

****
.SUBCKT POSTICGX1P4BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.26u L=0.06u
MN1 N1 M VSS VPW NCH W=0.26u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.29u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.51u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.29u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.32u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.3u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.205u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.98u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.205u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX1P4BA10TR

****
.SUBCKT POSTICGX1P7BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.3u L=0.06u
MN1 N1 M VSS VPW NCH W=0.3u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.295u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.61u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.295u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.365u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.3u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.21u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=1.19u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.21u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX1P7BA10TR

****
.SUBCKT POSTICGX2BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.34u L=0.06u
MN1 N1 M VSS VPW NCH W=0.34u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.3u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.72u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.3u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.41u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.3u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.215u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=1.4u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.215u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX2BA10TR

****
.SUBCKT POSTICGX2P5BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.455u L=0.06u
MN1 N1 M VSS VPW NCH W=0.455u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.155u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.365u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.9u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.365u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.155u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.55u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.305u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.265u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=1.74u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.265u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.155u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX2P5BA10TR

****
.SUBCKT POSTICGX3BA10TR  VDD VSS VPW VNW ECK   CK E SEN
MN0 NOUT CK N1 VPW NCH W=0.52u L=0.06u
MN1 N1 M VSS VPW NCH W=0.52u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.16u L=0.06u
MNA1020 M NM N1_9 VPW NCH W=0.37u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=1.08u L=0.06u
MNA2 N1_9 SEN VSS VPW NCH W=0.37u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.16u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.63u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.31u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.27u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=2.1u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.27u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.16u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	POSTICGX3BA10TR

****

****

****

****

****

****

****
.SUBCKT PREICGX0P5BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.15u L=0.06u
MN1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.18u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.18u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.35u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX0P5BA10TR

****
.SUBCKT PREICGX0P6BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.15u L=0.06u
MN1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.215u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.18u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.42u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX0P6BA10TR

****
.SUBCKT PREICGX0P7BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.15u L=0.06u
MN1 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.255u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.18u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.49u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX0P7BA10TR

****
.SUBCKT PREICGX0P8BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.155u L=0.06u
MN1 N1 M VSS VPW NCH W=0.155u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.29u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.185u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.56u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX0P8BA10TR

****

****

****

****
.SUBCKT PREICGX1BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.18u L=0.06u
MN1 N1 M VSS VPW NCH W=0.18u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.36u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.22u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.19u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX1BA10TR

****
.SUBCKT PREICGX1P2BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.235u L=0.06u
MN1 N1 M VSS VPW NCH W=0.235u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.155u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.29u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.2u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX1P2BA10TR

****
.SUBCKT PREICGX1P4BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.26u L=0.06u
MN1 N1 M VSS VPW NCH W=0.26u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.16u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.51u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.32u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.205u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.98u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX1P4BA10TR

****
.SUBCKT PREICGX1P7BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.3u L=0.06u
MN1 N1 M VSS VPW NCH W=0.3u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.165u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.61u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.365u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.21u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=1.19u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX1P7BA10TR

****
.SUBCKT PREICGX2BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.34u L=0.06u
MN1 N1 M VSS VPW NCH W=0.34u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.17u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.15u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.72u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.15u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.15u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.41u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.215u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=1.4u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.15u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX2BA10TR

****
.SUBCKT PREICGX2P5BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.455u L=0.06u
MN1 N1 M VSS VPW NCH W=0.455u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.21u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.155u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.9u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.155u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.155u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.55u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.265u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=1.74u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.155u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX2P5BA10TR

****
.SUBCKT PREICGX3BA10TR  VDD VSS VPW VNW ECK   CK E SE
MN0 NOUT CK N1 VPW NCH W=0.52u L=0.06u
MN1 N1 M VSS VPW NCH W=0.52u L=0.06u
MNA1 N1_6 M VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.22u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.16u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=1.08u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.16u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.16u L=0.06u
MNOE05 NM CK N1_6 VPW NCH W=0.15u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.63u L=0.06u
MPA1 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.27u L=0.06u
MPA1023 NEN E P1_9 VNW PCH W=0.2u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=2.1u L=0.06u
MPA2 P1_9 SE VDD VNW PCH W=0.56u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.16u L=0.06u
MPOEN07 NM NCLK_ P1 VNW PCH W=0.15u L=0.06u
.ENDS	PREICGX3BA10TR

****

****

****

****

****

****

****
.SUBCKT RF1R1WSX1MA10TR  VDD VSS VPW VNW RBL   RWL WBL WWL
MNA1 NRDWL RWL VSS VPW NCH W=0.17u L=0.06u
MNA1016 NWRWL WWL VSS VPW NCH W=0.2u L=0.06u
MNA102 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NWRBL WBL VSS VPW NCH W=0.4u L=0.06u
MNA1024 RDBL_INT NM VSS VPW NCH W=0.51u L=0.06u
MNA108 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM WWL NWRBL VPW NCH W=0.4u L=0.06u
MNOE012 NM NWRWL N1 VPW NCH W=0.15u L=0.06u
MNOE028 RBL RWL RDBL_INT VPW NCH W=0.51u L=0.06u
MPA1 NRDWL RWL VDD VNW PCH W=0.23u L=0.06u
MPA1010 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1018 NWRWL WWL VDD VNW PCH W=0.27u L=0.06u
MPA1022 NWRBL WBL VDD VNW PCH W=0.6u L=0.06u
MPA1026 RDBL_INT NM VDD VNW PCH W=0.77u L=0.06u
MPA104 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NWRWL NWRBL VNW PCH W=0.4u L=0.06u
MPOEN014 NM WWL P1 VNW PCH W=0.15u L=0.06u
MPOEN030 RBL NRDWL RDBL_INT VNW PCH W=0.51u L=0.06u
.ENDS	RF1R1WSX1MA10TR

****
.SUBCKT RF1R1WSX1P4MA10TR  VDD VSS VPW VNW RBL   RWL WBL WWL
MNA1 NRDWL RWL VSS VPW NCH W=0.28u L=0.06u
MNA1016 NWRWL WWL VSS VPW NCH W=0.22u L=0.06u
MNA102 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NWRBL WBL VSS VPW NCH W=0.47u L=0.06u
MNA1024 RDBL_INT NM VSS VPW NCH W=0.72u L=0.06u
MNA108 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM WWL NWRBL VPW NCH W=0.47u L=0.06u
MNOE012 NM NWRWL N1 VPW NCH W=0.15u L=0.06u
MNOE028 RBL RWL RDBL_INT VPW NCH W=0.72u L=0.06u
MPA1 NRDWL RWL VDD VNW PCH W=0.38u L=0.06u
MPA1010 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1018 NWRWL WWL VDD VNW PCH W=0.3u L=0.06u
MPA1022 NWRBL WBL VDD VNW PCH W=0.7u L=0.06u
MPA1026 RDBL_INT NM VDD VNW PCH W=1.08u L=0.06u
MPA104 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NWRWL NWRBL VNW PCH W=0.47u L=0.06u
MPOEN014 NM WWL P1 VNW PCH W=0.15u L=0.06u
MPOEN030 RBL NRDWL RDBL_INT VNW PCH W=0.72u L=0.06u
.ENDS	RF1R1WSX1P4MA10TR

****
.SUBCKT RF1R1WSX2MA10TR  VDD VSS VPW VNW RBL   RWL WBL WWL
MNA1 NRDWL RWL VSS VPW NCH W=0.35u L=0.06u
MNA1016 NWRWL WWL VSS VPW NCH W=0.23u L=0.06u
MNA102 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1020 NWRBL WBL VSS VPW NCH W=0.51u L=0.06u
MNA1024 RDBL_INT NM VSS VPW NCH W=1.02u L=0.06u
MNA108 N1 M VSS VPW NCH W=0.15u L=0.06u
MNOE NM WWL NWRBL VPW NCH W=0.51u L=0.06u
MNOE012 NM NWRWL N1 VPW NCH W=0.15u L=0.06u
MNOE028 RBL RWL RDBL_INT VPW NCH W=1.02u L=0.06u
MPA1 NRDWL RWL VDD VNW PCH W=0.46u L=0.06u
MPA1010 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1018 NWRWL WWL VDD VNW PCH W=0.31u L=0.06u
MPA1022 NWRBL WBL VDD VNW PCH W=0.77u L=0.06u
MPA1026 RDBL_INT NM VDD VNW PCH W=1.54u L=0.06u
MPA104 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NWRWL NWRBL VNW PCH W=0.51u L=0.06u
MPOEN014 NM WWL P1 VNW PCH W=0.15u L=0.06u
MPOEN030 RBL NRDWL RDBL_INT VNW PCH W=1.02u L=0.06u
.ENDS	RF1R1WSX2MA10TR

****
.SUBCKT RF1R2WSX1MA10TR  VDD VSS VPW VNW RBL   RWL WBL1 WBL2 WWL1 WWL2
MN2 NET29 NWRWL2 NET32 VPW NCH W=0.2u L=0.06u
MN3 NET32 M VSS VPW NCH W=0.2u L=0.06u
MN4 NM NWRWL1 NET29 VPW NCH W=0.2u L=0.06u
MNA1 NRDWL RWL VSS VPW NCH W=0.17u L=0.06u
MNA1018 NWRWL2 WWL2 VSS VPW NCH W=0.2u L=0.06u
MNA1022 NWRWL1 WWL1 VSS VPW NCH W=0.2u L=0.06u
MNA1026 NWRBL2 WBL2 VSS VPW NCH W=0.4u L=0.06u
MNA1030 NWRBL1 WBL1 VSS VPW NCH W=0.4u L=0.06u
MNA1034 RDBL_INT NM VSS VPW NCH W=0.51u L=0.06u
MNA106 M NM VSS VPW NCH W=0.15u L=0.06u
MNOE NM WWL2 NWRBL2 VPW NCH W=0.4u L=0.06u
MNOE014 NM WWL1 NWRBL1 VPW NCH W=0.4u L=0.06u
MNOE038 RBL RWL RDBL_INT VPW NCH W=0.51u L=0.06u
MP2 NET39 WWL2 NET42 VNW PCH W=0.2u L=0.06u
MP3 NM WWL1 NET39 VNW PCH W=0.2u L=0.06u
MP5 NET42 M VDD VNW PCH W=0.2u L=0.06u
MPA1 NRDWL RWL VDD VNW PCH W=0.23u L=0.06u
MPA1020 NWRWL2 WWL2 VDD VNW PCH W=0.27u L=0.06u
MPA1024 NWRWL1 WWL1 VDD VNW PCH W=0.27u L=0.06u
MPA1028 NWRBL2 WBL2 VDD VNW PCH W=0.6u L=0.06u
MPA1032 NWRBL1 WBL1 VDD VNW PCH W=0.6u L=0.06u
MPA1036 RDBL_INT NM VDD VNW PCH W=0.77u L=0.06u
MPA108 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NWRWL2 NWRBL2 VNW PCH W=0.4u L=0.06u
MPOEN016 NM NWRWL1 NWRBL1 VNW PCH W=0.4u L=0.06u
MPOEN040 RBL NRDWL RDBL_INT VNW PCH W=0.51u L=0.06u
.ENDS	RF1R2WSX1MA10TR

****
.SUBCKT RF1R2WSX1P4MA10TR  VDD VSS VPW VNW RBL   RWL WBL1 WBL2 WWL1 WWL2
MN2 NET29 NWRWL2 NET32 VPW NCH W=0.2u L=0.06u
MN3 NET32 M VSS VPW NCH W=0.2u L=0.06u
MN4 NM NWRWL1 NET29 VPW NCH W=0.2u L=0.06u
MNA1 NRDWL RWL VSS VPW NCH W=0.28u L=0.06u
MNA1018 NWRWL2 WWL2 VSS VPW NCH W=0.22u L=0.06u
MNA1022 NWRWL1 WWL1 VSS VPW NCH W=0.22u L=0.06u
MNA1026 NWRBL2 WBL2 VSS VPW NCH W=0.4u L=0.06u
MNA1030 NWRBL1 WBL1 VSS VPW NCH W=0.4u L=0.06u
MNA1034 RDBL_INT NM VSS VPW NCH W=0.72u L=0.06u
MNA106 M NM VSS VPW NCH W=0.15u L=0.06u
MNOE NM WWL2 NWRBL2 VPW NCH W=0.47u L=0.06u
MNOE014 NM WWL1 NWRBL1 VPW NCH W=0.47u L=0.06u
MNOE038 RBL RWL RDBL_INT VPW NCH W=0.72u L=0.06u
MP2 NET39 WWL2 NET42 VNW PCH W=0.2u L=0.06u
MP3 NM WWL1 NET39 VNW PCH W=0.2u L=0.06u
MP5 NET42 M VDD VNW PCH W=0.2u L=0.06u
MPA1 NRDWL RWL VDD VNW PCH W=0.38u L=0.06u
MPA1020 NWRWL2 WWL2 VDD VNW PCH W=0.3u L=0.06u
MPA1024 NWRWL1 WWL1 VDD VNW PCH W=0.3u L=0.06u
MPA1028 NWRBL2 WBL2 VDD VNW PCH W=0.6u L=0.06u
MPA1032 NWRBL1 WBL1 VDD VNW PCH W=0.6u L=0.06u
MPA1036 RDBL_INT NM VDD VNW PCH W=1.08u L=0.06u
MPA108 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NWRWL2 NWRBL2 VNW PCH W=0.47u L=0.06u
MPOEN016 NM NWRWL1 NWRBL1 VNW PCH W=0.47u L=0.06u
MPOEN040 RBL NRDWL RDBL_INT VNW PCH W=0.72u L=0.06u
.ENDS	RF1R2WSX1P4MA10TR

****
.SUBCKT RF1R2WSX2MA10TR  VDD VSS VPW VNW RBL   RWL WBL1 WBL2 WWL1 WWL2
MN2 NET29 NWRWL2 NET32 VPW NCH W=0.2u L=0.06u
MN3 NET32 M VSS VPW NCH W=0.2u L=0.06u
MN4 NM NWRWL1 NET29 VPW NCH W=0.2u L=0.06u
MNA1 NRDWL RWL VSS VPW NCH W=0.35u L=0.06u
MNA1018 NWRWL2 WWL2 VSS VPW NCH W=0.23u L=0.06u
MNA1022 NWRWL1 WWL1 VSS VPW NCH W=0.23u L=0.06u
MNA1026 NWRBL2 WBL2 VSS VPW NCH W=0.4u L=0.06u
MNA1030 NWRBL1 WBL1 VSS VPW NCH W=0.4u L=0.06u
MNA1034 RDBL_INT NM VSS VPW NCH W=1.02u L=0.06u
MNA106 M NM VSS VPW NCH W=0.15u L=0.06u
MNOE NM WWL2 NWRBL2 VPW NCH W=0.51u L=0.06u
MNOE014 NM WWL1 NWRBL1 VPW NCH W=0.51u L=0.06u
MNOE038 RBL RWL RDBL_INT VPW NCH W=1.02u L=0.06u
MP2 NET39 WWL2 NET42 VNW PCH W=0.2u L=0.06u
MP3 NM WWL1 NET39 VNW PCH W=0.2u L=0.06u
MP5 NET42 M VDD VNW PCH W=0.2u L=0.06u
MPA1 NRDWL RWL VDD VNW PCH W=0.46u L=0.06u
MPA1020 NWRWL2 WWL2 VDD VNW PCH W=0.31u L=0.06u
MPA1024 NWRWL1 WWL1 VDD VNW PCH W=0.31u L=0.06u
MPA1028 NWRBL2 WBL2 VDD VNW PCH W=0.6u L=0.06u
MPA1032 NWRBL1 WBL1 VDD VNW PCH W=0.6u L=0.06u
MPA1036 RDBL_INT NM VDD VNW PCH W=1.54u L=0.06u
MPA108 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NWRWL2 NWRBL2 VNW PCH W=0.51u L=0.06u
MPOEN016 NM NWRWL1 NWRBL1 VNW PCH W=0.51u L=0.06u
MPOEN040 RBL NRDWL RDBL_INT VNW PCH W=1.02u L=0.06u
.ENDS	RF1R2WSX2MA10TR

****
.SUBCKT RF2R1WSX1MA10TR  VDD VSS VPW VNW RBL1 RBL2   RWL1 RWL2 WBL WWL
MNA1 NRDWL1 RWL1 VSS VPW NCH W=0.17u L=0.06u
MNA1016 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA102 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1024 NWRWL WWL VSS VPW NCH W=0.23u L=0.06u
MNA1028 NRDWL2 RWL2 VSS VPW NCH W=0.17u L=0.06u
MNA1032 NWRBL WBL VSS VPW NCH W=0.5u L=0.06u
MNA1036 RDBL1_INT NM VSS VPW NCH W=0.51u L=0.06u
MNA108 RDBL2_INT NM VSS VPW NCH W=0.51u L=0.06u
MNOE RBL2 RWL2 RDBL2_INT VPW NCH W=0.51u L=0.06u
MNOE012 NM WWL NWRBL VPW NCH W=0.5u L=0.06u
MNOE020 NM NWRWL N1 VPW NCH W=0.15u L=0.06u
MNOE040 RBL1 RWL1 RDBL1_INT VPW NCH W=0.51u L=0.06u
MPA1 NRDWL1 RWL1 VDD VNW PCH W=0.23u L=0.06u
MPA1010 RDBL2_INT NM VDD VNW PCH W=0.77u L=0.06u
MPA1018 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1026 NWRWL WWL VDD VNW PCH W=0.3u L=0.06u
MPA1030 NRDWL2 RWL2 VDD VNW PCH W=0.23u L=0.06u
MPA1034 NWRBL WBL VDD VNW PCH W=0.74u L=0.06u
MPA1038 RDBL1_INT NM VDD VNW PCH W=0.77u L=0.06u
MPA104 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN RBL2 NRDWL2 RDBL2_INT VNW PCH W=0.51u L=0.06u
MPOEN014 NM NWRWL NWRBL VNW PCH W=0.5u L=0.06u
MPOEN022 NM WWL P1 VNW PCH W=0.15u L=0.06u
MPOEN042 RBL1 NRDWL1 RDBL1_INT VNW PCH W=0.51u L=0.06u
.ENDS	RF2R1WSX1MA10TR

****
.SUBCKT RF2R1WSX1P4MA10TR  VDD VSS VPW VNW RBL1 RBL2   RWL1 RWL2 WBL WWL
MNA1 NRDWL1 RWL1 VSS VPW NCH W=0.28u L=0.06u
MNA1016 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA102 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1024 NWRWL WWL VSS VPW NCH W=0.23u L=0.06u
MNA1028 NRDWL2 RWL2 VSS VPW NCH W=0.28u L=0.06u
MNA1032 NWRBL WBL VSS VPW NCH W=0.5u L=0.06u
MNA1036 RDBL1_INT NM VSS VPW NCH W=0.72u L=0.06u
MNA108 RDBL2_INT NM VSS VPW NCH W=0.72u L=0.06u
MNOE RBL2 RWL2 RDBL2_INT VPW NCH W=0.72u L=0.06u
MNOE012 NM WWL NWRBL VPW NCH W=0.5u L=0.06u
MNOE020 NM NWRWL N1 VPW NCH W=0.15u L=0.06u
MNOE040 RBL1 RWL1 RDBL1_INT VPW NCH W=0.72u L=0.06u
MPA1 NRDWL1 RWL1 VDD VNW PCH W=0.38u L=0.06u
MPA1010 RDBL2_INT NM VDD VNW PCH W=1.08u L=0.06u
MPA1018 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1026 NWRWL WWL VDD VNW PCH W=0.31u L=0.06u
MPA1030 NRDWL2 RWL2 VDD VNW PCH W=0.38u L=0.06u
MPA1034 NWRBL WBL VDD VNW PCH W=0.75u L=0.06u
MPA1038 RDBL1_INT NM VDD VNW PCH W=1.08u L=0.06u
MPA104 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN RBL2 NRDWL2 RDBL2_INT VNW PCH W=0.72u L=0.06u
MPOEN014 NM NWRWL NWRBL VNW PCH W=0.5u L=0.06u
MPOEN022 NM WWL P1 VNW PCH W=0.15u L=0.06u
MPOEN042 RBL1 NRDWL1 RDBL1_INT VNW PCH W=0.72u L=0.06u
.ENDS	RF2R1WSX1P4MA10TR

****
.SUBCKT RF2R1WSX2MA10TR  VDD VSS VPW VNW RBL1 RBL2   RWL1 RWL2 WBL WWL
MNA1 NRDWL1 RWL1 VSS VPW NCH W=0.35u L=0.06u
MNA1016 N1 M VSS VPW NCH W=0.15u L=0.06u
MNA102 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1024 NWRWL WWL VSS VPW NCH W=0.24u L=0.06u
MNA1028 NRDWL2 RWL2 VSS VPW NCH W=0.35u L=0.06u
MNA1032 NWRBL WBL VSS VPW NCH W=0.47u L=0.06u
MNA1036 RDBL1_INT NM VSS VPW NCH W=1.02u L=0.06u
MNA108 RDBL2_INT NM VSS VPW NCH W=1.02u L=0.06u
MNOE RBL2 RWL2 RDBL2_INT VPW NCH W=1.02u L=0.06u
MNOE012 NM WWL NWRBL VPW NCH W=0.58u L=0.06u
MNOE020 NM NWRWL N1 VPW NCH W=0.15u L=0.06u
MNOE040 RBL1 RWL1 RDBL1_INT VPW NCH W=1.02u L=0.06u
MPA1 NRDWL1 RWL1 VDD VNW PCH W=0.46u L=0.06u
MPA1010 RDBL2_INT NM VDD VNW PCH W=1.54u L=0.06u
MPA1018 P1 M VDD VNW PCH W=0.15u L=0.06u
MPA1026 NWRWL WWL VDD VNW PCH W=0.32u L=0.06u
MPA1030 NRDWL2 RWL2 VDD VNW PCH W=0.46u L=0.06u
MPA1034 NWRBL WBL VDD VNW PCH W=0.7u L=0.06u
MPA1038 RDBL1_INT NM VDD VNW PCH W=1.54u L=0.06u
MPA104 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN RBL2 NRDWL2 RDBL2_INT VNW PCH W=1.02u L=0.06u
MPOEN014 NM NWRWL NWRBL VNW PCH W=0.58u L=0.06u
MPOEN022 NM WWL P1 VNW PCH W=0.15u L=0.06u
MPOEN042 RBL1 NRDWL1 RDBL1_INT VNW PCH W=1.02u L=0.06u
.ENDS	RF2R1WSX2MA10TR

****
.SUBCKT RF2R2WSX1MA10TR  VDD VSS VPW VNW RBL1 RBL2   RWL1 RWL2 WBL1 WBL2 WWL1 WWL2
MN2 NET29 NWRWL2 NET32 VPW NCH W=0.2u L=0.06u
MN3 NET32 M VSS VPW NCH W=0.2u L=0.06u
MN4 NM NWRWL1 NET29 VPW NCH W=0.2u L=0.06u
MNA1 NRDWL1 RWL1 VSS VPW NCH W=0.17u L=0.06u
MNA1011 RDBL2_INT NM VSS VPW NCH W=0.51u L=0.06u
MNA1018 NRDWL2 RWL2 VSS VPW NCH W=0.17u L=0.06u
MNA1026 NWRWL2 WWL2 VSS VPW NCH W=0.2u L=0.06u
MNA1030 NWRWL1 WWL1 VSS VPW NCH W=0.2u L=0.06u
MNA1034 NWRBL2 WBL2 VSS VPW NCH W=0.4u L=0.06u
MNA1038 NWRBL1 WBL1 VSS VPW NCH W=0.4u L=0.06u
MNA1042 RDBL1_INT NM VSS VPW NCH W=0.51u L=0.06u
MNA106 M NM VSS VPW NCH W=0.15u L=0.06u
MNOE NM WWL2 NWRBL2 VPW NCH W=0.4u L=0.06u
MNOE022 NM WWL1 NWRBL1 VPW NCH W=0.4u L=0.06u
MNOE046 RBL1 RWL1 RDBL1_INT VPW NCH W=0.51u L=0.06u
MNOE050 RBL2 RWL2 RDBL2_INT VPW NCH W=0.51u L=0.06u
MP2 NET39 WWL2 NET42 VNW PCH W=0.2u L=0.06u
MP3 NM WWL1 NET39 VNW PCH W=0.2u L=0.06u
MP5 NET42 M VDD VNW PCH W=0.2u L=0.06u
MPA1 NRDWL1 RWL1 VDD VNW PCH W=0.23u L=0.06u
MPA1013 RDBL2_INT NM VDD VNW PCH W=0.77u L=0.06u
MPA1020 NRDWL2 RWL2 VDD VNW PCH W=0.23u L=0.06u
MPA1028 NWRWL2 WWL2 VDD VNW PCH W=0.27u L=0.06u
MPA1032 NWRWL1 WWL1 VDD VNW PCH W=0.27u L=0.06u
MPA1036 NWRBL2 WBL2 VDD VNW PCH W=0.6u L=0.06u
MPA1040 NWRBL1 WBL1 VDD VNW PCH W=0.6u L=0.06u
MPA1044 RDBL1_INT NM VDD VNW PCH W=0.77u L=0.06u
MPA108 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NWRWL2 NWRBL2 VNW PCH W=0.4u L=0.06u
MPOEN024 NM NWRWL1 NWRBL1 VNW PCH W=0.4u L=0.06u
MPOEN048 RBL1 NRDWL1 RDBL1_INT VNW PCH W=0.51u L=0.06u
MPOEN052 RBL2 NRDWL2 RDBL2_INT VNW PCH W=0.51u L=0.06u
.ENDS	RF2R2WSX1MA10TR

****
.SUBCKT RF2R2WSX1P4MA10TR  VDD VSS VPW VNW RBL1 RBL2   RWL1 RWL2 WBL1 WBL2 WWL1 WWL2
MN2 NET29 NWRWL2 NET32 VPW NCH W=0.2u L=0.06u
MN3 NET32 M VSS VPW NCH W=0.2u L=0.06u
MN4 NM NWRWL1 NET29 VPW NCH W=0.2u L=0.06u
MNA1 NRDWL1 RWL1 VSS VPW NCH W=0.275u L=0.06u
MNA1011 RDBL2_INT NM VSS VPW NCH W=0.72u L=0.06u
MNA1018 NRDWL2 RWL2 VSS VPW NCH W=0.275u L=0.06u
MNA1026 NWRWL2 WWL2 VSS VPW NCH W=0.22u L=0.06u
MNA1030 NWRWL1 WWL1 VSS VPW NCH W=0.22u L=0.06u
MNA1034 NWRBL2 WBL2 VSS VPW NCH W=0.4u L=0.06u
MNA1038 NWRBL1 WBL1 VSS VPW NCH W=0.4u L=0.06u
MNA1042 RDBL1_INT NM VSS VPW NCH W=0.72u L=0.06u
MNA106 M NM VSS VPW NCH W=0.15u L=0.06u
MNOE NM WWL2 NWRBL2 VPW NCH W=0.47u L=0.06u
MNOE022 NM WWL1 NWRBL1 VPW NCH W=0.47u L=0.06u
MNOE046 RBL1 RWL1 RDBL1_INT VPW NCH W=0.72u L=0.06u
MNOE050 RBL2 RWL2 RDBL2_INT VPW NCH W=0.72u L=0.06u
MP2 NET39 WWL2 NET42 VNW PCH W=0.2u L=0.06u
MP3 NM WWL1 NET39 VNW PCH W=0.2u L=0.06u
MP5 NET42 M VDD VNW PCH W=0.2u L=0.06u
MPA1 NRDWL1 RWL1 VDD VNW PCH W=0.38u L=0.06u
MPA1013 RDBL2_INT NM VDD VNW PCH W=1.08u L=0.06u
MPA1020 NRDWL2 RWL2 VDD VNW PCH W=0.38u L=0.06u
MPA1028 NWRWL2 WWL2 VDD VNW PCH W=0.3u L=0.06u
MPA1032 NWRWL1 WWL1 VDD VNW PCH W=0.3u L=0.06u
MPA1036 NWRBL2 WBL2 VDD VNW PCH W=0.6u L=0.06u
MPA1040 NWRBL1 WBL1 VDD VNW PCH W=0.6u L=0.06u
MPA1044 RDBL1_INT NM VDD VNW PCH W=1.08u L=0.06u
MPA108 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NWRWL2 NWRBL2 VNW PCH W=0.47u L=0.06u
MPOEN024 NM NWRWL1 NWRBL1 VNW PCH W=0.47u L=0.06u
MPOEN048 RBL1 NRDWL1 RDBL1_INT VNW PCH W=0.72u L=0.06u
MPOEN052 RBL2 NRDWL2 RDBL2_INT VNW PCH W=0.72u L=0.06u
.ENDS	RF2R2WSX1P4MA10TR

****
.SUBCKT RF2R2WSX2MA10TR  VDD VSS VPW VNW RBL1 RBL2   RWL1 RWL2 WBL1 WBL2 WWL1 WWL2
MN2 NET29 NWRWL2 NET32 VPW NCH W=0.2u L=0.06u
MN3 NET32 M VSS VPW NCH W=0.2u L=0.06u
MN4 NM NWRWL1 NET29 VPW NCH W=0.2u L=0.06u
MNA1 NRDWL1 RWL1 VSS VPW NCH W=0.35u L=0.06u
MNA1011 RDBL2_INT NM VSS VPW NCH W=1.02u L=0.06u
MNA1018 NRDWL2 RWL2 VSS VPW NCH W=0.35u L=0.06u
MNA1026 NWRWL2 WWL2 VSS VPW NCH W=0.24u L=0.06u
MNA1030 NWRWL1 WWL1 VSS VPW NCH W=0.24u L=0.06u
MNA1034 NWRBL2 WBL2 VSS VPW NCH W=0.4u L=0.06u
MNA1038 NWRBL1 WBL1 VSS VPW NCH W=0.4u L=0.06u
MNA1042 RDBL1_INT NM VSS VPW NCH W=1.02u L=0.06u
MNA106 M NM VSS VPW NCH W=0.15u L=0.06u
MNOE NM WWL2 NWRBL2 VPW NCH W=0.57u L=0.06u
MNOE022 NM WWL1 NWRBL1 VPW NCH W=0.57u L=0.06u
MNOE046 RBL1 RWL1 RDBL1_INT VPW NCH W=1.02u L=0.06u
MNOE050 RBL2 RWL2 RDBL2_INT VPW NCH W=1.02u L=0.06u
MP2 NET39 WWL2 NET42 VNW PCH W=0.2u L=0.06u
MP3 NM WWL1 NET39 VNW PCH W=0.2u L=0.06u
MP5 NET42 M VDD VNW PCH W=0.2u L=0.06u
MPA1 NRDWL1 RWL1 VDD VNW PCH W=0.46u L=0.06u
MPA1013 RDBL2_INT NM VDD VNW PCH W=1.54u L=0.06u
MPA1020 NRDWL2 RWL2 VDD VNW PCH W=0.46u L=0.06u
MPA1028 NWRWL2 WWL2 VDD VNW PCH W=0.32u L=0.06u
MPA1032 NWRWL1 WWL1 VDD VNW PCH W=0.32u L=0.06u
MPA1036 NWRBL2 WBL2 VDD VNW PCH W=0.6u L=0.06u
MPA1040 NWRBL1 WBL1 VDD VNW PCH W=0.6u L=0.06u
MPA1044 RDBL1_INT NM VDD VNW PCH W=1.54u L=0.06u
MPA108 M NM VDD VNW PCH W=0.15u L=0.06u
MPOEN NM NWRWL2 NWRBL2 VNW PCH W=0.57u L=0.06u
MPOEN024 NM NWRWL1 NWRBL1 VNW PCH W=0.57u L=0.06u
MPOEN048 RBL1 NRDWL1 RDBL1_INT VNW PCH W=1.02u L=0.06u
MPOEN052 RBL2 NRDWL2 RDBL2_INT VNW PCH W=1.02u L=0.06u
.ENDS	RF2R2WSX2MA10TR

****
.SUBCKT SDFFNQX1MA10TR  VDD VSS VPW VNW Q   CKN D SE SI
MN0 NMUX D N1 VPW NCH W=0.25u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.25u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.15u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.3u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.2u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.35u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.15u L=0.06u
MNOE017 S BCLK_ N1_10 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK_ N1_14 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM BCLK_ NMUX VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.55u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.55u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.35u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.45u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.25u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.45u L=0.06u
MPOEN019 S NCLK_ P1_12 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK_ P1_16 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.2u L=0.06u
MPOEN046 NM NCLK_ NMUX VNW PCH W=0.45u L=0.06u
.ENDS	SDFFNQX1MA10TR

****
.SUBCKT SDFFNQX2MA10TR  VDD VSS VPW VNW Q   CKN D SE SI
MN0 NMUX D N1 VPW NCH W=0.35u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.35u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.16u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.24u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.58u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.2u L=0.06u
MNOE017 S BCLK_ N1_10 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK_ N1_14 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM BCLK_ NMUX VPW NCH W=0.2u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.7u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.7u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.32u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.58u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.6u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.3u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.6u L=0.06u
MPOEN019 S NCLK_ P1_12 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK_ P1_16 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.2u L=0.06u
MPOEN046 NM NCLK_ NMUX VNW PCH W=0.6u L=0.06u
.ENDS	SDFFNQX2MA10TR

****
.SUBCKT SDFFNQX3MA10TR  VDD VSS VPW VNW Q   CKN D SE SI
MN0 NMUX D N1 VPW NCH W=0.35u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.35u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.18u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.45u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.28u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA108 NS S VSS VPW NCH W=0.58u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.25u L=0.06u
MNOE017 S BCLK_ N1_10 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK_ N1_14 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM BCLK_ NMUX VPW NCH W=0.25u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.7u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.7u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.36u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.58u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.34u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.7u L=0.06u
MPOEN019 S NCLK_ P1_12 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK_ P1_16 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.2u L=0.06u
MPOEN046 NM NCLK_ NMUX VNW PCH W=0.7u L=0.06u
.ENDS	SDFFNQX3MA10TR

****
.SUBCKT SDFFNRPQX1MA10TR  VDD VSS VPW VNW Q   CKN R D SE SI
MN0 NMUX D N1 VPW NCH W=0.25u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.25u L=0.06u
MN2 NET47 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.15u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.15u L=0.06u
MNA1018 M R VSS VPW NCH W=0.25u L=0.06u
MNA1028 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.2u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.36u L=0.06u
MNA2 M NM VSS VPW NCH W=0.25u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.15u L=0.06u
MNOE032 NM NCLK_ N1_15 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE044 NM BCLK_ NMUX VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.55u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.55u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.36u L=0.06u
MPA1021 M R P1_13 VNW PCH W=0.6u L=0.06u
MPA1030 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.25u L=0.06u
MPA2 P1_13 NM VDD VNW PCH W=0.6u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.445u L=0.06u
MPOEN034 NM BCLK_ P1_17 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN046 NM NCLK_ NMUX VNW PCH W=0.45u L=0.06u
.ENDS	SDFFNRPQX1MA10TR

****
.SUBCKT SDFFNRPQX2MA10TR  VDD VSS VPW VNW Q   CKN R D SE SI
MN0 NMUX D N1 VPW NCH W=0.35u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.35u L=0.06u
MN2 NET47 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.15u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.16u L=0.06u
MNA1018 M R VSS VPW NCH W=0.3u L=0.06u
MNA1028 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.24u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.58u L=0.06u
MNA2 M NM VSS VPW NCH W=0.3u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.2u L=0.06u
MNOE032 NM NCLK_ N1_15 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE044 NM BCLK_ NMUX VPW NCH W=0.2u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.7u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.7u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.32u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.58u L=0.06u
MPA1021 M R P1_13 VNW PCH W=0.8u L=0.06u
MPA1030 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.3u L=0.06u
MPA2 P1_13 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.6u L=0.06u
MPOEN034 NM BCLK_ P1_17 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN046 NM NCLK_ NMUX VNW PCH W=0.6u L=0.06u
.ENDS	SDFFNRPQX2MA10TR

****
.SUBCKT SDFFNRPQX3MA10TR  VDD VSS VPW VNW Q   CKN R D SE SI
MN5 NMUX D N1 VPW NCH W=0.35u L=0.06u
MN6 N1 NSE VSS VPW NCH W=0.35u L=0.06u
MN7 S R VSS VPW NCH W=0.15u L=0.06u
MN8 S BCLK_ NET49 VPW NCH W=0.15u L=0.06u
MN9 NET49 NS VSS VPW NCH W=0.15u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.18u L=0.06u
MNA1010 M R VSS VPW NCH W=0.3u L=0.06u
MNA102 BCLK_ NCLK_ VSS VPW NCH W=0.28u L=0.06u
MNA1025 N1_15 SI VSS VPW NCH W=0.15u L=0.06u
MNA1031 N1_19 M VSS VPW NCH W=0.15u L=0.06u
MNA1047 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1051 NS S VSS VPW NCH W=0.58u L=0.06u
MNA106 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA2 M NM VSS VPW NCH W=0.3u L=0.06u
MNOE NMUX SE N1_15 VPW NCH W=0.15u L=0.06u
MNOE035 NM NCLK_ N1_19 VPW NCH W=0.15u L=0.06u
MNOE039 NM BCLK_ NMUX VPW NCH W=0.25u L=0.06u
MNOE043 S NCLK_ M VPW NCH W=0.25u L=0.06u
MP10 NET69 NS NET63 VNW PCH W=0.2u L=0.06u
MP6 P1 SE VDD VNW PCH W=0.7u L=0.06u
MP7 NMUX D P1 VNW PCH W=0.7u L=0.06u
MP8 S NCLK_ NET69 VNW PCH W=0.2u L=0.06u
MP9 NET63 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.36u L=0.06u
MPA1013 M R P1_13 VNW PCH W=0.8u L=0.06u
MPA1027 P1_17 SI VDD VNW PCH W=0.2u L=0.06u
MPA1033 P1_21 M VDD VNW PCH W=0.15u L=0.06u
MPA104 BCLK_ NCLK_ VDD VNW PCH W=0.34u L=0.06u
MPA1049 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1053 NS S VDD VNW PCH W=0.58u L=0.06u
MPA108 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA2 P1_13 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN NMUX NSE P1_17 VNW PCH W=0.2u L=0.06u
MPOEN037 NM BCLK_ P1_21 VNW PCH W=0.15u L=0.06u
MPOEN041 NM NCLK_ NMUX VNW PCH W=0.7u L=0.06u
MPOEN045 S BCLK_ M VNW PCH W=0.7u L=0.06u
.ENDS	SDFFNRPQX3MA10TR

****
.SUBCKT SDFFNSQX1MA10TR  VDD VSS VPW VNW Q   CKN D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.25u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.25u L=0.06u
MN2 NET50 NS NET47 VPW NCH W=0.2u L=0.06u
MN3 NET47 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET50 VPW NCH W=0.2u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.15u L=0.06u
MNA1022 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1030 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.2u L=0.06u
MNA1042 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1046 M SN N1_21 VPW NCH W=0.5u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.37u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.5u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK_ N1_13 VPW NCH W=0.15u L=0.06u
MNOE034 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE038 NM BCLK_ NMUX VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.55u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.55u L=0.06u
MP2 NET58 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.37u L=0.06u
MPA1024 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1044 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1049 M SN VDD VNW PCH W=0.45u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.25u L=0.06u
MPA2 M NM VDD VNW PCH W=0.45u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.45u L=0.06u
MPOEN028 NM BCLK_ P1_15 VNW PCH W=0.15u L=0.06u
MPOEN036 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN040 NM NCLK_ NMUX VNW PCH W=0.45u L=0.06u
.ENDS	SDFFNSQX1MA10TR

****
.SUBCKT SDFFNSQX2MA10TR  VDD VSS VPW VNW Q   CKN D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.35u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.35u L=0.06u
MN2 NET50 NS NET47 VPW NCH W=0.2u L=0.06u
MN3 NET47 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET50 VPW NCH W=0.2u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.16u L=0.06u
MNA1022 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1030 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.24u L=0.06u
MNA1042 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1046 M SN N1_21 VPW NCH W=0.6u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.58u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.6u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.2u L=0.06u
MNOE026 NM NCLK_ N1_13 VPW NCH W=0.15u L=0.06u
MNOE034 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE038 NM BCLK_ NMUX VPW NCH W=0.2u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.7u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.7u L=0.06u
MP2 NET58 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.32u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.58u L=0.06u
MPA1024 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1044 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1049 M SN VDD VNW PCH W=0.5u L=0.06u
MPA1054 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.3u L=0.06u
MPA2 M NM VDD VNW PCH W=0.5u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.6u L=0.06u
MPOEN028 NM BCLK_ P1_15 VNW PCH W=0.15u L=0.06u
MPOEN036 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN040 NM NCLK_ NMUX VNW PCH W=0.6u L=0.06u
.ENDS	SDFFNSQX2MA10TR

****
.SUBCKT SDFFNSQX3MA10TR  VDD VSS VPW VNW Q   CKN D SE SN SI
MN5 NMUX D N1 VPW NCH W=0.35u L=0.06u
MN6 N1 NSE VSS VPW NCH W=0.35u L=0.06u
MN7 NET55 SN VSS VPW NCH W=0.2u L=0.06u
MN8 NET52 NS NET55 VPW NCH W=0.2u L=0.06u
MN9 S BCLK_ NET52 VPW NCH W=0.2u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.18u L=0.06u
MNA102 BCLK_ NCLK_ VSS VPW NCH W=0.28u L=0.06u
MNA1020 N1_13 SI VSS VPW NCH W=0.15u L=0.06u
MNA1026 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1042 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1046 NS S VSS VPW NCH W=0.58u L=0.06u
MNA1050 M SN N1_21 VPW NCH W=0.6u L=0.06u
MNA106 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.6u L=0.06u
MNOE NMUX SE N1_13 VPW NCH W=0.15u L=0.06u
MNOE030 NM NCLK_ N1_17 VPW NCH W=0.15u L=0.06u
MNOE034 NM BCLK_ NMUX VPW NCH W=0.25u L=0.06u
MNOE038 S NCLK_ M VPW NCH W=0.25u L=0.06u
MP5 NET66 NS VDD VNW PCH W=0.2u L=0.06u
MP6 P1 SE VDD VNW PCH W=0.7u L=0.06u
MP7 NMUX D P1 VNW PCH W=0.7u L=0.06u
MP8 S NCLK_ NET66 VNW PCH W=0.2u L=0.06u
MP9 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.36u L=0.06u
MPA1022 P1_15 SI VDD VNW PCH W=0.2u L=0.06u
MPA1028 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA104 BCLK_ NCLK_ VDD VNW PCH W=0.34u L=0.06u
MPA1044 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1048 NS S VDD VNW PCH W=0.58u L=0.06u
MPA1053 M SN VDD VNW PCH W=0.5u L=0.06u
MPA108 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA2 M NM VDD VNW PCH W=0.5u L=0.06u
MPOEN NMUX NSE P1_15 VNW PCH W=0.2u L=0.06u
MPOEN032 NM BCLK_ P1_19 VNW PCH W=0.15u L=0.06u
MPOEN036 NM NCLK_ NMUX VNW PCH W=0.7u L=0.06u
MPOEN040 S BCLK_ M VNW PCH W=0.7u L=0.06u
.ENDS	SDFFNSQX3MA10TR

****
.SUBCKT SDFFNSRPQX1MA10TR  VDD VSS VPW VNW Q   CKN R D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.25u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.25u L=0.06u
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.3u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.3u L=0.06u
MN9 M R NET046 VPW NCH W=0.3u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.15u L=0.06u
MNA1031 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1039 N1_21 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.2u L=0.06u
MNA1051 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1055 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.37u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.15u L=0.06u
MNOE035 NM NCLK_ N1_17 VPW NCH W=0.15u L=0.06u
MNOE043 NMUX SE N1_21 VPW NCH W=0.15u L=0.06u
MNOE047 NM BCLK_ NMUX VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.55u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.55u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.45u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.45u L=0.06u
MP9 M SN VDD VNW PCH W=0.45u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.37u L=0.06u
MPA1033 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA1041 P1_23 SI VDD VNW PCH W=0.2u L=0.06u
MPA1053 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1057 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.25u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.45u L=0.06u
MPOEN037 NM BCLK_ P1_19 VNW PCH W=0.15u L=0.06u
MPOEN045 NMUX NSE P1_23 VNW PCH W=0.2u L=0.06u
MPOEN049 NM NCLK_ NMUX VNW PCH W=0.45u L=0.06u
.ENDS	SDFFNSRPQX1MA10TR

****
.SUBCKT SDFFNSRPQX2MA10TR  VDD VSS VPW VNW Q   CKN R D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.3u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.3u L=0.06u
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.4u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.4u L=0.06u
MN9 M R NET046 VPW NCH W=0.4u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.16u L=0.06u
MNA1031 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1039 N1_21 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK_ NCLK_ VSS VPW NCH W=0.24u L=0.06u
MNA1051 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1055 Q NS VSS VPW NCH W=1.06u L=0.06u
MNA108 NS S VSS VPW NCH W=0.52u L=0.06u
MNOE S NCLK_ M VPW NCH W=0.2u L=0.06u
MNOE035 NM NCLK_ N1_17 VPW NCH W=0.15u L=0.06u
MNOE043 NMUX SE N1_21 VPW NCH W=0.15u L=0.06u
MNOE047 NM BCLK_ NMUX VPW NCH W=0.2u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.7u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.7u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.6u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.6u L=0.06u
MP9 M SN VDD VNW PCH W=0.6u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.32u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.52u L=0.06u
MPA1033 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA1041 P1_23 SI VDD VNW PCH W=0.2u L=0.06u
MPA1053 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1057 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK_ NCLK_ VDD VNW PCH W=0.3u L=0.06u
MPOEN S BCLK_ M VNW PCH W=0.6u L=0.06u
MPOEN037 NM BCLK_ P1_19 VNW PCH W=0.15u L=0.06u
MPOEN045 NMUX NSE P1_23 VNW PCH W=0.2u L=0.06u
MPOEN049 NM NCLK_ NMUX VNW PCH W=0.6u L=0.06u
.ENDS	SDFFNSRPQX2MA10TR

****
.SUBCKT SDFFNSRPQX3MA10TR  VDD VSS VPW VNW Q   CKN R D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.3u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.3u L=0.06u
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S BCLK_ NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.4u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.4u L=0.06u
MN9 M R NET046 VPW NCH W=0.4u L=0.06u
MNA1 NCLK_ CKN VSS VPW NCH W=0.18u L=0.06u
MNA1031 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1039 N1_21 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA1047 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1055 NS S VSS VPW NCH W=0.58u L=0.06u
MNA109 BCLK_ NCLK_ VSS VPW NCH W=0.28u L=0.06u
MNOE NM BCLK_ NMUX VPW NCH W=0.25u L=0.06u
MNOE035 NM NCLK_ N1_17 VPW NCH W=0.15u L=0.06u
MNOE043 NMUX SE N1_21 VPW NCH W=0.15u L=0.06u
MNOE051 S NCLK_ M VPW NCH W=0.25u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.7u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.7u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S NCLK_ NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.6u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.6u L=0.06u
MP9 M SN VDD VNW PCH W=0.6u L=0.06u
MPA1 NCLK_ CKN VDD VNW PCH W=0.36u L=0.06u
MPA1011 BCLK_ NCLK_ VDD VNW PCH W=0.34u L=0.06u
MPA1033 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA1041 P1_23 SI VDD VNW PCH W=0.2u L=0.06u
MPA1049 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1057 NS S VDD VNW PCH W=0.58u L=0.06u
MPA106 Q NS VDD VNW PCH W=2.1u L=0.06u
MPOEN NM NCLK_ NMUX VNW PCH W=0.7u L=0.06u
MPOEN037 NM BCLK_ P1_19 VNW PCH W=0.15u L=0.06u
MPOEN045 NMUX NSE P1_23 VNW PCH W=0.2u L=0.06u
MPOEN053 S BCLK_ M VNW PCH W=0.7u L=0.06u
.ENDS	SDFFNSRPQX3MA10TR

****
.SUBCKT SDFFQNX0P5MA10TR  VDD VSS VPW VNW QN   CK D SE SI
MN2 NMUX D N1 VPW NCH W=0.26u L=0.06u
MN3 N1 NSE VSS VPW NCH W=0.26u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_18 M VSS VPW NCH W=0.15u L=0.06u
MNA102 N1_10 SI VSS VPW NCH W=0.15u L=0.06u
MNA1036 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1048 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1052 QN S VSS VPW NCH W=0.28u L=0.06u
MNA109 N1_14 NS VSS VPW NCH W=0.15u L=0.06u
MNOE NMUX SE N1_10 VPW NCH W=0.15u L=0.06u
MNOE013 S NCLK N1_14 VPW NCH W=0.15u L=0.06u
MNOE022 NM BCLK N1_18 VPW NCH W=0.15u L=0.06u
MNOE027 NM NCLK NMUX VPW NCH W=0.15u L=0.06u
MNOE032 S BCLK M VPW NCH W=0.15u L=0.06u
MP2 P1 SE VDD VNW PCH W=0.29u L=0.06u
MP3 NMUX D P1 VNW PCH W=0.29u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1011 P1_16 NS VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_20 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA104 P1_12 SI VDD VNW PCH W=0.15u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1050 M NM VDD VNW PCH W=0.22u L=0.06u
MPA1054 QN S VDD VNW PCH W=0.37u L=0.06u
MPOEN NMUX NSE P1_12 VNW PCH W=0.15u L=0.06u
MPOEN015 S BCLK P1_16 VNW PCH W=0.15u L=0.06u
MPOEN024 NM NCLK P1_20 VNW PCH W=0.15u L=0.06u
MPOEN029 NM BCLK NMUX VNW PCH W=0.15u L=0.06u
MPOEN034 S NCLK M VNW PCH W=0.15u L=0.06u
.ENDS	SDFFQNX0P5MA10TR

****
.SUBCKT SDFFQNX1MA10TR  VDD VSS VPW VNW QN   CK D SE SI
MN2 NMUX D N1 VPW NCH W=0.4u L=0.06u
MN3 N1 NSE VSS VPW NCH W=0.4u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1010 N1_14 NS VSS VPW NCH W=0.15u L=0.06u
MNA1019 N1_18 M VSS VPW NCH W=0.15u L=0.06u
MNA103 N1_10 SI VSS VPW NCH W=0.15u L=0.06u
MNA1036 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1048 M NM VSS VPW NCH W=0.32u L=0.06u
MNA1052 QN S VSS VPW NCH W=0.53u L=0.06u
MNOE NMUX SE N1_10 VPW NCH W=0.15u L=0.06u
MNOE014 S NCLK N1_14 VPW NCH W=0.15u L=0.06u
MNOE023 NM BCLK N1_18 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MNOE032 S BCLK M VPW NCH W=0.28u L=0.06u
MP2 P1 SE VDD VNW PCH W=0.48u L=0.06u
MP3 NMUX D P1 VNW PCH W=0.48u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1012 P1_16 NS VDD VNW PCH W=0.15u L=0.06u
MPA1021 P1_20 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA105 P1_12 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 M NM VDD VNW PCH W=0.5u L=0.06u
MPA1054 QN S VDD VNW PCH W=0.7u L=0.06u
MPOEN NMUX NSE P1_12 VNW PCH W=0.2u L=0.06u
MPOEN016 S BCLK P1_16 VNW PCH W=0.15u L=0.06u
MPOEN025 NM NCLK P1_20 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NMUX VNW PCH W=0.28u L=0.06u
MPOEN034 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	SDFFQNX1MA10TR

****
.SUBCKT SDFFQNX2MA10TR  VDD VSS VPW VNW QN   CK D SE SI
MN2 NMUX D N1 VPW NCH W=0.57u L=0.06u
MN3 N1 NSE VSS VPW NCH W=0.57u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1010 N1_14 NS VSS VPW NCH W=0.15u L=0.06u
MNA1019 N1_18 M VSS VPW NCH W=0.15u L=0.06u
MNA103 N1_10 SI VSS VPW NCH W=0.15u L=0.06u
MNA1036 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1048 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1052 QN S VSS VPW NCH W=1.06u L=0.06u
MNOE NMUX SE N1_10 VPW NCH W=0.15u L=0.06u
MNOE014 S NCLK N1_14 VPW NCH W=0.15u L=0.06u
MNOE023 NM BCLK N1_18 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MNOE032 S BCLK M VPW NCH W=0.4u L=0.06u
MP2 P1 SE VDD VNW PCH W=0.63u L=0.06u
MP3 NMUX D P1 VNW PCH W=0.63u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1012 P1_16 NS VDD VNW PCH W=0.15u L=0.06u
MPA1021 P1_20 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA105 P1_12 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 M NM VDD VNW PCH W=0.56u L=0.06u
MPA1054 QN S VDD VNW PCH W=1.4u L=0.06u
MPOEN NMUX NSE P1_12 VNW PCH W=0.2u L=0.06u
MPOEN016 S BCLK P1_16 VNW PCH W=0.15u L=0.06u
MPOEN025 NM NCLK P1_20 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
MPOEN034 S NCLK M VNW PCH W=0.4u L=0.06u
.ENDS	SDFFQNX2MA10TR

****
.SUBCKT SDFFQNX3MA10TR  VDD VSS VPW VNW QN   CK D SE SI
MN2 NMUX D N1 VPW NCH W=0.57u L=0.06u
MN3 N1 NSE VSS VPW NCH W=0.57u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1010 N1_14 NS VSS VPW NCH W=0.15u L=0.06u
MNA1019 N1_18 M VSS VPW NCH W=0.15u L=0.06u
MNA103 N1_10 SI VSS VPW NCH W=0.15u L=0.06u
MNA1036 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1048 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1052 QN S VSS VPW NCH W=1.59u L=0.06u
MNOE NMUX SE N1_10 VPW NCH W=0.15u L=0.06u
MNOE014 S NCLK N1_14 VPW NCH W=0.15u L=0.06u
MNOE023 NM BCLK N1_18 VPW NCH W=0.15u L=0.06u
MNOE028 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE032 S BCLK M VPW NCH W=0.58u L=0.06u
MP2 P1 SE VDD VNW PCH W=0.63u L=0.06u
MP3 NMUX D P1 VNW PCH W=0.63u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1012 P1_16 NS VDD VNW PCH W=0.15u L=0.06u
MPA1021 P1_20 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA105 P1_12 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1054 QN S VDD VNW PCH W=2.1u L=0.06u
MPOEN NMUX NSE P1_12 VNW PCH W=0.2u L=0.06u
MPOEN016 S BCLK P1_16 VNW PCH W=0.15u L=0.06u
MPOEN025 NM NCLK P1_20 VNW PCH W=0.15u L=0.06u
MPOEN030 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN034 S NCLK M VNW PCH W=0.58u L=0.06u
.ENDS	SDFFQNX3MA10TR

****
.SUBCKT SDFFQX0P5MA10TR  VDD VSS VPW VNW Q   CK D SE SI
MN0 NMUX D N1 VPW NCH W=0.26u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.26u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.31u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE017 S NCLK N1_10 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_14 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.29u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.29u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.25u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.22u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.15u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN019 S BCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_16 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.15u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.15u L=0.06u
.ENDS	SDFFQX0P5MA10TR

****
.SUBCKT SDFFQX1MA10TR  VDD VSS VPW VNW Q   CK D SE SI
MN0 NMUX D N1 VPW NCH W=0.4u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.4u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.28u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA108 NS S VSS VPW NCH W=0.3u L=0.06u
MNOE S BCLK M VPW NCH W=0.28u L=0.06u
MNOE017 S NCLK N1_10 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_14 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.48u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.48u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.47u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.4u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPOEN S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN019 S BCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_16 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.2u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.28u L=0.06u
.ENDS	SDFFQX1MA10TR

****
.SUBCKT SDFFQX2MA10TR  VDD VSS VPW VNW Q   CK D SE SI
MN0 NMUX D N1 VPW NCH W=0.58u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.58u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.46u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE017 S NCLK N1_10 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_14 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.62u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.62u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.57u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN019 S BCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_16 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.2u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
.ENDS	SDFFQX2MA10TR

****
.SUBCKT SDFFQX3MA10TR  VDD VSS VPW VNW Q   CK D SE SI
MN0 NMUX D N1 VPW NCH W=0.58u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.58u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.51u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA108 NS S VSS VPW NCH W=0.47u L=0.06u
MNOE S BCLK M VPW NCH W=0.45u L=0.06u
MNOE017 S NCLK N1_10 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_14 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.62u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.62u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.77u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPOEN S NCLK M VNW PCH W=0.45u L=0.06u
MPOEN019 S BCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_16 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.2u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
.ENDS	SDFFQX3MA10TR

****
.SUBCKT SDFFQX4MA10TR  VDD VSS VPW VNW Q   CK D SE SI
MN0 NMUX D N1 VPW NCH W=0.58u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.58u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.15u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.58u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA108 NS S VSS VPW NCH W=0.7u L=0.06u
MNOE S BCLK M VPW NCH W=0.58u L=0.06u
MNOE017 S NCLK N1_10 VPW NCH W=0.15u L=0.06u
MNOE028 NM BCLK N1_14 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.62u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.62u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1010 NS S VDD VNW PCH W=1.1u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.15u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPOEN S NCLK M VNW PCH W=0.58u L=0.06u
MPOEN019 S BCLK P1_12 VNW PCH W=0.15u L=0.06u
MPOEN030 NM NCLK P1_16 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.2u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
.ENDS	SDFFQX4MA10TR

****
.SUBCKT SDFFRPQNX0P5MA10TR  VDD VSS VPW VNW QN   CK R D SE SI
MN0 NMUX D N1 VPW NCH W=0.27u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.27u L=0.06u
MN2 NET50 NET40 VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.15u L=0.06u
MNA1 NET40 S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA1034 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1038 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1042 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1046 QN S VSS VPW NCH W=0.31u L=0.06u
MNA1050 M NM VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.15u L=0.06u
MNOE NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE022 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NMUX VPW NCH W=0.15u L=0.06u
MNOE030 S BCLK M VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.28u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.28u L=0.06u
MP2 NET39 NET40 NET36 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET39 VNW PCH W=0.2u L=0.06u
MP5 NET36 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NET40 S VDD VNW PCH W=0.15u L=0.06u
MPA1014 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_19 SI VDD VNW PCH W=0.15u L=0.06u
MPA1036 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1040 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1044 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1048 QN S VDD VNW PCH W=0.37u L=0.06u
MPA1053 M NM P1_21 VNW PCH W=0.3u L=0.06u
MPA2 P1_21 R VDD VNW PCH W=0.3u L=0.06u
MPOEN NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN024 NMUX NSE P1_19 VNW PCH W=0.15u L=0.06u
MPOEN028 NM BCLK NMUX VNW PCH W=0.15u L=0.06u
MPOEN032 S NCLK M VNW PCH W=0.15u L=0.06u
.ENDS	SDFFRPQNX0P5MA10TR

****
.SUBCKT SDFFRPQNX1MA10TR  VDD VSS VPW VNW QN   CK R D SE SI
MN0 NMUX D N1 VPW NCH W=0.44u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.44u L=0.06u
MN2 NET53 NET37 VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET53 VPW NCH W=0.15u L=0.06u
MNA1 NET37 S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA1034 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1038 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1042 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1046 QN S VSS VPW NCH W=0.53u L=0.06u
MNA1050 M R VSS VPW NCH W=0.32u L=0.06u
MNA2 M NM VSS VPW NCH W=0.32u L=0.06u
MNOE NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE022 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MNOE030 S BCLK M VPW NCH W=0.28u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.48u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.48u L=0.06u
MP2 NET36 NET37 NET39 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET36 VNW PCH W=0.2u L=0.06u
MP5 NET39 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NET37 S VDD VNW PCH W=0.15u L=0.06u
MPA1014 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1036 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1040 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1044 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1048 QN S VDD VNW PCH W=0.7u L=0.06u
MPA1053 M R P1_21 VNW PCH W=0.64u L=0.06u
MPA2 P1_21 NM VDD VNW PCH W=0.64u L=0.06u
MPOEN NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN024 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN028 NM BCLK NMUX VNW PCH W=0.28u L=0.06u
MPOEN032 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	SDFFRPQNX1MA10TR

****
.SUBCKT SDFFRPQNX2MA10TR  VDD VSS VPW VNW QN   CK R D SE SI
MN0 NMUX D N1 VPW NCH W=0.53u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.53u L=0.06u
MN2 NET53 NET37 VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET53 VPW NCH W=0.15u L=0.06u
MNA1 NET37 S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA1034 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1038 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1042 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1046 QN S VSS VPW NCH W=1.16u L=0.06u
MNA1050 M R VSS VPW NCH W=0.4u L=0.06u
MNA2 M NM VSS VPW NCH W=0.4u L=0.06u
MNOE NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE022 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MNOE030 S BCLK M VPW NCH W=0.4u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.67u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.67u L=0.06u
MP2 NET36 NET37 NET39 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET36 VNW PCH W=0.2u L=0.06u
MP5 NET39 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NET37 S VDD VNW PCH W=0.15u L=0.06u
MPA1014 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1036 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1040 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1044 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1048 QN S VDD VNW PCH W=1.4u L=0.06u
MPA1053 M R P1_21 VNW PCH W=0.8u L=0.06u
MPA2 P1_21 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN024 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN028 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
MPOEN032 S NCLK M VNW PCH W=0.4u L=0.06u
.ENDS	SDFFRPQNX2MA10TR

****
.SUBCKT SDFFRPQNX3MA10TR  VDD VSS VPW VNW QN   CK R D SE SI
MN0 NMUX D N1 VPW NCH W=0.53u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.53u L=0.06u
MN2 NET53 NET37 VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET53 VPW NCH W=0.15u L=0.06u
MNA1 NET37 S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA1034 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1038 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1042 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA1046 QN S VSS VPW NCH W=1.59u L=0.06u
MNA1050 M R VSS VPW NCH W=0.4u L=0.06u
MNA2 M NM VSS VPW NCH W=0.4u L=0.06u
MNOE NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE022 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE030 S BCLK M VPW NCH W=0.51u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.67u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.67u L=0.06u
MP2 NET36 NET37 NET39 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET36 VNW PCH W=0.2u L=0.06u
MP5 NET39 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NET37 S VDD VNW PCH W=0.15u L=0.06u
MPA1014 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1036 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1040 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1044 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA1048 QN S VDD VNW PCH W=2.1u L=0.06u
MPA1053 M R P1_21 VNW PCH W=0.8u L=0.06u
MPA2 P1_21 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN024 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN028 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN032 S NCLK M VNW PCH W=0.59u L=0.06u
.ENDS	SDFFRPQNX3MA10TR

****
.SUBCKT SDFFRPQX0P5MA10TR  VDD VSS VPW VNW Q   CK R D SE SI
MN0 NMUX D N1 VPW NCH W=0.27u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.27u L=0.06u
MN2 NET63 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET63 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1018 M NM VSS VPW NCH W=0.15u L=0.06u
MNA1028 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.3u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNA2 M R VSS VPW NCH W=0.15u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE032 NM BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.28u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.28u L=0.06u
MP2 NET83 NS NET77 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET83 VNW PCH W=0.2u L=0.06u
MP5 NET77 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.2u L=0.06u
MPA1021 M NM P1_13 VNW PCH W=0.3u L=0.06u
MPA1030 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 P1_21 SI VDD VNW PCH W=0.15u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA2 P1_13 R VDD VNW PCH W=0.3u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN034 NM NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_21 VNW PCH W=0.15u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.15u L=0.06u
.ENDS	SDFFRPQX0P5MA10TR

****
.SUBCKT SDFFRPQX1MA10TR  VDD VSS VPW VNW Q   CK R D SE SI
MN0 NMUX D N1 VPW NCH W=0.38u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.38u L=0.06u
MN2 NET139 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET139 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1018 M R VSS VPW NCH W=0.28u L=0.06u
MNA1028 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA109 NS S VSS VPW NCH W=0.3u L=0.06u
MNA2 M NM VSS VPW NCH W=0.28u L=0.06u
MNOE S BCLK M VPW NCH W=0.28u L=0.06u
MNOE032 NM BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.45u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.45u L=0.06u
MP2 NET129 NS NET123 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET129 VNW PCH W=0.2u L=0.06u
MP5 NET123 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1011 NS S VDD VNW PCH W=0.47u L=0.06u
MPA1021 M R P1_13 VNW PCH W=0.7u L=0.06u
MPA1030 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA2 P1_13 NM VDD VNW PCH W=0.7u L=0.06u
MPOEN S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN034 NM NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.28u L=0.06u
.ENDS	SDFFRPQX1MA10TR

****
.SUBCKT SDFFRPQX2MA10TR  VDD VSS VPW VNW Q   CK R D SE SI
MN0 NMUX D N1 VPW NCH W=0.58u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.58u L=0.06u
MN2 NET47 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET47 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1018 M R VSS VPW NCH W=0.4u L=0.06u
MNA1028 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.47u L=0.06u
MNA2 M NM VSS VPW NCH W=0.4u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE032 NM BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.62u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.62u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.69u L=0.06u
MPA1021 M R P1_13 VNW PCH W=0.8u L=0.06u
MPA1030 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA2 P1_13 NM VDD VNW PCH W=0.8u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN034 NM NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
.ENDS	SDFFRPQX2MA10TR

****
.SUBCKT SDFFRPQX3MA10TR  VDD VSS VPW VNW Q   CK R D SE SI
MN0 NMUX D N1 VPW NCH W=0.565u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.565u L=0.06u
MN2 NET140 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET140 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1014 M R VSS VPW NCH W=0.42u L=0.06u
MNA1024 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1032 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1044 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1048 NS S VSS VPW NCH W=0.53u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA2 M NM VSS VPW NCH W=0.42u L=0.06u
MNOE S BCLK M VPW NCH W=0.45u L=0.06u
MNOE028 NM BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE036 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE040 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.635u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.635u L=0.06u
MP2 NET118 NS NET124 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET118 VNW PCH W=0.2u L=0.06u
MP5 NET124 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1017 M R P1_13 VNW PCH W=0.84u L=0.06u
MPA1026 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA1034 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1046 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1050 NS S VDD VNW PCH W=0.68u L=0.06u
MPA1054 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA2 P1_13 NM VDD VNW PCH W=0.84u L=0.06u
MPOEN S NCLK M VNW PCH W=0.45u L=0.06u
MPOEN030 NM NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN038 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN042 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
.ENDS	SDFFRPQX3MA10TR

****
.SUBCKT SDFFRPQX4MA10TR  VDD VSS VPW VNW Q   CK R D SE SI
MN0 NMUX D N1 VPW NCH W=0.54u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.54u L=0.06u
MN2 NET134 NS VSS VPW NCH W=0.15u L=0.06u
MN3 S R VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET134 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1018 M R VSS VPW NCH W=0.42u L=0.06u
MNA1028 N1_15 M VSS VPW NCH W=0.15u L=0.06u
MNA1036 N1_19 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA109 NS S VSS VPW NCH W=0.9u L=0.06u
MNA2 M NM VSS VPW NCH W=0.42u L=0.06u
MNOE S BCLK M VPW NCH W=0.55u L=0.06u
MNOE032 NM BCLK N1_15 VPW NCH W=0.15u L=0.06u
MNOE040 NMUX SE N1_19 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.66u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.66u L=0.06u
MP2 NET124 NS NET118 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET124 VNW PCH W=0.2u L=0.06u
MP5 NET118 R VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1011 NS S VDD VNW PCH W=0.9u L=0.06u
MPA1021 M R P1_13 VNW PCH W=0.84u L=0.06u
MPA1030 P1_17 M VDD VNW PCH W=0.15u L=0.06u
MPA1038 P1_21 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPA2 P1_13 NM VDD VNW PCH W=0.84u L=0.06u
MPOEN S NCLK M VNW PCH W=0.55u L=0.06u
MPOEN034 NM NCLK P1_17 VNW PCH W=0.15u L=0.06u
MPOEN042 NMUX NSE P1_21 VNW PCH W=0.2u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
.ENDS	SDFFRPQX4MA10TR

****
.SUBCKT SDFFSQNX0P5MA10TR  VDD VSS VPW VNW QN   CK D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.3u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.3u L=0.06u
MN2 NET65 NS NET59 VPW NCH W=0.15u L=0.06u
MN3 NET59 SN VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET65 VPW NCH W=0.15u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA1034 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1038 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1042 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1046 QN S VSS VPW NCH W=0.28u L=0.06u
MNA1050 M NM N1_21 VPW NCH W=0.35u L=0.06u
MNA2 N1_21 SN VSS VPW NCH W=0.35u L=0.06u
MNOE NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE022 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NMUX VPW NCH W=0.15u L=0.06u
MNOE030 S BCLK M VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.26u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.26u L=0.06u
MP2 NET45 NS VDD VNW PCH W=0.15u L=0.06u
MP3 S BCLK NET45 VNW PCH W=0.15u L=0.06u
MP4 S SN VDD VNW PCH W=0.15u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_19 SI VDD VNW PCH W=0.15u L=0.06u
MPA1036 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1040 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1044 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA1048 QN S VDD VNW PCH W=0.37u L=0.06u
MPA1053 M NM VDD VNW PCH W=0.22u L=0.06u
MPA2 M SN VDD VNW PCH W=0.22u L=0.06u
MPOEN NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN024 NMUX NSE P1_19 VNW PCH W=0.15u L=0.06u
MPOEN028 NM BCLK NMUX VNW PCH W=0.15u L=0.06u
MPOEN032 S NCLK M VNW PCH W=0.15u L=0.06u
.ENDS	SDFFSQNX0P5MA10TR

****
.SUBCKT SDFFSQNX1MA10TR  VDD VSS VPW VNW QN   CK D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.4u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.4u L=0.06u
MN2 NET50 NS NET53 VPW NCH W=0.2u L=0.06u
MN3 NET53 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.2u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA1034 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1038 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1042 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1046 QN S VSS VPW NCH W=0.53u L=0.06u
MNA1050 M SN N1_21 VPW NCH W=0.58u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.58u L=0.06u
MNOE NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE022 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MNOE030 S BCLK M VPW NCH W=0.28u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.4u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.4u L=0.06u
MP2 NET42 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET42 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1036 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1040 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1044 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1048 QN S VDD VNW PCH W=0.7u L=0.06u
MPA1053 M SN VDD VNW PCH W=0.45u L=0.06u
MPA2 M NM VDD VNW PCH W=0.45u L=0.06u
MPOEN NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN024 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN028 NM BCLK NMUX VNW PCH W=0.28u L=0.06u
MPOEN032 S NCLK M VNW PCH W=0.28u L=0.06u
.ENDS	SDFFSQNX1MA10TR

****
.SUBCKT SDFFSQNX2MA10TR  VDD VSS VPW VNW QN   CK D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.6u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.6u L=0.06u
MN2 NET50 NS NET53 VPW NCH W=0.2u L=0.06u
MN3 NET53 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.2u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1018 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA1034 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1038 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1042 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1046 QN S VSS VPW NCH W=1.06u L=0.06u
MNA1050 M SN N1_21 VPW NCH W=0.6u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.6u L=0.06u
MNOE NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE022 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE026 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MNOE030 S BCLK M VPW NCH W=0.4u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.6u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.6u L=0.06u
MP2 NET42 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET42 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1020 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1036 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1040 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1044 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA1048 QN S VDD VNW PCH W=1.4u L=0.06u
MPA1053 M SN VDD VNW PCH W=0.57u L=0.06u
MPA2 M NM VDD VNW PCH W=0.57u L=0.06u
MPOEN NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN024 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN028 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
MPOEN032 S NCLK M VNW PCH W=0.39u L=0.06u
.ENDS	SDFFSQNX2MA10TR

****
.SUBCKT SDFFSQNX3MA10TR  VDD VSS VPW VNW QN   CK D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.56u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.56u L=0.06u
MN2 NET50 NS NET53 VPW NCH W=0.2u L=0.06u
MN3 NET53 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.2u L=0.06u
MNA1 NS S VSS VPW NCH W=0.15u L=0.06u
MNA1012 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1016 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1022 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA1038 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1042 QN S VSS VPW NCH W=1.59u L=0.06u
MNA1046 M SN N1_21 VPW NCH W=0.6u L=0.06u
MNA1052 BCLK NCLK VSS VPW NCH W=0.24u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.6u L=0.06u
MNOE NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE026 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE030 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE034 S BCLK M VPW NCH W=0.52u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.64u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.64u L=0.06u
MP2 NET42 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET42 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NS S VDD VNW PCH W=0.15u L=0.06u
MPA1014 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1018 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1024 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1040 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1044 QN S VDD VNW PCH W=2.1u L=0.06u
MPA1049 M SN VDD VNW PCH W=0.58u L=0.06u
MPA1054 BCLK NCLK VDD VNW PCH W=0.48u L=0.06u
MPA2 M NM VDD VNW PCH W=0.58u L=0.06u
MPOEN NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN028 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN032 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN036 S NCLK M VNW PCH W=0.52u L=0.06u
.ENDS	SDFFSQNX3MA10TR

****
.SUBCKT SDFFSQX0P5MA10TR  VDD VSS VPW VNW Q   CK D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.3u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.3u L=0.06u
MN2 NET69 NS NET72 VPW NCH W=0.15u L=0.06u
MN3 NET72 SN VSS VPW NCH W=0.15u L=0.06u
MN4 S NCLK NET69 VPW NCH W=0.15u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1022 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1030 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1042 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1046 M NM N1_21 VPW NCH W=0.25u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.31u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNA2 N1_21 SN VSS VPW NCH W=0.25u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE026 NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE034 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE038 NM NCLK NMUX VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.3u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.3u L=0.06u
MP2 NET83 NS VDD VNW PCH W=0.15u L=0.06u
MP3 S BCLK NET83 VNW PCH W=0.15u L=0.06u
MP4 S SN VDD VNW PCH W=0.15u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.3u L=0.06u
MPA1024 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 P1_19 SI VDD VNW PCH W=0.15u L=0.06u
MPA1044 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1049 M NM VDD VNW PCH W=0.22u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.2u L=0.06u
MPA2 M SN VDD VNW PCH W=0.22u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN028 NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN036 NMUX NSE P1_19 VNW PCH W=0.15u L=0.06u
MPOEN040 NM BCLK NMUX VNW PCH W=0.15u L=0.06u
.ENDS	SDFFSQX0P5MA10TR

****
.SUBCKT SDFFSQX1MA10TR  VDD VSS VPW VNW Q   CK D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.4u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.4u L=0.06u
MN2 NET44 NS NET47 VPW NCH W=0.2u L=0.06u
MN3 NET47 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET44 VPW NCH W=0.2u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1022 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1030 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1042 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1046 M SN N1_21 VPW NCH W=0.4u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA108 NS S VSS VPW NCH W=0.3u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.4u L=0.06u
MNOE S BCLK M VPW NCH W=0.28u L=0.06u
MNOE026 NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE034 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE038 NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.4u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.4u L=0.06u
MP2 NET58 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET58 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.5u L=0.06u
MPA1024 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1044 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1049 M SN VDD VNW PCH W=0.4u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA2 M NM VDD VNW PCH W=0.4u L=0.06u
MPOEN S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN028 NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN036 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN040 NM BCLK NMUX VNW PCH W=0.28u L=0.06u
.ENDS	SDFFSQX1MA10TR

****
.SUBCKT SDFFSQX2MA10TR  VDD VSS VPW VNW Q   CK D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.6u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.6u L=0.06u
MN2 NET50 NS NET47 VPW NCH W=0.2u L=0.06u
MN3 NET47 SN VSS VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET50 VPW NCH W=0.2u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1022 N1_13 M VSS VPW NCH W=0.15u L=0.06u
MNA1030 N1_17 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1042 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1046 M SN N1_21 VPW NCH W=0.6u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.46u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.6u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE026 NM BCLK N1_13 VPW NCH W=0.15u L=0.06u
MNOE034 NMUX SE N1_17 VPW NCH W=0.15u L=0.06u
MNOE038 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.6u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.6u L=0.06u
MP2 NET58 NS VDD VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET58 VNW PCH W=0.2u L=0.06u
MP4 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1024 P1_15 M VDD VNW PCH W=0.15u L=0.06u
MPA1032 P1_19 SI VDD VNW PCH W=0.2u L=0.06u
MPA1044 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1049 M SN VDD VNW PCH W=0.57u L=0.06u
MPA1054 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPA2 M NM VDD VNW PCH W=0.57u L=0.06u
MPOEN S NCLK M VNW PCH W=0.39u L=0.06u
MPOEN028 NM NCLK P1_15 VNW PCH W=0.15u L=0.06u
MPOEN036 NMUX NSE P1_19 VNW PCH W=0.2u L=0.06u
MPOEN040 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
.ENDS	SDFFSQX2MA10TR

****
.SUBCKT SDFFSQX3MA10TR  VDD VSS VPW VNW Q   CK D SE SN SI
MN5 NMUX D N1 VPW NCH W=0.58u L=0.06u
MN6 N1 NSE VSS VPW NCH W=0.58u L=0.06u
MN7 S NCLK NET49 VPW NCH W=0.2u L=0.06u
MN8 NET52 SN VSS VPW NCH W=0.2u L=0.06u
MN9 NET49 NS NET52 VPW NCH W=0.2u L=0.06u
MNA1 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1016 N1_13 SI VSS VPW NCH W=0.15u L=0.06u
MNA102 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA1022 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1038 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1042 NS S VSS VPW NCH W=0.47u L=0.06u
MNA1046 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1050 M SN N1_21 VPW NCH W=0.66u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.66u L=0.06u
MNOE NMUX SE N1_13 VPW NCH W=0.15u L=0.06u
MNOE026 NM BCLK N1_17 VPW NCH W=0.15u L=0.06u
MNOE030 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE034 S BCLK M VPW NCH W=0.44u L=0.06u
MP5 P1 SE VDD VNW PCH W=0.62u L=0.06u
MP6 NMUX D P1 VNW PCH W=0.62u L=0.06u
MP7 NET66 NS VDD VNW PCH W=0.2u L=0.06u
MP8 S BCLK NET66 VNW PCH W=0.2u L=0.06u
MP9 S SN VDD VNW PCH W=0.2u L=0.06u
MPA1 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA1018 P1_15 SI VDD VNW PCH W=0.2u L=0.06u
MPA1024 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA104 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1040 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1044 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1048 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1053 M SN VDD VNW PCH W=0.62u L=0.06u
MPA2 M NM VDD VNW PCH W=0.62u L=0.06u
MPOEN NMUX NSE P1_15 VNW PCH W=0.2u L=0.06u
MPOEN028 NM NCLK P1_19 VNW PCH W=0.15u L=0.06u
MPOEN032 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN036 S NCLK M VNW PCH W=0.44u L=0.06u
.ENDS	SDFFSQX3MA10TR

****
.SUBCKT SDFFSQX4MA10TR  VDD VSS VPW VNW Q   CK D SE SN SI
MN10 NET55 SN VSS VPW NCH W=0.2u L=0.06u
MN11 NET52 NS NET55 VPW NCH W=0.2u L=0.06u
MN12 S NCLK NET52 VPW NCH W=0.2u L=0.06u
MN5 NMUX D N1 VPW NCH W=0.55u L=0.06u
MN6 N1 NSE VSS VPW NCH W=0.55u L=0.06u
MNA1 N1_13 SI VSS VPW NCH W=0.15u L=0.06u
MNA1017 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1025 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1029 NS S VSS VPW NCH W=0.8u L=0.06u
MNA1033 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1037 M SN N1_21 VPW NCH W=0.66u L=0.06u
MNA1043 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1047 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA2 N1_21 NM VSS VPW NCH W=0.66u L=0.06u
MNOE NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE013 NMUX SE N1_13 VPW NCH W=0.15u L=0.06u
MNOE021 NM BCLK N1_17 VPW NCH W=0.15u L=0.06u
MNOE06 S BCLK M VPW NCH W=0.53u L=0.06u
MP10 NET66 NS VDD VNW PCH W=0.2u L=0.06u
MP11 S BCLK NET66 VNW PCH W=0.2u L=0.06u
MP12 S SN VDD VNW PCH W=0.2u L=0.06u
MP5 P1 SE VDD VNW PCH W=0.65u L=0.06u
MP6 NMUX D P1 VNW PCH W=0.65u L=0.06u
MPA1 P1_15 SI VDD VNW PCH W=0.2u L=0.06u
MPA1019 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA1027 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1031 NS S VDD VNW PCH W=1u L=0.06u
MPA1035 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1040 M SN VDD VNW PCH W=0.62u L=0.06u
MPA1045 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPA1049 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA2 M NM VDD VNW PCH W=0.62u L=0.06u
MPOEN NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN015 NMUX NSE P1_15 VNW PCH W=0.2u L=0.06u
MPOEN023 NM NCLK P1_19 VNW PCH W=0.15u L=0.06u
MPOEN08 S NCLK M VNW PCH W=0.53u L=0.06u
.ENDS	SDFFSQX4MA10TR

****
.SUBCKT SDFFSRPQX0P5MA10TR  VDD VSS VPW VNW Q   CK R D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.26u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.26u L=0.06u
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.2u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.2u L=0.06u
MN9 M R NET046 VPW NCH W=0.2u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.15u L=0.06u
MNA1031 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1039 N1_21 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1051 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1055 Q NS VSS VPW NCH W=0.31u L=0.06u
MNA108 NS S VSS VPW NCH W=0.15u L=0.06u
MNOE S BCLK M VPW NCH W=0.15u L=0.06u
MNOE035 NM BCLK N1_17 VPW NCH W=0.15u L=0.06u
MNOE043 NMUX SE N1_21 VPW NCH W=0.15u L=0.06u
MNOE047 NM NCLK NMUX VPW NCH W=0.15u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.29u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.29u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.3u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.3u L=0.06u
MP9 M SN VDD VNW PCH W=0.3u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.2u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.22u L=0.06u
MPA1033 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA1041 P1_23 SI VDD VNW PCH W=0.15u L=0.06u
MPA1053 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1057 Q NS VDD VNW PCH W=0.37u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.22u L=0.06u
MPOEN S NCLK M VNW PCH W=0.15u L=0.06u
MPOEN037 NM NCLK P1_19 VNW PCH W=0.15u L=0.06u
MPOEN045 NMUX NSE P1_23 VNW PCH W=0.15u L=0.06u
MPOEN049 NM BCLK NMUX VNW PCH W=0.15u L=0.06u
.ENDS	SDFFSRPQX0P5MA10TR

****
.SUBCKT SDFFSRPQX1MA10TR  VDD VSS VPW VNW Q   CK R D SE SN SI
MN10 NMUX D N1 VPW NCH W=0.4u L=0.06u
MN11 N1 NSE VSS VPW NCH W=0.4u L=0.06u
MN12 M NM NET79 VPW NCH W=0.32u L=0.06u
MN13 NET79 SN VSS VPW NCH W=0.32u L=0.06u
MN14 M R NET79 VPW NCH W=0.32u L=0.06u
MN15 S R NET64 VPW NCH W=0.2u L=0.06u
MN16 NET70 SN VSS VPW NCH W=0.2u L=0.06u
MN17 S NCLK NET61 VPW NCH W=0.2u L=0.06u
MN18 NET64 SN VSS VPW NCH W=0.2u L=0.06u
MN19 NET61 NS NET70 VPW NCH W=0.2u L=0.06u
MNA1 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1021 NCLK CK VSS VPW NCH W=0.17u L=0.06u
MNA1025 BCLK NCLK VSS VPW NCH W=0.15u L=0.06u
MNA1029 Q NS VSS VPW NCH W=0.58u L=0.06u
MNA1033 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1041 N1_21 SI VSS VPW NCH W=0.15u L=0.06u
MNA1049 NS S VSS VPW NCH W=0.28u L=0.06u
MNOE NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MNOE015 S BCLK M VPW NCH W=0.28u L=0.06u
MNOE037 NM BCLK N1_17 VPW NCH W=0.15u L=0.06u
MNOE045 NMUX SE N1_21 VPW NCH W=0.15u L=0.06u
MP10 P1 SE VDD VNW PCH W=0.5u L=0.06u
MP11 NMUX D P1 VNW PCH W=0.5u L=0.06u
MP12 M NM NET108 VNW PCH W=0.6u L=0.06u
MP13 NET108 R VDD VNW PCH W=0.6u L=0.06u
MP14 M SN VDD VNW PCH W=0.6u L=0.06u
MP15 S BCLK NET99 VNW PCH W=0.2u L=0.06u
MP16 NET90 R VDD VNW PCH W=0.2u L=0.06u
MP17 S SN VDD VNW PCH W=0.2u L=0.06u
MP18 NET99 NS NET90 VNW PCH W=0.2u L=0.06u
MPA1 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1023 NCLK CK VDD VNW PCH W=0.22u L=0.06u
MPA1027 BCLK NCLK VDD VNW PCH W=0.3u L=0.06u
MPA1031 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA1035 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA1043 P1_23 SI VDD VNW PCH W=0.2u L=0.06u
MPA1051 NS S VDD VNW PCH W=0.62u L=0.06u
MPOEN NM BCLK NMUX VNW PCH W=0.28u L=0.06u
MPOEN017 S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN039 NM NCLK P1_19 VNW PCH W=0.15u L=0.06u
MPOEN047 NMUX NSE P1_23 VNW PCH W=0.2u L=0.06u
.ENDS	SDFFSRPQX1MA10TR

****
.SUBCKT SDFFSRPQX2MA10TR  VDD VSS VPW VNW Q   CK R D SE SN SI
MN0 NMUX D N1 VPW NCH W=0.54u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.54u L=0.06u
MN2 NET47 NS NET058 VPW NCH W=0.2u L=0.06u
MN3 S R NET064 VPW NCH W=0.2u L=0.06u
MN4 S NCLK NET47 VPW NCH W=0.2u L=0.06u
MN5 NET058 SN VSS VPW NCH W=0.2u L=0.06u
MN6 NET064 SN VSS VPW NCH W=0.2u L=0.06u
MN7 M NM NET046 VPW NCH W=0.35u L=0.06u
MN8 NET046 SN VSS VPW NCH W=0.35u L=0.06u
MN9 M R NET046 VPW NCH W=0.35u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.21u L=0.06u
MNA1031 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1039 N1_21 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.18u L=0.06u
MNA1051 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1055 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.37u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE035 NM BCLK N1_17 VPW NCH W=0.15u L=0.06u
MNOE043 NMUX SE N1_21 VPW NCH W=0.15u L=0.06u
MNOE047 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.66u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.66u L=0.06u
MP2 NET58 NS NET61 VNW PCH W=0.2u L=0.06u
MP3 S BCLK NET58 VNW PCH W=0.2u L=0.06u
MP5 NET61 R VDD VNW PCH W=0.2u L=0.06u
MP6 S SN VDD VNW PCH W=0.2u L=0.06u
MP7 M NM NET081 VNW PCH W=0.7u L=0.06u
MP8 NET081 R VDD VNW PCH W=0.7u L=0.06u
MP9 M SN VDD VNW PCH W=0.7u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.26u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1033 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA1041 P1_23 SI VDD VNW PCH W=0.2u L=0.06u
MPA1053 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1057 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.36u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN037 NM NCLK P1_19 VNW PCH W=0.15u L=0.06u
MPOEN045 NMUX NSE P1_23 VNW PCH W=0.2u L=0.06u
MPOEN049 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
.ENDS	SDFFSRPQX2MA10TR

****
.SUBCKT SDFFSRPQX3MA10TR  VDD VSS VPW VNW Q   CK R D SE SN SI
MN13 NMUX D N1 VPW NCH W=0.545u L=0.06u
MN14 N1 NSE VSS VPW NCH W=0.545u L=0.06u
MN15 S R NET67 VPW NCH W=0.2u L=0.06u
MN16 NET70 SN VSS VPW NCH W=0.2u L=0.06u
MN17 S NCLK NET79 VPW NCH W=0.2u L=0.06u
MN18 NET67 SN VSS VPW NCH W=0.2u L=0.06u
MN19 NET79 NS NET70 VPW NCH W=0.2u L=0.06u
MN20 M NM NET88 VPW NCH W=0.4u L=0.06u
MN21 NET88 SN VSS VPW NCH W=0.4u L=0.06u
MN22 M R NET88 VPW NCH W=0.4u L=0.06u
MNA1 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1023 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1027 NS S VSS VPW NCH W=0.47u L=0.06u
MNA1031 NCLK CK VSS VPW NCH W=0.24u L=0.06u
MNA1035 BCLK NCLK VSS VPW NCH W=0.21u L=0.06u
MNA1039 Q NS VSS VPW NCH W=1.74u L=0.06u
MNA1048 N1_21 SI VSS VPW NCH W=0.15u L=0.06u
MNOE NM BCLK N1_17 VPW NCH W=0.15u L=0.06u
MNOE015 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE019 S BCLK M VPW NCH W=0.45u L=0.06u
MNOE052 NMUX SE N1_21 VPW NCH W=0.15u L=0.06u
MP10 P1 SE VDD VNW PCH W=0.655u L=0.06u
MP11 NMUX D P1 VNW PCH W=0.655u L=0.06u
MP15 S BCLK NET96 VNW PCH W=0.2u L=0.06u
MP16 NET105 R VDD VNW PCH W=0.2u L=0.06u
MP17 S SN VDD VNW PCH W=0.2u L=0.06u
MP18 NET96 NS NET105 VNW PCH W=0.2u L=0.06u
MP19 M NM NET108 VNW PCH W=0.7u L=0.06u
MP20 NET108 R VDD VNW PCH W=0.7u L=0.06u
MP21 M SN VDD VNW PCH W=0.7u L=0.06u
MPA1 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA1025 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1029 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1033 NCLK CK VDD VNW PCH W=0.3u L=0.06u
MPA1037 BCLK NCLK VDD VNW PCH W=0.42u L=0.06u
MPA1041 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA1050 P1_23 SI VDD VNW PCH W=0.2u L=0.06u
MPOEN NM NCLK P1_19 VNW PCH W=0.15u L=0.06u
MPOEN017 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN021 S NCLK M VNW PCH W=0.45u L=0.06u
MPOEN054 NMUX NSE P1_23 VNW PCH W=0.2u L=0.06u
.ENDS	SDFFSRPQX3MA10TR

****
.SUBCKT SDFFSRPQX4MA10TR  VDD VSS VPW VNW Q   CK R D SE SN SI
MN10 NMUX D N1 VPW NCH W=0.53u L=0.06u
MN11 N1 NSE VSS VPW NCH W=0.53u L=0.06u
MN12 S R NET73 VPW NCH W=0.2u L=0.06u
MN13 NET79 SN VSS VPW NCH W=0.2u L=0.06u
MN14 S NCLK NET70 VPW NCH W=0.2u L=0.06u
MN15 NET73 SN VSS VPW NCH W=0.2u L=0.06u
MN16 NET70 NS NET79 VPW NCH W=0.2u L=0.06u
MN17 M NM NET64 VPW NCH W=0.4u L=0.06u
MN18 NET64 SN VSS VPW NCH W=0.4u L=0.06u
MN19 M R NET64 VPW NCH W=0.4u L=0.06u
MNA1 N1_17 M VSS VPW NCH W=0.15u L=0.06u
MNA1025 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1029 NS S VSS VPW NCH W=0.8u L=0.06u
MNA1033 NCLK CK VSS VPW NCH W=0.28u L=0.06u
MNA1037 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1041 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA1045 N1_21 SI VSS VPW NCH W=0.15u L=0.06u
MNOE NM BCLK N1_17 VPW NCH W=0.15u L=0.06u
MNOE017 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE021 S BCLK M VPW NCH W=0.44u L=0.06u
MNOE049 NMUX SE N1_21 VPW NCH W=0.15u L=0.06u
MP10 P1 SE VDD VNW PCH W=0.67u L=0.06u
MP11 NMUX D P1 VNW PCH W=0.67u L=0.06u
MP12 S BCLK NET108 VNW PCH W=0.2u L=0.06u
MP13 NET99 R VDD VNW PCH W=0.2u L=0.06u
MP14 S SN VDD VNW PCH W=0.2u L=0.06u
MP15 NET108 NS NET99 VNW PCH W=0.2u L=0.06u
MP16 M NM NET96 VNW PCH W=0.7u L=0.06u
MP17 NET96 R VDD VNW PCH W=0.7u L=0.06u
MP18 M SN VDD VNW PCH W=0.7u L=0.06u
MPA1 P1_19 M VDD VNW PCH W=0.15u L=0.06u
MPA1027 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1031 NS S VDD VNW PCH W=1u L=0.06u
MPA1035 NCLK CK VDD VNW PCH W=0.35u L=0.06u
MPA1039 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPA1043 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA1047 P1_23 SI VDD VNW PCH W=0.2u L=0.06u
MPOEN NM NCLK P1_19 VNW PCH W=0.15u L=0.06u
MPOEN019 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN023 S NCLK M VNW PCH W=0.58u L=0.06u
MPOEN051 NMUX NSE P1_23 VNW PCH W=0.2u L=0.06u
.ENDS	SDFFSRPQX4MA10TR

****
.SUBCKT SDFFYQX1MA10TR  VDD VSS VPW VNW Q   CK D SE SI
MN0 NMUX D N1 VPW NCH W=0.4u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.4u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.29u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.4u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.4u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.32u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.25u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=0.53u L=0.06u
MNA108 NS S VSS VPW NCH W=0.32u L=0.06u
MNOE S BCLK M VPW NCH W=0.28u L=0.06u
MNOE017 S NCLK N1_10 VPW NCH W=0.4u L=0.06u
MNOE028 NM BCLK N1_14 VPW NCH W=0.4u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.28u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.56u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.56u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.36u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.5u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.4u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.4u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.5u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=0.7u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.5u L=0.06u
MPOEN S NCLK M VNW PCH W=0.28u L=0.06u
MPOEN019 S BCLK P1_12 VNW PCH W=0.4u L=0.06u
MPOEN030 NM NCLK P1_16 VNW PCH W=0.4u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.2u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.28u L=0.06u
.ENDS	SDFFYQX1MA10TR

****
.SUBCKT SDFFYQX2MA10TR  VDD VSS VPW VNW Q   CK D SE SI
MN0 NMUX D N1 VPW NCH W=0.515u L=0.06u
MN1 N1 NSE VSS VPW NCH W=0.515u L=0.06u
MNA1 NCLK CK VSS VPW NCH W=0.42u L=0.06u
MNA1013 N1_10 NS VSS VPW NCH W=0.4u L=0.06u
MNA1024 N1_14 M VSS VPW NCH W=0.4u L=0.06u
MNA1032 M NM VSS VPW NCH W=0.4u L=0.06u
MNA1036 N1_18 SI VSS VPW NCH W=0.15u L=0.06u
MNA104 BCLK NCLK VSS VPW NCH W=0.34u L=0.06u
MNA1048 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.16u L=0.06u
MNA108 NS S VSS VPW NCH W=0.53u L=0.06u
MNOE S BCLK M VPW NCH W=0.4u L=0.06u
MNOE017 S NCLK N1_10 VPW NCH W=0.4u L=0.06u
MNOE028 NM BCLK N1_14 VPW NCH W=0.4u L=0.06u
MNOE040 NMUX SE N1_18 VPW NCH W=0.15u L=0.06u
MNOE044 NM NCLK NMUX VPW NCH W=0.4u L=0.06u
MP0 NMUX D P1 VNW PCH W=0.685u L=0.06u
MP1 P1 SE VDD VNW PCH W=0.685u L=0.06u
MPA1 NCLK CK VDD VNW PCH W=0.52u L=0.06u
MPA1010 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1015 P1_12 NS VDD VNW PCH W=0.4u L=0.06u
MPA1026 P1_16 M VDD VNW PCH W=0.4u L=0.06u
MPA1034 M NM VDD VNW PCH W=0.6u L=0.06u
MPA1038 P1_20 SI VDD VNW PCH W=0.2u L=0.06u
MPA1050 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1054 Q NS VDD VNW PCH W=1.4u L=0.06u
MPA106 BCLK NCLK VDD VNW PCH W=0.68u L=0.06u
MPOEN S NCLK M VNW PCH W=0.4u L=0.06u
MPOEN019 S BCLK P1_12 VNW PCH W=0.4u L=0.06u
MPOEN030 NM NCLK P1_16 VNW PCH W=0.4u L=0.06u
MPOEN042 NMUX NSE P1_20 VNW PCH W=0.2u L=0.06u
MPOEN046 NM BCLK NMUX VNW PCH W=0.4u L=0.06u
.ENDS	SDFFYQX2MA10TR

****
.SUBCKT SDFFYQX3MA10TR  VDD VSS VPW VNW Q   CK D SE SI
MN4 NMUX D N1 VPW NCH W=0.5u L=0.06u
MN5 N1 NSE VSS VPW NCH W=0.5u L=0.06u
MNA1 N1_10 SI VSS VPW NCH W=0.15u L=0.06u
MNA1016 N1_18 M VSS VPW NCH W=0.4u L=0.06u
MNA1032 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1036 NS S VSS VPW NCH W=0.4u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.3u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.26u L=0.06u
MNA1048 M NM VSS VPW NCH W=0.38u L=0.06u
MNA105 N1_14 NS VSS VPW NCH W=0.4u L=0.06u
MNA1052 Q NS VSS VPW NCH W=1.74u L=0.06u
MNOE NMUX SE N1_10 VPW NCH W=0.15u L=0.06u
MNOE020 NM BCLK N1_18 VPW NCH W=0.4u L=0.06u
MNOE024 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.45u L=0.06u
MNOE09 S NCLK N1_14 VPW NCH W=0.4u L=0.06u
MP4 P1 SE VDD VNW PCH W=0.7u L=0.06u
MP5 NMUX D P1 VNW PCH W=0.7u L=0.06u
MPA1 P1_12 SI VDD VNW PCH W=0.2u L=0.06u
MPA1018 P1_20 M VDD VNW PCH W=0.4u L=0.06u
MPA1034 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1038 NS S VDD VNW PCH W=0.7u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.37u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.52u L=0.06u
MPA1050 M NM VDD VNW PCH W=0.76u L=0.06u
MPA1054 Q NS VDD VNW PCH W=2.1u L=0.06u
MPA107 P1_16 NS VDD VNW PCH W=0.4u L=0.06u
MPOEN NMUX NSE P1_12 VNW PCH W=0.2u L=0.06u
MPOEN011 S BCLK P1_16 VNW PCH W=0.4u L=0.06u
MPOEN022 NM NCLK P1_20 VNW PCH W=0.4u L=0.06u
MPOEN026 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.45u L=0.06u
.ENDS	SDFFYQX3MA10TR

****
.SUBCKT SDFFYQX4MA10TR  VDD VSS VPW VNW Q   CK D SE SI
MN2 NMUX D N1 VPW NCH W=0.5u L=0.06u
MN3 N1 NSE VSS VPW NCH W=0.5u L=0.06u
MNA1 N1_10 SI VSS VPW NCH W=0.15u L=0.06u
MNA1016 N1_18 M VSS VPW NCH W=0.4u L=0.06u
MNA1032 NSE SE VSS VPW NCH W=0.15u L=0.06u
MNA1036 NS S VSS VPW NCH W=1.05u L=0.06u
MNA1040 NCLK CK VSS VPW NCH W=0.38u L=0.06u
MNA1044 BCLK NCLK VSS VPW NCH W=0.35u L=0.06u
MNA1048 M NM VSS VPW NCH W=0.45u L=0.06u
MNA1052 Q NS VSS VPW NCH W=2.32u L=0.06u
MNA107 N1_14 NS VSS VPW NCH W=0.4u L=0.06u
MNOE NMUX SE N1_10 VPW NCH W=0.15u L=0.06u
MNOE011 S NCLK N1_14 VPW NCH W=0.4u L=0.06u
MNOE020 NM BCLK N1_18 VPW NCH W=0.4u L=0.06u
MNOE024 NM NCLK NMUX VPW NCH W=0.45u L=0.06u
MNOE028 S BCLK M VPW NCH W=0.57u L=0.06u
MP2 P1 SE VDD VNW PCH W=0.7u L=0.06u
MP3 NMUX D P1 VNW PCH W=0.7u L=0.06u
MPA1 P1_12 SI VDD VNW PCH W=0.2u L=0.06u
MPA1018 P1_20 M VDD VNW PCH W=0.4u L=0.06u
MPA1034 NSE SE VDD VNW PCH W=0.2u L=0.06u
MPA1038 NS S VDD VNW PCH W=1.25u L=0.06u
MPA1042 NCLK CK VDD VNW PCH W=0.47u L=0.06u
MPA1046 BCLK NCLK VDD VNW PCH W=0.7u L=0.06u
MPA1050 M NM VDD VNW PCH W=0.7u L=0.06u
MPA1054 Q NS VDD VNW PCH W=2.8u L=0.06u
MPA109 P1_16 NS VDD VNW PCH W=0.4u L=0.06u
MPOEN NMUX NSE P1_12 VNW PCH W=0.2u L=0.06u
MPOEN013 S BCLK P1_16 VNW PCH W=0.4u L=0.06u
MPOEN022 NM NCLK P1_20 VNW PCH W=0.4u L=0.06u
MPOEN026 NM BCLK NMUX VNW PCH W=0.45u L=0.06u
MPOEN030 S NCLK M VNW PCH W=0.57u L=0.06u
.ENDS	SDFFYQX4MA10TR

****

****

****
.SUBCKT XNOR2X0P5MA10TR  VDD VSS VPW VNW Y   A B
MNA1 NIN2 B VSS VPW NCH W=0.235u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.235u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.275u L=0.06u
MNOE Y NIN1 NIN2 VPW NCH W=0.235u L=0.06u
MNOE02 Y A BIN2 VPW NCH W=0.235u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.35u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.37u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.35u L=0.06u
MPOEN Y A NIN2 VNW PCH W=0.235u L=0.06u
MPOEN04 Y NIN1 BIN2 VNW PCH W=0.235u L=0.06u
.ENDS	XNOR2X0P5MA10TR

****
.SUBCKT XNOR2X0P7MA10TR  VDD VSS VPW VNW Y   A B
MNA1 NIN2 B VSS VPW NCH W=0.33u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.33u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.31u L=0.06u
MNOE Y NIN1 NIN2 VPW NCH W=0.33u L=0.06u
MNOE02 Y A BIN2 VPW NCH W=0.33u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.49u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.42u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.49u L=0.06u
MPOEN Y A NIN2 VNW PCH W=0.33u L=0.06u
MPOEN04 Y NIN1 BIN2 VNW PCH W=0.33u L=0.06u
.ENDS	XNOR2X0P7MA10TR

****
.SUBCKT XNOR2X1MA10TR  VDD VSS VPW VNW Y   A B
MNA1 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.38u L=0.06u
MNOE Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MNOE02 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.49u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MPOEN Y A NIN2 VNW PCH W=0.47u L=0.06u
MPOEN04 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
.ENDS	XNOR2X1MA10TR

****

****

****

****

****
.SUBCKT XNOR3X0P5MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 NIN3 C VSS VPW NCH W=0.26u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.2u L=0.06u
MNA1020 NIN2 B VSS VPW NCH W=0.26u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.2u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.26u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=0.265u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.26u L=0.06u
MNOE012 NOUT A XNOR23 VPW NCH W=0.2u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.26u L=0.06u
MNOE08 NOUT NIN1 XOR23 VPW NCH W=0.2u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=0.39u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.3u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.35u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.27u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=0.39u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=0.35u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.32u L=0.06u
MPOEN010 NOUT A XOR23 VNW PCH W=0.24u L=0.06u
MPOEN014 NOUT NIN1 XNOR23 VNW PCH W=0.24u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.32u L=0.06u
.ENDS	XNOR3X0P5MA10TR

****

****

****

****

****
.SUBCKT XNOR3X3MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 NIN3 C VSS VPW NCH W=1.335u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.89u L=0.06u
MNA1020 NIN2 B VSS VPW NCH W=0.98u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.66u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=1.335u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=1.59u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=1.335u L=0.06u
MNOE012 NOUT A XNOR23 VPW NCH W=0.89u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=1.335u L=0.06u
MNOE08 NOUT NIN1 XOR23 VPW NCH W=0.89u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=2.01u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=1.33u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=1.3u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.88u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=2.01u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=2.1u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=1.335u L=0.06u
MPOEN010 NOUT A XOR23 VNW PCH W=1.09u L=0.06u
MPOEN014 NOUT NIN1 XNOR23 VNW PCH W=1.09u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=1.335u L=0.06u
.ENDS	XNOR3X3MA10TR

****
.SUBCKT XNOR3X4MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 NIN3 C VSS VPW NCH W=1.68u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=1.13u L=0.06u
MNA1020 NIN2 B VSS VPW NCH W=1.23u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.82u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=1.68u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=2.12u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=1.68u L=0.06u
MNOE012 NOUT A XNOR23 VPW NCH W=1.13u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=1.68u L=0.06u
MNOE08 NOUT NIN1 XOR23 VPW NCH W=1.13u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=2.52u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=1.695u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=1.65u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=1.1u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=2.52u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=2.8u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=1.68u L=0.06u
MPOEN010 NOUT A XOR23 VNW PCH W=1.41u L=0.06u
MPOEN014 NOUT NIN1 XNOR23 VNW PCH W=1.41u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=1.68u L=0.06u
.ENDS	XNOR3X4MA10TR

****
.SUBCKT XOR2X0P5MA10TR  VDD VSS VPW VNW Y   A B
MNA1 NIN2 B VSS VPW NCH W=0.235u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.235u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.275u L=0.06u
MNOE Y A NIN2 VPW NCH W=0.235u L=0.06u
MNOE02 Y NIN1 BIN2 VPW NCH W=0.235u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.35u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.37u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.35u L=0.06u
MPOEN Y NIN1 NIN2 VNW PCH W=0.235u L=0.06u
MPOEN04 Y A BIN2 VNW PCH W=0.235u L=0.06u
.ENDS	XOR2X0P5MA10TR

****
.SUBCKT XOR2X0P7MA10TR  VDD VSS VPW VNW Y   A B
MNA1 NIN2 B VSS VPW NCH W=0.33u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.33u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.31u L=0.06u
MNOE Y A NIN2 VPW NCH W=0.33u L=0.06u
MNOE02 Y NIN1 BIN2 VPW NCH W=0.33u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.49u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.42u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.49u L=0.06u
MPOEN Y NIN1 NIN2 VNW PCH W=0.33u L=0.06u
MPOEN04 Y A BIN2 VNW PCH W=0.33u L=0.06u
.ENDS	XOR2X0P7MA10TR

****
.SUBCKT XOR2X1MA10TR  VDD VSS VPW VNW Y   A B
MNA1 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.38u L=0.06u
MNOE Y A NIN2 VPW NCH W=0.47u L=0.06u
MNOE02 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.49u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MPOEN Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MPOEN04 Y A BIN2 VNW PCH W=0.47u L=0.06u
.ENDS	XOR2X1MA10TR

****

****

****

****

****
.SUBCKT XOR3X0P5MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 NIN3 C VSS VPW NCH W=0.26u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.2u L=0.06u
MNA1020 NIN2 B VSS VPW NCH W=0.265u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.2u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.26u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=0.265u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.26u L=0.06u
MNOE012 NOUT NIN1 XNOR23 VPW NCH W=0.2u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.26u L=0.06u
MNOE08 NOUT A XOR23 VPW NCH W=0.2u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=0.39u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.3u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.35u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.27u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=0.39u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=0.35u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.32u L=0.06u
MPOEN010 NOUT NIN1 XOR23 VNW PCH W=0.24u L=0.06u
MPOEN014 NOUT A XNOR23 VNW PCH W=0.24u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.32u L=0.06u
.ENDS	XOR3X0P5MA10TR

****

****

****

****
.SUBCKT XOR3X2MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 NIN3 C VSS VPW NCH W=0.89u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.63u L=0.06u
MNA1020 NIN2 B VSS VPW NCH W=0.72u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.47u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.89u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=1.06u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.89u L=0.06u
MNOE012 NOUT NIN1 XNOR23 VPW NCH W=0.63u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.89u L=0.06u
MNOE08 NOUT A XOR23 VPW NCH W=0.63u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=1.33u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.94u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.96u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.63u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=1.33u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=1.4u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.89u L=0.06u
MPOEN010 NOUT NIN1 XOR23 VNW PCH W=0.77u L=0.06u
MPOEN014 NOUT A XNOR23 VNW PCH W=0.77u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.89u L=0.06u
.ENDS	XOR3X2MA10TR

****
.SUBCKT XOR3X3MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 NIN3 C VSS VPW NCH W=1.335u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.89u L=0.06u
MNA1020 NIN2 B VSS VPW NCH W=0.98u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.66u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=1.335u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=1.59u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=1.335u L=0.06u
MNOE012 NOUT NIN1 XNOR23 VPW NCH W=0.89u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=1.335u L=0.06u
MNOE08 NOUT A XOR23 VPW NCH W=0.89u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=2.01u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=1.33u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=1.3u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.88u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=2.01u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=2.1u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=1.335u L=0.06u
MPOEN010 NOUT NIN1 XOR23 VNW PCH W=1.09u L=0.06u
MPOEN014 NOUT A XNOR23 VNW PCH W=1.09u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=1.335u L=0.06u
.ENDS	XOR3X3MA10TR

****
.SUBCKT XOR3X4MA10TR  VDD VSS VPW VNW Y   A B C
MNA1 NIN3 C VSS VPW NCH W=1.68u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=1.13u L=0.06u
MNA1020 NIN2 B VSS VPW NCH W=1.23u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.82u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=1.68u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=2.12u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=1.68u L=0.06u
MNOE012 NOUT NIN1 XNOR23 VPW NCH W=1.13u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=1.68u L=0.06u
MNOE08 NOUT A XOR23 VPW NCH W=1.13u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=2.52u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=1.695u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=1.65u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=1.1u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=2.52u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=2.8u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=1.68u L=0.06u
MPOEN010 NOUT NIN1 XOR23 VNW PCH W=1.41u L=0.06u
MPOEN014 NOUT A XNOR23 VNW PCH W=1.41u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=1.68u L=0.06u
.ENDS	XOR3X4MA10TR
****
.SUBCKT	FILL128A10TR	VDD	VSS	VPW	VNW
.ENDS FILL128A10TR

****
.SUBCKT	FILL16A10TR	VDD	VSS	VPW	VNW
.ENDS FILL16A10TR

****
.SUBCKT	FILL18CAP128A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_18 W=22.8u L=0.705u
.ENDS FILL18CAP128A10TR

****
.SUBCKT	FILL18CAP12A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_18 W=0.95u L=0.85u
.ENDS FILL18CAP12A10TR

****
.SUBCKT	FILL18CAP16A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_18 W=1.9u L=0.67u
.ENDS FILL18CAP16A10TR

****
.SUBCKT	FILL18CAP32A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_18 W=4.75u L=0.72u
.ENDS FILL18CAP32A10TR

****
.SUBCKT	FILL18CAP64A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_18 W=10.45u L=0.74u
.ENDS FILL18CAP64A10TR

****
.SUBCKT	FILL18CAPTIE128A10TR	VDD	VSS
MN0 VSS VDD VSS VSS NCH_18 W=21.85u L=0.73u
.ENDS FILL18CAPTIE128A10TR

****
.SUBCKT	FILL18CAPTIE12A10TR	VDD	VSS
MN0 VSS VDD VSS VSS NCH_18 W=0.95u L=0.47u
.ENDS FILL18CAPTIE12A10TR

****
.SUBCKT	FILL18CAPTIE16A10TR	VDD	VSS
MN0 VSS VDD VSS VSS NCH_18 W=0.95u L=1.27u
.ENDS FILL18CAPTIE16A10TR

****
.SUBCKT	FILL18CAPTIE32A10TR	VDD     VSS
MN0 VSS VDD VSS VSS NCH_18 W=3.8u L=0.885u
.ENDS FILL18CAPTIE32A10TR

****
.SUBCKT	FILL18CAPTIE64A10TR	VDD	VSS
MN0 VSS VDD VSS VSS NCH_18 W=10.45u L=0.705u
.ENDS FILL18CAPTIE64A10TR

****
.SUBCKT	FILL1A10TR	VDD	VSS	VPW	VNW
.ENDS FILL1A10TR

****
.SUBCKT	FILL25CAP128A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_25 W=22.8u L=0.705u
.ENDS FILL25CAP128A10TR

****
.SUBCKT	FILL25CAP12A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_25 W=0.95u L=0.85u
.ENDS FILL25CAP12A10TR

****
.SUBCKT	FILL25CAP16A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_25 W=1.9u L=0.67u
.ENDS FILL25CAP16A10TR

****
.SUBCKT	FILL25CAP32A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_25 W=4.75u L=0.72u
.ENDS FILL25CAP32A10TR

****
.SUBCKT	FILL25CAP64A10TR	VDD	VSS	VPW	VNW
MN0 VSS VDD VSS VPW NCH_25 W=10.45u L=0.74u
.ENDS FILL25CAP64A10TR

****
.SUBCKT	FILL25CAPTIE128A10TR	VDD	VSS
MN0 VSS VDD VSS VSS NCH_25 W=21.85u L=0.73u
.ENDS FILL25CAPTIE128A10TR

****
.SUBCKT	FILL25CAPTIE12A10TR	VDD	VSS
MN0 VSS VDD VSS VSS NCH_25 W=0.95u L=0.47u
.ENDS FILL25CAPTIE12A10TR

****
.SUBCKT	FILL25CAPTIE16A10TR	VDD	VSS
MN0 VSS VDD VSS VSS NCH_25 W=0.95u L=1.27u
.ENDS FILL25CAPTIE16A10TR

****
.SUBCKT	FILL25CAPTIE32A10TR	VDD	VSS
MN0 VSS VDD VSS VSS NCH_25 W=3.8u L=0.885u
.ENDS FILL25CAPTIE32A10TR

****
.SUBCKT	FILL25CAPTIE64A10TR	VDD	VSS
MN0 VSS VDD VSS VSS NCH_25 W=10.45u L=0.705u
.ENDS FILL25CAPTIE64A10TR

****
.SUBCKT	FILL2A10TR	VDD	VSS	VPW	VNW
.ENDS FILL2A10TR

****
.SUBCKT	FILL32A10TR	VDD	VSS	VPW	VNW
.ENDS FILL32A10TR

****
.SUBCKT	FILL4A10TR	VDD	VSS	VPW	VNW
.ENDS FILL4A10TR

****
.SUBCKT	FILL64A10TR	VDD	VSS	VPW	VNW
.ENDS FILL64A10TR

****
.SUBCKT	FILL8A10TR	VDD	VSS	VPW	VNW
.ENDS FILL8A10TR

****
.SUBCKT	FILLCAP128A10TR	VDD	VSS	VPW	VNW
MN1 NET10 NET9 VSS VPW NCH W=45.59u L=0.06u
MP0 NET9 NET10 VDD VNW PCH W=67.9u L=0.06u
.ENDS FILLCAP128A10TR

****
.SUBCKT	FILLCAP16A10TR	VDD	VSS	VPW	VNW
MN1 NET10 NET9 VSS VPW NCH W=5.17u L=0.06u
MP0 NET9 NET10 VDD VNW PCH W=7.7u L=0.06u
.ENDS FILLCAP16A10TR

****
.SUBCKT	FILLCAP32A10TR	VDD	VSS	VPW	VNW
MN1 NET10 NET9 VSS VPW NCH W=10.81u L=0.06u
MP0 NET9 NET10 VDD VNW PCH W=16.1u L=0.06u
.ENDS FILLCAP32A10TR

****
.SUBCKT	FILLCAP3A10TR	VDD	VSS	VPW	VNW
MN1 NET10 NET9 VSS VPW NCH W=0.47u L=0.06u
MP0 NET9 NET10 VDD VNW PCH W=0.7u L=0.06u
.ENDS FILLCAP3A10TR

****
.SUBCKT	FILLCAP4A10TR	VDD	VSS	VPW	VNW
MN1 NET10 NET9 VSS VPW NCH W=0.94u L=0.06u
MP0 NET9 NET10 VDD VNW PCH W=1.4u L=0.06u
.ENDS FILLCAP4A10TR

****
.SUBCKT	FILLCAP64A10TR	VDD	VSS	VPW	VNW
MN1 NET10 NET9 VSS VPW NCH W=22.56u L=0.06u
MP0 NET9 NET10 VDD VNW PCH W=33.6u L=0.06u
.ENDS FILLCAP64A10TR

****
.SUBCKT	FILLCAP8A10TR	VDD	VSS	VPW	VNW
MN1 NET10 NET9 VSS VPW NCH W=2.35u L=0.06u
MP0 NET9 NET10 VDD VNW PCH W=3.5u L=0.06u
.ENDS FILLCAP8A10TR

****
.SUBCKT	FILLCAPTIE128A10TR	VDD	VSS
MN1 NET10 NET9 VSS VSS NCH W=44.18u L=0.06u
MP0 NET9 NET10 VDD VDD PCH W=65.8u L=0.06u
.ENDS FILLCAPTIE128A10TR

****
.SUBCKT	FILLCAPTIE16A10TR	VDD	VSS
MN1 NET10 NET9 VSS VSS NCH W=3.76u L=0.06u
MP0 NET9 NET10 VDD VDD PCH W=5.6u L=0.06u
.ENDS FILLCAPTIE16A10TR

****
.SUBCKT	FILLCAPTIE32A10TR	VDD	VSS
MN1 NET10 NET9 VSS VSS NCH W=9.4u L=0.06u
MP0 NET9 NET10 VDD VDD PCH W=14u L=0.06u
.ENDS FILLCAPTIE32A10TR

****
.SUBCKT	FILLCAPTIE64A10TR	VDD	VSS
MN1 NET10 NET9 VSS VSS NCH W=21.15u L=0.06u
MP0 NET9 NET10 VDD VDD PCH W=31.5u L=0.06u
.ENDS FILLCAPTIE64A10TR

****
.SUBCKT	FILLCAPTIE6A10TR	VDD	VSS
MN1 NET10 NET9 VSS VSS NCH W=0.94u L=0.06u
MP0 NET9 NET10 VDD VDD PCH W=1.4u L=0.06u
.ENDS FILLCAPTIE6A10TR

****
.SUBCKT	FILLCAPTIE8A10TR	VDD	VSS
MN1 NET10 NET9 VSS VSS NCH W=0.94u L=0.06u
MP0 NET9 NET10 VDD VDD PCH W=1.4u L=0.06u
.ENDS FILLCAPTIE8A10TR

****
.SUBCKT	FILLTIE128A10TR	VDD	VSS
.ENDS FILLTIE128A10TR

****
.SUBCKT	FILLTIE16A10TR	VDD	VSS
.ENDS FILLTIE16A10TR

****
.SUBCKT	FILLTIE2A10TR	VDD	VSS
.ENDS FILLTIE2A10TR

****
.SUBCKT	FILLTIE32A10TR	VDD	VSS
.ENDS FILLTIE32A10TR

****
.SUBCKT	FILLTIE4A10TR	VDD	VSS
.ENDS FILLTIE4A10TR

****
.SUBCKT	FILLTIE64A10TR	VDD	VSS
.ENDS FILLTIE64A10TR

****
.SUBCKT	FILLTIE8A10TR	VDD	VSS
.ENDS FILLTIE8A10TR


****
.SUBCKT AND2X11MA10TR VDD VSS VPW VNW Y A B
MPA2_6 INT B VDD VNW PCH W=0.435u L=0.06u
MNA2_3 VSS B N_53 VPW NCH W=0.53u L=0.06u
MPA1_3 INT A VDD VNW PCH W=0.435u L=0.06u
MNA1_3 INT A N_53 VPW NCH W=0.53u L=0.06u
MNA1 INT A N_55 VPW NCH W=0.53u L=0.06u
MPA1_2 INT A VDD VNW PCH W=0.435u L=0.06u
MPA2_5 INT B VDD VNW PCH W=0.435u L=0.06u
MNA2 VSS B N_55 VPW NCH W=0.53u L=0.06u
MNA2_6 VSS B N_57 VPW NCH W=0.53u L=0.06u
MPA2_4 INT B VDD VNW PCH W=0.435u L=0.06u
MNA1_6 INT A N_57 VPW NCH W=0.53u L=0.06u
MPA1 INT A VDD VNW PCH W=0.435u L=0.06u
MNA1_4 INT A N_59 VPW NCH W=0.53u L=0.06u
MPA1_6 INT A VDD VNW PCH W=0.435u L=0.06u
MPA2_3 INT B VDD VNW PCH W=0.435u L=0.06u
MNA2_4 VSS B N_59 VPW NCH W=0.53u L=0.06u
MNA2_2 VSS B N_61 VPW NCH W=0.535u L=0.06u
MPA2_2 INT B VDD VNW PCH W=0.435u L=0.06u
MNA1_2 INT A N_61 VPW NCH W=0.535u L=0.06u
MPA1_5 INT A VDD VNW PCH W=0.435u L=0.06u
MNA1_5 INT A N_64 VPW NCH W=0.535u L=0.06u
MPA1_4 INT A VDD VNW PCH W=0.44u L=0.06u
MNA2_5 N_64 B VSS VPW NCH W=0.535u L=0.06u
MPA2 INT B VDD VNW PCH W=0.44u L=0.06u
MNA104_7 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_5 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_10 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_8 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_10 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_6 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_8 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_6 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_11 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_9 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_11 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_7 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_9 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_5 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AND2X11MA10TR

****
.SUBCKT AND2X3MA10TR VDD VSS VPW VNW Y A B
MPA2 INT B VDD VNW PCH W=0.36u L=0.06u
MNA2 VSS B N_17 VPW NCH W=0.44u L=0.06u
MPA1 INT A VDD VNW PCH W=0.36u L=0.06u
MNA1 INT A N_17 VPW NCH W=0.44u L=0.06u
MNA1_2 INT A N_19 VPW NCH W=0.44u L=0.06u
MPA1_2 INT A VDD VNW PCH W=0.36u L=0.06u
MNA2_2 N_19 B VSS VPW NCH W=0.44u L=0.06u
MPA2_2 INT B VDD VNW PCH W=0.36u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AND2X3MA10TR

****
.SUBCKT NAND2X3MA10TR VDD VSS VPW VNW Y A B
MPA2_3 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS B N_19 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1 Y A N_19 VPW NCH W=0.58u L=0.06u
MNA1_3 Y A N_21 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_3 VSS B N_21 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_2 VSS B N_17 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_2 N_17 A Y VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2X3MA10TR

****
.SUBCKT AND2X4MA10TR VDD VSS VPW VNW Y A B
MPA2_2 INT B VDD VNW PCH W=0.47u L=0.06u
MNA2 VSS B N_24 VPW NCH W=0.58u L=0.06u
MPA1_2 INT A VDD VNW PCH W=0.47u L=0.06u
MNA1 N_24 A INT VPW NCH W=0.58u L=0.06u
MNA1_2 INT A N_26 VPW NCH W=0.575u L=0.06u
MPA1 INT A VDD VNW PCH W=0.475u L=0.06u
MNA2_2 N_26 B VSS VPW NCH W=0.575u L=0.06u
MPA2 INT B VDD VNW PCH W=0.475u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_4 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AND2X4MA10TR

****
.SUBCKT NAND2X4MA10TR VDD VSS VPW VNW Y A B
MPA2_4 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS B N_23 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1 Y A N_23 VPW NCH W=0.58u L=0.06u
MNA1_3 Y A N_25 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_3 VSS B N_25 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_2 VSS B N_27 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y A N_27 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_4 Y A N_21 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_4 N_21 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2X4MA10TR

****
.SUBCKT AND2X6MA10TR VDD VSS VPW VNW Y A B
MPA1_2 INT A VDD VNW PCH W=0.475u L=0.06u
MNA1_3 INT A N_32 VPW NCH W=0.58u L=0.06u
MPA2_3 INT B VDD VNW PCH W=0.475u L=0.06u
MNA2_3 N_32 B VSS VPW NCH W=0.58u L=0.06u
MNA2 VSS B N_33 VPW NCH W=0.575u L=0.06u
MPA2 INT B VDD VNW PCH W=0.475u L=0.06u
MNA1 INT A N_33 VPW NCH W=0.575u L=0.06u
MPA1_3 INT A VDD VNW PCH W=0.475u L=0.06u
MNA1_2 INT A N_36 VPW NCH W=0.575u L=0.06u
MPA1 INT A VDD VNW PCH W=0.47u L=0.06u
MNA2_2 N_36 B VSS VPW NCH W=0.575u L=0.06u
MPA2_2 INT B VDD VNW PCH W=0.47u L=0.06u
MNA104_5 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_5 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_6 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_6 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AND2X6MA10TR

****
.SUBCKT NAND2X6MA10TR VDD VSS VPW VNW Y A B
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_5 VSS B N_31 VPW NCH W=0.58u L=0.06u
MPA1_6 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_5 Y A N_31 VPW NCH W=0.58u L=0.06u
MNA1_6 Y A N_33 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_4 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_6 VSS B N_33 VPW NCH W=0.58u L=0.06u
MNA2 VSS B N_35 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1 Y A N_35 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y A N_37 VPW NCH W=0.58u L=0.06u
MPA1_5 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_6 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_3 VSS B N_37 VPW NCH W=0.58u L=0.06u
MNA2_4 VSS B N_39 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_4 Y A N_39 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y A N_29 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_2 N_29 B VSS VPW NCH W=0.58u L=0.06u
MPA2_5 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2X6MA10TR

****
.SUBCKT AND2X8MA10TR VDD VSS VPW VNW Y A B
MPA2_4 INT B VDD VNW PCH W=0.47u L=0.06u
MNA2 VSS B N_22 VPW NCH W=0.575u L=0.06u
MPA1_4 INT A VDD VNW PCH W=0.47u L=0.06u
MNA1 INT A N_22 VPW NCH W=0.575u L=0.06u
MPA1_2 INT A VDD VNW PCH W=0.475u L=0.06u
MNA1_3 INT A N_24 VPW NCH W=0.575u L=0.06u
MPA2_3 INT B VDD VNW PCH W=0.475u L=0.06u
MNA2_3 N_24 B VSS VPW NCH W=0.575u L=0.06u
MNA2_4 VSS B N_26 VPW NCH W=0.58u L=0.06u
MPA2_2 INT B VDD VNW PCH W=0.475u L=0.06u
MNA1_4 INT A N_26 VPW NCH W=0.58u L=0.06u
MPA1_3 INT A VDD VNW PCH W=0.475u L=0.06u
MNA1_2 INT A N_29 VPW NCH W=0.58u L=0.06u
MPA1 INT A VDD VNW PCH W=0.475u L=0.06u
MNA2_2 N_29 B VSS VPW NCH W=0.58u L=0.06u
MPA2 INT B VDD VNW PCH W=0.475u L=0.06u
MNA104_5 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_5 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_7 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_7 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_6 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_6 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_8 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_8 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AND2X8MA10TR

****
.SUBCKT NAND2X8MA10TR VDD VSS VPW VNW Y A B
MPA2_8 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS B N_39 VPW NCH W=0.58u L=0.06u
MPA1_8 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1 Y A N_39 VPW NCH W=0.58u L=0.06u
MNA1_8 Y A N_41 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_7 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_8 VSS B N_41 VPW NCH W=0.58u L=0.06u
MNA2_2 VSS B N_43 VPW NCH W=0.58u L=0.06u
MPA2_4 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y A N_43 VPW NCH W=0.58u L=0.06u
MPA1_7 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_6 Y A N_45 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_6 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_6 VSS B N_45 VPW NCH W=0.58u L=0.06u
MNA2_7 VSS B N_47 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_7 Y A N_47 VPW NCH W=0.58u L=0.06u
MPA1_6 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_4 Y A N_49 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_5 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_4 VSS B N_49 VPW NCH W=0.58u L=0.06u
MNA2_5 VSS B N_51 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_5 Y A N_51 VPW NCH W=0.58u L=0.06u
MPA1_5 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y A N_37 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_3 N_37 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2X8MA10TR

****
.SUBCKT AND3X2MA10TR VDD VSS VPW VNW Y A B C
MNA3 N_17 C VSS VPW NCH W=0.47u L=0.06u
MNA2 N_17 B N_18 VPW NCH W=0.47u L=0.06u
MNA102 N_18 A INT VPW NCH W=0.47u L=0.06u
MPA105 INT A VDD VNW PCH W=0.58u L=0.06u
MNA102_2 INT A N_20 VPW NCH W=0.475u L=0.06u
MNA2_2 N_20 B N_21 VPW NCH W=0.475u L=0.06u
MPA2 INT B VDD VNW PCH W=0.58u L=0.06u
MNA3_2 N_21 C VSS VPW NCH W=0.475u L=0.06u
MPA3 INT C VDD VNW PCH W=0.58u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AND3X2MA10TR

****
.SUBCKT NAND3X2MA10TR VDD VSS VPW VNW Y A B C
MPA3_2 Y C VDD VNW PCH W=0.36u L=0.06u
MNA3 VSS C N_19 VPW NCH W=0.58u L=0.06u
MNA2 N_19 B N_20 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.36u L=0.06u
MNA1 Y A N_20 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.36u L=0.06u
MNA1_2 Y A N_22 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.36u L=0.06u
MNA2_2 N_22 B N_17 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.36u L=0.06u
MNA3_2 N_17 C VSS VPW NCH W=0.58u L=0.06u
MPA3 Y C VDD VNW PCH W=0.36u L=0.06u
.ENDS NAND3X2MA10TR

****
.SUBCKT AND3X3MA10TR VDD VSS VPW VNW Y A B C
MNA102 INT A N_25 VPW NCH W=0.45u L=0.06u
MNA2 N_25 B N_26 VPW NCH W=0.45u L=0.06u
MPA3 INT C VDD VNW PCH W=0.415u L=0.06u
MNA3 VSS C N_26 VPW NCH W=0.45u L=0.06u
MNA3_3 VSS C N_28 VPW NCH W=0.45u L=0.06u
MPA2_2 INT B VDD VNW PCH W=0.415u L=0.06u
MNA2_3 N_28 B N_29 VPW NCH W=0.45u L=0.06u
MPA105 INT A VDD VNW PCH W=0.415u L=0.06u
MNA102_3 N_29 A INT VPW NCH W=0.45u L=0.06u
MPA105_2 INT A VDD VNW PCH W=0.415u L=0.06u
MNA102_2 INT A N_31 VPW NCH W=0.455u L=0.06u
MNA2_2 N_31 B N_32 VPW NCH W=0.455u L=0.06u
MPA2 INT B VDD VNW PCH W=0.415u L=0.06u
MNA3_2 N_32 C VSS VPW NCH W=0.455u L=0.06u
MPA3_2 INT C VDD VNW PCH W=0.415u L=0.06u
MNA1_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AND3X3MA10TR

****
.SUBCKT NAND3X3MA10TR VDD VSS VPW VNW Y A B C
MNA3_2 N_15 C VSS VPW NCH W=0.58u L=0.06u
MPA3 Y C VDD VNW PCH W=0.36u L=0.06u
MNA3 VSS C N_15 VPW NCH W=0.58u L=0.06u
MPA3_3 Y C VDD VNW PCH W=0.36u L=0.06u
MNA3_3 VSS C N_15 VPW NCH W=0.58u L=0.06u
MPA3_2 Y C VDD VNW PCH W=0.36u L=0.06u
MNA2 N_13 B N_15 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.36u L=0.06u
MNA2_3 N_15 B N_13 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.36u L=0.06u
MNA2_2 N_15 B N_13 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.36u L=0.06u
MNA1_2 Y A N_13 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.36u L=0.06u
MNA1 N_13 A Y VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.36u L=0.06u
MNA1_3 Y A N_13 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.36u L=0.06u
.ENDS NAND3X3MA10TR

****
.SUBCKT AND4X1P4MA10TR VDD VSS VPW VNW Y A B C D
MPA4_2 INT D VDD VNW PCH W=0.255u L=0.06u
MNA4_2 VSS D N_27 VPW NCH W=0.5u L=0.06u
MPA3 INT C VDD VNW PCH W=0.255u L=0.06u
MNA3_2 N_27 C N_28 VPW NCH W=0.5u L=0.06u
MNA2_2 N_28 B N_29 VPW NCH W=0.5u L=0.06u
MPA2_2 INT B VDD VNW PCH W=0.255u L=0.06u
MNA102_2 INT A N_29 VPW NCH W=0.5u L=0.06u
MPA105 INT A VDD VNW PCH W=0.255u L=0.06u
MNA102 INT A N_31 VPW NCH W=0.5u L=0.06u
MPA105_2 INT A VDD VNW PCH W=0.255u L=0.06u
MNA2 N_31 B N_32 VPW NCH W=0.5u L=0.06u
MPA2 INT B VDD VNW PCH W=0.255u L=0.06u
MNA3 N_32 C N_33 VPW NCH W=0.5u L=0.06u
MPA3_2 INT C VDD VNW PCH W=0.255u L=0.06u
MNA4 N_33 D VSS VPW NCH W=0.5u L=0.06u
MPA4 INT D VDD VNW PCH W=0.255u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS AND4X1P4MA10TR

****
.SUBCKT NAND4X1P4MA10TR VDD VSS VPW VNW Y A B C D
MPA4_2 Y D VDD VNW PCH W=0.2u L=0.06u
MNA4 VSS D N_23 VPW NCH W=0.41u L=0.06u
MPA3 Y C VDD VNW PCH W=0.2u L=0.06u
MNA3 N_23 C N_24 VPW NCH W=0.41u L=0.06u
MNA2 N_24 B N_25 VPW NCH W=0.41u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.2u L=0.06u
MNA1 Y A N_25 VPW NCH W=0.41u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.2u L=0.06u
MNA1_2 Y A N_27 VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.2u L=0.06u
MNA2_2 N_27 B N_28 VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.2u L=0.06u
MNA3_2 N_28 C N_21 VPW NCH W=0.41u L=0.06u
MPA3_2 Y C VDD VNW PCH W=0.2u L=0.06u
MNA4_2 N_21 D VSS VPW NCH W=0.41u L=0.06u
MPA4 Y D VDD VNW PCH W=0.2u L=0.06u
.ENDS NAND4X1P4MA10TR

****
.SUBCKT AO1B2X1P4MA10TR VDD VSS VPW VNW Y A0N B0 B1
MPA1 INT B0 VDD VNW PCH W=0.41u L=0.06u
MNA1 INT B0 N_19 VPW NCH W=0.335u L=0.06u
MPA2 INT B1 VDD VNW PCH W=0.41u L=0.06u
MNA2 N_19 B1 VSS VPW NCH W=0.335u L=0.06u
MNA206 VSS A0N N_21 VPW NCH W=0.405u L=0.06u
MPA2010_2 Y A0N VDD VNW PCH W=0.49u L=0.06u
MNA104 Y INT N_21 VPW NCH W=0.405u L=0.06u
MPA108_2 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA104_2 Y INT N_17 VPW NCH W=0.405u L=0.06u
MPA108 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA206_2 N_17 A0N VSS VPW NCH W=0.405u L=0.06u
MPA2010 Y A0N VDD VNW PCH W=0.49u L=0.06u
.ENDS AO1B2X1P4MA10TR

****
.SUBCKT AO1B2X2MA10TR VDD VSS VPW VNW Y A0N B0 B1
MPA1 INT B0 VDD VNW PCH W=0.55u L=0.06u
MNA1 INT B0 N_19 VPW NCH W=0.45u L=0.06u
MPA2 INT B1 VDD VNW PCH W=0.55u L=0.06u
MNA2 N_19 B1 VSS VPW NCH W=0.45u L=0.06u
MNA206 VSS A0N N_21 VPW NCH W=0.575u L=0.06u
MPA2010_2 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT N_21 VPW NCH W=0.575u L=0.06u
MPA108_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT N_17 VPW NCH W=0.575u L=0.06u
MPA108 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA206_2 N_17 A0N VSS VPW NCH W=0.575u L=0.06u
MPA2010 Y A0N VDD VNW PCH W=0.7u L=0.06u
.ENDS AO1B2X2MA10TR

****
.SUBCKT AO1B2X3MA10TR VDD VSS VPW VNW Y A0N B0 B1
MNA2_2 VSS B1 N_27 VPW NCH W=0.345u L=0.06u
MPA2_2 INT B1 VDD VNW PCH W=0.42u L=0.06u
MNA1_2 INT B0 N_27 VPW NCH W=0.345u L=0.06u
MPA1_2 INT B0 VDD VNW PCH W=0.42u L=0.06u
MNA1 INT B0 N_29 VPW NCH W=0.345u L=0.06u
MPA1 INT B0 VDD VNW PCH W=0.42u L=0.06u
MPA2 INT B1 VDD VNW PCH W=0.42u L=0.06u
MNA2 N_29 B1 VSS VPW NCH W=0.345u L=0.06u
MNA206_2 VSS A0N N_31 VPW NCH W=0.575u L=0.06u
MPA2010_2 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT N_31 VPW NCH W=0.575u L=0.06u
MPA108_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT N_33 VPW NCH W=0.575u L=0.06u
MPA108 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA2010_3 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA206 VSS A0N N_33 VPW NCH W=0.575u L=0.06u
MNA206_3 VSS A0N N_25 VPW NCH W=0.575u L=0.06u
MPA2010 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA104_3 N_25 INT Y VPW NCH W=0.575u L=0.06u
MPA108_2 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AO1B2X3MA10TR

****
.SUBCKT AO1B2X4MA10TR VDD VSS VPW VNW Y A0N B0 B1
MNA2 VSS B1 N_31 VPW NCH W=0.45u L=0.06u
MPA2_2 INT B1 VDD VNW PCH W=0.55u L=0.06u
MNA1 INT B0 N_31 VPW NCH W=0.45u L=0.06u
MPA1_2 INT B0 VDD VNW PCH W=0.55u L=0.06u
MNA1_2 INT B0 N_33 VPW NCH W=0.45u L=0.06u
MPA1 INT B0 VDD VNW PCH W=0.55u L=0.06u
MPA2 INT B1 VDD VNW PCH W=0.55u L=0.06u
MNA2_2 N_33 B1 VSS VPW NCH W=0.45u L=0.06u
MNA206 VSS A0N N_35 VPW NCH W=0.575u L=0.06u
MPA2010_2 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT N_35 VPW NCH W=0.575u L=0.06u
MPA108_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT N_37 VPW NCH W=0.575u L=0.06u
MPA108_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA2010_4 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA206_2 VSS A0N N_37 VPW NCH W=0.575u L=0.06u
MNA206_3 VSS A0N N_39 VPW NCH W=0.575u L=0.06u
MPA2010 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT N_39 VPW NCH W=0.575u L=0.06u
MPA108_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y INT N_29 VPW NCH W=0.575u L=0.06u
MPA108 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA206_4 N_29 A0N VSS VPW NCH W=0.575u L=0.06u
MPA2010_3 Y A0N VDD VNW PCH W=0.7u L=0.06u
.ENDS AO1B2X4MA10TR

****
.SUBCKT AO1B2X6MA10TR VDD VSS VPW VNW Y A0N B0 B1
MNA1_3 INT B0 N_43 VPW NCH W=0.45u L=0.06u
MPA1_3 INT B0 VDD VNW PCH W=0.55u L=0.06u
MPA2_3 INT B1 VDD VNW PCH W=0.55u L=0.06u
MNA2_3 VSS B1 N_43 VPW NCH W=0.45u L=0.06u
MNA2_2 VSS B1 N_45 VPW NCH W=0.45u L=0.06u
MPA2_2 INT B1 VDD VNW PCH W=0.55u L=0.06u
MNA1_2 INT B0 N_45 VPW NCH W=0.45u L=0.06u
MPA1_2 INT B0 VDD VNW PCH W=0.55u L=0.06u
MNA1 INT B0 N_47 VPW NCH W=0.45u L=0.06u
MPA1 INT B0 VDD VNW PCH W=0.55u L=0.06u
MPA2 INT B1 VDD VNW PCH W=0.55u L=0.06u
MNA2 N_47 B1 VSS VPW NCH W=0.45u L=0.06u
MNA206_4 VSS A0N N_49 VPW NCH W=0.575u L=0.06u
MPA2010_6 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y INT N_49 VPW NCH W=0.575u L=0.06u
MPA108_6 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT N_51 VPW NCH W=0.575u L=0.06u
MPA108_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA2010_5 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA206_3 VSS A0N N_51 VPW NCH W=0.575u L=0.06u
MNA206_2 VSS A0N N_53 VPW NCH W=0.575u L=0.06u
MPA2010_3 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT N_53 VPW NCH W=0.575u L=0.06u
MPA108_5 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT N_55 VPW NCH W=0.575u L=0.06u
MPA108_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MPA2010_4 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA206 VSS A0N N_55 VPW NCH W=0.575u L=0.06u
MNA206_6 VSS A0N N_57 VPW NCH W=0.575u L=0.06u
MPA2010_2 Y A0N VDD VNW PCH W=0.7u L=0.06u
MNA104_6 Y INT N_57 VPW NCH W=0.575u L=0.06u
MPA108_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_5 Y INT N_41 VPW NCH W=0.575u L=0.06u
MPA108 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA206_5 N_41 A0N VSS VPW NCH W=0.575u L=0.06u
MPA2010 Y A0N VDD VNW PCH W=0.7u L=0.06u
.ENDS AO1B2X6MA10TR

****
.SUBCKT AO21BX1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0N
MPA1 INT A0 VDD VNW PCH W=0.41u L=0.06u
MNA1 INT A0 N_19 VPW NCH W=0.335u L=0.06u
MPA2 INT A1 VDD VNW PCH W=0.41u L=0.06u
MNA2 N_19 A1 VSS VPW NCH W=0.335u L=0.06u
MNA206 VSS INT N_21 VPW NCH W=0.405u L=0.06u
MPA2010_2 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA104 Y B0N N_21 VPW NCH W=0.405u L=0.06u
MPA108_2 Y B0N VDD VNW PCH W=0.49u L=0.06u
MNA104_2 Y B0N N_17 VPW NCH W=0.405u L=0.06u
MPA108 Y B0N VDD VNW PCH W=0.49u L=0.06u
MNA206_2 N_17 INT VSS VPW NCH W=0.405u L=0.06u
MPA2010 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS AO21BX1P4MA10TR

****
.SUBCKT AO21BX2MA10TR VDD VSS VPW VNW Y A0 A1 B0N
MPA1 INT A0 VDD VNW PCH W=0.55u L=0.06u
MNA1 INT A0 N_19 VPW NCH W=0.45u L=0.06u
MPA2 INT A1 VDD VNW PCH W=0.55u L=0.06u
MNA2 N_19 A1 VSS VPW NCH W=0.45u L=0.06u
MNA206 VSS INT N_21 VPW NCH W=0.575u L=0.06u
MPA2010_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y B0N N_21 VPW NCH W=0.575u L=0.06u
MPA108_2 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y B0N N_17 VPW NCH W=0.575u L=0.06u
MPA108 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA206_2 N_17 INT VSS VPW NCH W=0.575u L=0.06u
MPA2010 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AO21BX2MA10TR

****
.SUBCKT AO21BX3MA10TR VDD VSS VPW VNW Y A0 A1 B0N
MNA2_2 VSS A1 N_27 VPW NCH W=0.345u L=0.06u
MPA2_2 INT A1 VDD VNW PCH W=0.42u L=0.06u
MNA1_2 INT A0 N_27 VPW NCH W=0.345u L=0.06u
MPA1_2 INT A0 VDD VNW PCH W=0.42u L=0.06u
MNA1 INT A0 N_29 VPW NCH W=0.345u L=0.06u
MPA1 INT A0 VDD VNW PCH W=0.42u L=0.06u
MPA2 INT A1 VDD VNW PCH W=0.42u L=0.06u
MNA2 N_29 A1 VSS VPW NCH W=0.345u L=0.06u
MNA206_2 VSS INT N_31 VPW NCH W=0.575u L=0.06u
MPA2010_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y B0N N_31 VPW NCH W=0.575u L=0.06u
MPA108_3 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA104 Y B0N N_33 VPW NCH W=0.575u L=0.06u
MPA108 Y B0N VDD VNW PCH W=0.7u L=0.06u
MPA2010_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA206 VSS INT N_33 VPW NCH W=0.575u L=0.06u
MNA206_3 VSS INT N_25 VPW NCH W=0.575u L=0.06u
MPA2010 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 N_25 B0N Y VPW NCH W=0.575u L=0.06u
MPA108_2 Y B0N VDD VNW PCH W=0.7u L=0.06u
.ENDS AO21BX3MA10TR

****
.SUBCKT AO21BX4MA10TR VDD VSS VPW VNW Y A0 A1 B0N
MNA2 VSS A1 N_31 VPW NCH W=0.45u L=0.06u
MPA2_2 INT A1 VDD VNW PCH W=0.55u L=0.06u
MNA1 INT A0 N_31 VPW NCH W=0.45u L=0.06u
MPA1_2 INT A0 VDD VNW PCH W=0.55u L=0.06u
MNA1_2 INT A0 N_33 VPW NCH W=0.45u L=0.06u
MPA1 INT A0 VDD VNW PCH W=0.55u L=0.06u
MPA2 INT A1 VDD VNW PCH W=0.55u L=0.06u
MNA2_2 N_33 A1 VSS VPW NCH W=0.45u L=0.06u
MNA206 VSS INT N_35 VPW NCH W=0.575u L=0.06u
MPA2010_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y B0N N_35 VPW NCH W=0.575u L=0.06u
MPA108_2 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y B0N N_37 VPW NCH W=0.575u L=0.06u
MPA108_4 Y B0N VDD VNW PCH W=0.7u L=0.06u
MPA2010_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA206_2 VSS INT N_37 VPW NCH W=0.575u L=0.06u
MNA206_3 VSS INT N_39 VPW NCH W=0.575u L=0.06u
MPA2010 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y B0N N_39 VPW NCH W=0.575u L=0.06u
MPA108_3 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y B0N N_29 VPW NCH W=0.575u L=0.06u
MPA108 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA206_4 N_29 INT VSS VPW NCH W=0.575u L=0.06u
MPA2010_3 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AO21BX4MA10TR

****
.SUBCKT AO21BX6MA10TR VDD VSS VPW VNW Y A0 A1 B0N
MNA1_3 INT A0 N_43 VPW NCH W=0.45u L=0.06u
MPA1_3 INT A0 VDD VNW PCH W=0.55u L=0.06u
MPA2_3 INT A1 VDD VNW PCH W=0.55u L=0.06u
MNA2_3 VSS A1 N_43 VPW NCH W=0.45u L=0.06u
MNA2_2 VSS A1 N_45 VPW NCH W=0.45u L=0.06u
MPA2_2 INT A1 VDD VNW PCH W=0.55u L=0.06u
MNA1_2 INT A0 N_45 VPW NCH W=0.45u L=0.06u
MPA1_2 INT A0 VDD VNW PCH W=0.55u L=0.06u
MNA1 INT A0 N_47 VPW NCH W=0.45u L=0.06u
MPA1 INT A0 VDD VNW PCH W=0.55u L=0.06u
MPA2 INT A1 VDD VNW PCH W=0.55u L=0.06u
MNA2 N_47 A1 VSS VPW NCH W=0.45u L=0.06u
MNA206_4 VSS INT N_49 VPW NCH W=0.575u L=0.06u
MPA2010_6 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y B0N N_49 VPW NCH W=0.575u L=0.06u
MPA108_6 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y B0N N_51 VPW NCH W=0.575u L=0.06u
MPA108_3 Y B0N VDD VNW PCH W=0.7u L=0.06u
MPA2010_5 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA206_3 VSS INT N_51 VPW NCH W=0.575u L=0.06u
MNA206_2 VSS INT N_53 VPW NCH W=0.575u L=0.06u
MPA2010_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y B0N N_53 VPW NCH W=0.575u L=0.06u
MPA108_5 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA104 Y B0N N_55 VPW NCH W=0.575u L=0.06u
MPA108_2 Y B0N VDD VNW PCH W=0.7u L=0.06u
MPA2010_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA206 VSS INT N_55 VPW NCH W=0.575u L=0.06u
MNA206_6 VSS INT N_57 VPW NCH W=0.575u L=0.06u
MPA2010_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_6 Y B0N N_57 VPW NCH W=0.575u L=0.06u
MPA108_4 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA104_5 Y B0N N_41 VPW NCH W=0.575u L=0.06u
MPA108 Y B0N VDD VNW PCH W=0.7u L=0.06u
MNA206_5 N_41 INT VSS VPW NCH W=0.575u L=0.06u
MPA2010 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AO21BX6MA10TR

****
.SUBCKT AO21X2MA10TR VDD VSS VPW VNW Y A0 A1 B0
MNB2_2 VSS A1 N_25 VPW NCH W=0.36u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.53u L=0.06u
MNB1_2 INT A0 N_25 VPW NCH W=0.36u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.53u L=0.06u
MNB1 N_27 A0 INT VPW NCH W=0.36u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.53u L=0.06u
MNB2 VSS A1 N_27 VPW NCH W=0.36u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.53u L=0.06u
MNA106 INT B0 VSS VPW NCH W=0.435u L=0.06u
MPA108_2 INT B0 P1 VNW PCH W=0.53u L=0.06u
MPA108 INT B0 P1 VNW PCH W=0.53u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AO21X2MA10TR

****
.SUBCKT AO21X3MA10TR VDD VSS VPW VNW Y A0 A1 B0
MPB1_2 P1 A0 VDD VNW PCH W=0.52u L=0.06u
MNB1_2 INT A0 N_33 VPW NCH W=0.35u L=0.06u
MPB2_3 P1 A1 VDD VNW PCH W=0.515u L=0.06u
MNB2_2 VSS A1 N_33 VPW NCH W=0.35u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.515u L=0.06u
MNB2_3 VSS A1 N_35 VPW NCH W=0.35u L=0.06u
MPB1_3 P1 A0 VDD VNW PCH W=0.515u L=0.06u
MNB1_3 INT A0 N_35 VPW NCH W=0.35u L=0.06u
MNB1 INT A0 N_38 VPW NCH W=0.35u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.515u L=0.06u
MNB2 N_38 A1 VSS VPW NCH W=0.35u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.52u L=0.06u
MNA106_2 INT B0 VSS VPW NCH W=0.32u L=0.06u
MPA108_3 INT B0 P1 VNW PCH W=0.52u L=0.06u
MNA106 INT B0 VSS VPW NCH W=0.315u L=0.06u
MPA108_2 INT B0 P1 VNW PCH W=0.515u L=0.06u
MPA108 INT B0 P1 VNW PCH W=0.515u L=0.06u
MNA1_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AO21X3MA10TR

****
.SUBCKT AO21X4MA10TR VDD VSS VPW VNW Y A0 A1 B0
MPB2_3 P1 A1 VDD VNW PCH W=0.68u L=0.06u
MNB2_3 VSS A1 N_20 VPW NCH W=0.46u L=0.06u
MPB1_3 P1 A0 VDD VNW PCH W=0.685u L=0.06u
MNB1_3 N_20 A0 INT VPW NCH W=0.46u L=0.06u
MNB1 INT A0 N_22 VPW NCH W=0.465u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.685u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.685u L=0.06u
MNB2 VSS A1 N_22 VPW NCH W=0.465u L=0.06u
MNB2_2 VSS A1 N_25 VPW NCH W=0.465u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.685u L=0.06u
MNB1_2 N_25 A0 INT VPW NCH W=0.465u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.68u L=0.06u
MNA106 INT B0 VSS VPW NCH W=0.42u L=0.06u
MPA108_2 INT B0 P1 VNW PCH W=0.685u L=0.06u
MNA106_2 INT B0 VSS VPW NCH W=0.42u L=0.06u
MPA108 INT B0 P1 VNW PCH W=0.685u L=0.06u
MPA108_3 INT B0 P1 VNW PCH W=0.68u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_4 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AO21X4MA10TR

****
.SUBCKT AO22X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1
MNB2_2 VSS A1 N_29 VPW NCH W=0.28u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.42u L=0.06u
MNB1_2 INT A0 N_29 VPW NCH W=0.28u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.42u L=0.06u
MNB1 INT A0 N_31 VPW NCH W=0.28u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.42u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.42u L=0.06u
MNB2 N_31 A1 VSS VPW NCH W=0.28u L=0.06u
MNA2 VSS B1 N_33 VPW NCH W=0.28u L=0.06u
MPA2_2 INT B1 P1 VNW PCH W=0.42u L=0.06u
MNA106 INT B0 N_33 VPW NCH W=0.28u L=0.06u
MPA109_2 INT B0 P1 VNW PCH W=0.42u L=0.06u
MNA106_2 INT B0 N_27 VPW NCH W=0.28u L=0.06u
MPA109 INT B0 P1 VNW PCH W=0.42u L=0.06u
MNA2_2 N_27 B1 VSS VPW NCH W=0.28u L=0.06u
MPA2 INT B1 P1 VNW PCH W=0.42u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS AO22X1P4MA10TR

****
.SUBCKT AO22X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1
MNB2_2 VSS A1 N_29 VPW NCH W=0.38u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.575u L=0.06u
MNB1_2 INT A0 N_29 VPW NCH W=0.38u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.575u L=0.06u
MNB1 INT A0 N_31 VPW NCH W=0.38u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.57u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.57u L=0.06u
MNB2 N_31 A1 VSS VPW NCH W=0.38u L=0.06u
MNA2 VSS B1 N_33 VPW NCH W=0.38u L=0.06u
MPA2_2 INT B1 P1 VNW PCH W=0.57u L=0.06u
MNA106 INT B0 N_33 VPW NCH W=0.38u L=0.06u
MPA109_2 INT B0 P1 VNW PCH W=0.57u L=0.06u
MNA106_2 INT B0 N_27 VPW NCH W=0.38u L=0.06u
MPA109 INT B0 P1 VNW PCH W=0.575u L=0.06u
MNA2_2 N_27 B1 VSS VPW NCH W=0.38u L=0.06u
MPA2 INT B1 P1 VNW PCH W=0.575u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS AO22X2MA10TR

****
.SUBCKT AOI211X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MN5 VSS A1 N_23 VPW NCH W=0.23u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
MN4 Y A0 N_23 VPW NCH W=0.23u L=0.06u
MP5_2 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MN4_2 Y A0 N_25 VPW NCH W=0.23u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MN5_2 N_25 A1 VSS VPW NCH W=0.23u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.49u L=0.06u
MP2 P1 B0 N_9 VNW PCH W=0.49u L=0.06u
MN3 Y B0 VSS VPW NCH W=0.29u L=0.06u
MN0 Y C0 VSS VPW NCH W=0.29u L=0.06u
MP1 Y C0 N_9 VNW PCH W=0.49u L=0.06u
MP1_2 Y C0 N_3 VNW PCH W=0.49u L=0.06u
MP2_2 N_3 B0 P1 VNW PCH W=0.49u L=0.06u
.ENDS AOI211X1P4MA10TR

****
.SUBCKT AOI211X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MN5 VSS A1 N_23 VPW NCH W=0.33u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4 Y A0 N_23 VPW NCH W=0.33u L=0.06u
MP5_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4_2 Y A0 N_25 VPW NCH W=0.33u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN5_2 N_25 A1 VSS VPW NCH W=0.33u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MP2 P1 B0 N_9 VNW PCH W=0.7u L=0.06u
MN3 Y B0 VSS VPW NCH W=0.41u L=0.06u
MN0 Y C0 VSS VPW NCH W=0.41u L=0.06u
MP1 Y C0 N_9 VNW PCH W=0.7u L=0.06u
MP1_2 Y C0 N_3 VNW PCH W=0.7u L=0.06u
MP2_2 N_3 B0 P1 VNW PCH W=0.7u L=0.06u
.ENDS AOI211X2MA10TR

****
.SUBCKT AOI211X3MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MP5_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4_3 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5_2 VSS A1 N_18 VPW NCH W=0.495u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4_2 Y A0 N_18 VPW NCH W=0.495u L=0.06u
MP5_3 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4 Y A0 N_21 VPW NCH W=0.495u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN5 N_21 A1 VSS VPW NCH W=0.495u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MP2_2 P1 B0 N_11 VNW PCH W=0.7u L=0.06u
MN3_2 Y B0 VSS VPW NCH W=0.305u L=0.06u
MP1_2 Y C0 N_11 VNW PCH W=0.7u L=0.06u
MN0_2 Y C0 VSS VPW NCH W=0.305u L=0.06u
MP1 Y C0 N_13 VNW PCH W=0.7u L=0.06u
MN0 Y C0 VSS VPW NCH W=0.31u L=0.06u
MP2 P1 B0 N_13 VNW PCH W=0.7u L=0.06u
MN3 Y B0 VSS VPW NCH W=0.31u L=0.06u
MP2_3 P1 B0 N_3 VNW PCH W=0.7u L=0.06u
MP1_3 N_3 C0 Y VNW PCH W=0.7u L=0.06u
.ENDS AOI211X3MA10TR

****
.SUBCKT AOI211X4MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MP4_4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MP5_3 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4_3 Y A0 N_39 VPW NCH W=0.44u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5_3 VSS A1 N_39 VPW NCH W=0.44u L=0.06u
MN5_2 VSS A1 N_41 VPW NCH W=0.44u L=0.06u
MP4_3 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4_2 Y A0 N_41 VPW NCH W=0.44u L=0.06u
MP5_4 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4 Y A0 N_44 VPW NCH W=0.44u L=0.06u
MP5_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN5 N_44 A1 VSS VPW NCH W=0.44u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MP2_3 P1 B0 N_13 VNW PCH W=0.7u L=0.06u
MN3_2 Y B0 VSS VPW NCH W=0.41u L=0.06u
MP1_3 Y C0 N_13 VNW PCH W=0.7u L=0.06u
MN0 Y C0 VSS VPW NCH W=0.41u L=0.06u
MP1 Y C0 N_15 VNW PCH W=0.7u L=0.06u
MN0_2 Y C0 VSS VPW NCH W=0.41u L=0.06u
MP2 P1 B0 N_15 VNW PCH W=0.7u L=0.06u
MN3 Y B0 VSS VPW NCH W=0.41u L=0.06u
MP2_2 P1 B0 N_17 VNW PCH W=0.7u L=0.06u
MP1_2 Y C0 N_17 VNW PCH W=0.7u L=0.06u
MP1_4 Y C0 N_3 VNW PCH W=0.7u L=0.06u
MP2_4 N_3 B0 P1 VNW PCH W=0.7u L=0.06u
.ENDS AOI211X4MA10TR

****
.SUBCKT AOI21BX1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0N
MNB2 VSS A1 N_23 VPW NCH W=0.32u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
MNB1 Y A0 N_23 VPW NCH W=0.32u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MNB1_2 Y A0 N_25 VPW NCH W=0.32u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MNB2_2 N_25 A1 VSS VPW NCH W=0.32u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
MNA106_2 Y NET28 VSS VPW NCH W=0.2u L=0.06u
MPA108 Y NET28 P1 VNW PCH W=0.49u L=0.06u
MNA106 Y NET28 VSS VPW NCH W=0.2u L=0.06u
MPA108_2 Y NET28 P1 VNW PCH W=0.49u L=0.06u
MNA1 NET28 B0N VSS VPW NCH W=0.21u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.275u L=0.06u
.ENDS AOI21BX1P4MA10TR

****
.SUBCKT AOI21BX2MA10TR VDD VSS VPW VNW Y A0 A1 B0N
MNB2 VSS A1 N_23 VPW NCH W=0.455u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MNB1 Y A0 N_23 VPW NCH W=0.455u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MNB1_2 Y A0 N_25 VPW NCH W=0.455u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MNB2_2 N_25 A1 VSS VPW NCH W=0.455u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MNA106_2 Y NET28 VSS VPW NCH W=0.285u L=0.06u
MPA108 Y NET28 P1 VNW PCH W=0.7u L=0.06u
MNA106 Y NET28 VSS VPW NCH W=0.285u L=0.06u
MPA108_2 Y NET28 P1 VNW PCH W=0.7u L=0.06u
MNA1 NET28 B0N VSS VPW NCH W=0.27u L=0.06u
MPA1 NET28 B0N VDD VNW PCH W=0.36u L=0.06u
.ENDS AOI21BX2MA10TR

****
.SUBCKT AOI21X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0
MNB2 VSS A1 N_19 VPW NCH W=0.32u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
MNB1 Y A0 N_19 VPW NCH W=0.32u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MNB1_2 Y A0 N_21 VPW NCH W=0.32u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MNB2_2 N_21 A1 VSS VPW NCH W=0.32u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
MNA1_2 Y B0 VSS VPW NCH W=0.2u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.49u L=0.06u
MNA1 Y B0 VSS VPW NCH W=0.2u L=0.06u
MPA1_2 Y B0 P1 VNW PCH W=0.49u L=0.06u
.ENDS AOI21X1P4MA10TR

****
.SUBCKT AOI21X2MA10TR VDD VSS VPW VNW Y A0 A1 B0
MNB2 VSS A1 N_19 VPW NCH W=0.455u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MNB1 Y A0 N_19 VPW NCH W=0.455u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MNB1_2 Y A0 N_21 VPW NCH W=0.455u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MNB2_2 N_21 A1 VSS VPW NCH W=0.455u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y B0 VSS VPW NCH W=0.285u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.7u L=0.06u
MNA1 Y B0 VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y B0 P1 VNW PCH W=0.7u L=0.06u
.ENDS AOI21X2MA10TR

****
.SUBCKT AOI221X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0
MN5_2 VSS A1 N_29 VPW NCH W=0.33u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4_2 Y A0 N_29 VPW NCH W=0.33u L=0.06u
MP5_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4 Y A0 N_27 VPW NCH W=0.33u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN5 N_27 A1 VSS VPW NCH W=0.33u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN2_2 VSS B1 N_34 VPW NCH W=0.33u L=0.06u
MP3_2 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN3_2 Y B0 N_34 VPW NCH W=0.33u L=0.06u
MP2_2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN3 Y B0 N_36 VPW NCH W=0.33u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN2 N_36 B1 VSS VPW NCH W=0.33u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN0 Y C0 VSS VPW NCH W=0.41u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.7u L=0.06u
MP1_2 Y C0 P2 VNW PCH W=0.7u L=0.06u
.ENDS AOI221X2MA10TR

****
.SUBCKT AOI221X3MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0
MP5_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4_3 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5_2 VSS A1 N_22 VPW NCH W=0.495u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4_2 Y A0 N_22 VPW NCH W=0.495u L=0.06u
MP5_3 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4 Y A0 N_24 VPW NCH W=0.495u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5 N_24 A1 VSS VPW NCH W=0.495u L=0.06u
MN2_2 VSS B1 N_26 VPW NCH W=0.495u L=0.06u
MP3_2 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN3_2 Y B0 N_26 VPW NCH W=0.495u L=0.06u
MP2_3 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN3 Y B0 N_20 VPW NCH W=0.495u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN2 N_20 B1 VSS VPW NCH W=0.495u L=0.06u
MP3_3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MP2_2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN0_2 Y C0 VSS VPW NCH W=0.31u L=0.06u
MP1_3 Y C0 P2 VNW PCH W=0.7u L=0.06u
MN0 Y C0 VSS VPW NCH W=0.305u L=0.06u
MP1_2 Y C0 P2 VNW PCH W=0.7u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.7u L=0.06u
.ENDS AOI221X3MA10TR

****
.SUBCKT AOI221X4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0
MN5_4 VSS A1 N_49 VPW NCH W=0.33u L=0.06u
MP4_4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4_4 Y A0 N_49 VPW NCH W=0.33u L=0.06u
MP5_4 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4_3 Y A0 N_51 VPW NCH W=0.33u L=0.06u
MP5_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4_3 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5_3 VSS A1 N_51 VPW NCH W=0.33u L=0.06u
MN5_2 VSS A1 N_53 VPW NCH W=0.33u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4_2 Y A0 N_53 VPW NCH W=0.33u L=0.06u
MP5_3 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4 Y A0 N_47 VPW NCH W=0.33u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN5 N_47 A1 VSS VPW NCH W=0.33u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN2_4 VSS B1 N_58 VPW NCH W=0.33u L=0.06u
MP3_4 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN3_4 Y B0 N_58 VPW NCH W=0.33u L=0.06u
MP2_4 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN3_3 Y B0 N_60 VPW NCH W=0.33u L=0.06u
MP2_2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MP3_3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN2_3 VSS B1 N_60 VPW NCH W=0.33u L=0.06u
MN2_2 VSS B1 N_62 VPW NCH W=0.33u L=0.06u
MP3_2 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN3_2 Y B0 N_62 VPW NCH W=0.33u L=0.06u
MP2_3 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN3 Y B0 N_64 VPW NCH W=0.33u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN2 N_64 B1 VSS VPW NCH W=0.33u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN0_2 Y C0 VSS VPW NCH W=0.41u L=0.06u
MP1_3 Y C0 P2 VNW PCH W=0.7u L=0.06u
MN0 Y C0 VSS VPW NCH W=0.41u L=0.06u
MP1_2 Y C0 P2 VNW PCH W=0.7u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.7u L=0.06u
MP1_4 Y C0 P2 VNW PCH W=0.7u L=0.06u
.ENDS AOI221X4MA10TR

****
.SUBCKT AOI222X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0 C1
MN5 VSS A1 N_33 VPW NCH W=0.33u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4 Y A0 N_33 VPW NCH W=0.33u L=0.06u
MP5_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4_2 Y A0 N_35 VPW NCH W=0.33u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5_2 N_35 A1 VSS VPW NCH W=0.33u L=0.06u
MN2 VSS B1 N_37 VPW NCH W=0.33u L=0.06u
MP3_2 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN3 Y B0 N_37 VPW NCH W=0.33u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN3_2 Y B0 N_31 VPW NCH W=0.33u L=0.06u
MP2_2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN2_2 N_31 B1 VSS VPW NCH W=0.33u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN1_2 VSS C1 N_42 VPW NCH W=0.33u L=0.06u
MP0_2 Y C1 P2 VNW PCH W=0.7u L=0.06u
MN0_2 Y C0 N_42 VPW NCH W=0.33u L=0.06u
MP1_2 Y C0 P2 VNW PCH W=0.7u L=0.06u
MN0 Y C0 N_40 VPW NCH W=0.33u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.7u L=0.06u
MN1 N_40 C1 VSS VPW NCH W=0.33u L=0.06u
MP0 Y C1 P2 VNW PCH W=0.7u L=0.06u
.ENDS AOI222X2MA10TR

****
.SUBCKT AOI222X3MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0 C1
MP5_3 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4_3 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5 VSS A1 N_45 VPW NCH W=0.495u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4 Y A0 N_45 VPW NCH W=0.495u L=0.06u
MP5_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4_2 Y A0 N_47 VPW NCH W=0.495u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5_2 N_47 A1 VSS VPW NCH W=0.495u L=0.06u
MN2 VSS B1 N_49 VPW NCH W=0.495u L=0.06u
MP3_3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN3 Y B0 N_49 VPW NCH W=0.495u L=0.06u
MP2_3 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN3_2 Y B0 N_43 VPW NCH W=0.495u L=0.06u
MP2_2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN2_2 N_43 B1 VSS VPW NCH W=0.495u L=0.06u
MP3_2 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN1 VSS C1 N_54 VPW NCH W=0.495u L=0.06u
MP0_3 Y C1 P2 VNW PCH W=0.7u L=0.06u
MN0 Y C0 N_54 VPW NCH W=0.495u L=0.06u
MP1_3 Y C0 P2 VNW PCH W=0.7u L=0.06u
MN0_2 Y C0 N_52 VPW NCH W=0.495u L=0.06u
MP1_2 Y C0 P2 VNW PCH W=0.7u L=0.06u
MN1_2 N_52 C1 VSS VPW NCH W=0.495u L=0.06u
MP0_2 Y C1 P2 VNW PCH W=0.7u L=0.06u
MP0 Y C1 P2 VNW PCH W=0.7u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.7u L=0.06u
.ENDS AOI222X3MA10TR

****
.SUBCKT AOI222X4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0 C1
MN5_3 VSS A1 N_57 VPW NCH W=0.33u L=0.06u
MP4_4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4_3 Y A0 N_57 VPW NCH W=0.33u L=0.06u
MP5 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4_4 Y A0 N_59 VPW NCH W=0.33u L=0.06u
MP5_4 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4_3 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5_4 VSS A1 N_59 VPW NCH W=0.33u L=0.06u
MN5 VSS A1 N_61 VPW NCH W=0.33u L=0.06u
MP4_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN4 Y A0 N_61 VPW NCH W=0.33u L=0.06u
MP5_3 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MN4_2 Y A0 N_63 VPW NCH W=0.33u L=0.06u
MP5_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MP4 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MN5_2 N_63 A1 VSS VPW NCH W=0.33u L=0.06u
MN2 VSS B1 N_65 VPW NCH W=0.33u L=0.06u
MP3_2 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN3 Y B0 N_65 VPW NCH W=0.33u L=0.06u
MP2_4 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN3_2 Y B0 N_67 VPW NCH W=0.33u L=0.06u
MP2_3 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MP3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN2_2 VSS B1 N_67 VPW NCH W=0.33u L=0.06u
MN2_3 VSS B1 N_69 VPW NCH W=0.33u L=0.06u
MP3_4 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN3_3 Y B0 N_69 VPW NCH W=0.33u L=0.06u
MP2_2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN3_4 Y B0 N_55 VPW NCH W=0.33u L=0.06u
MP2 P2 B0 P1 VNW PCH W=0.7u L=0.06u
MN2_4 N_55 B1 VSS VPW NCH W=0.33u L=0.06u
MP3_3 P2 B1 P1 VNW PCH W=0.7u L=0.06u
MN1_4 VSS C1 N_74 VPW NCH W=0.33u L=0.06u
MP0_4 Y C1 P2 VNW PCH W=0.7u L=0.06u
MN0_4 Y C0 N_74 VPW NCH W=0.33u L=0.06u
MP1_3 Y C0 P2 VNW PCH W=0.7u L=0.06u
MN0_2 Y C0 N_76 VPW NCH W=0.33u L=0.06u
MP1_2 Y C0 P2 VNW PCH W=0.7u L=0.06u
MP0_3 Y C1 P2 VNW PCH W=0.7u L=0.06u
MN1_2 VSS C1 N_76 VPW NCH W=0.33u L=0.06u
MN1 VSS C1 N_78 VPW NCH W=0.33u L=0.06u
MP0_2 Y C1 P2 VNW PCH W=0.7u L=0.06u
MN0 Y C0 N_78 VPW NCH W=0.33u L=0.06u
MP1 Y C0 P2 VNW PCH W=0.7u L=0.06u
MN0_3 Y C0 N_72 VPW NCH W=0.33u L=0.06u
MP1_4 Y C0 P2 VNW PCH W=0.7u L=0.06u
MN1_3 N_72 C1 VSS VPW NCH W=0.33u L=0.06u
MP0 Y C1 P2 VNW PCH W=0.7u L=0.06u
.ENDS AOI222X4MA10TR

****
.SUBCKT AOI22X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1
MNB2 VSS A1 N_23 VPW NCH W=0.32u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
MNB1 Y A0 N_23 VPW NCH W=0.32u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MNB1_2 Y A0 N_25 VPW NCH W=0.32u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.49u L=0.06u
MNB2_2 N_25 A1 VSS VPW NCH W=0.32u L=0.06u
MNA2 VSS B1 N_27 VPW NCH W=0.32u L=0.06u
MPA2_2 Y B1 P1 VNW PCH W=0.49u L=0.06u
MNA1 Y B0 N_27 VPW NCH W=0.32u L=0.06u
MPA1_2 Y B0 P1 VNW PCH W=0.49u L=0.06u
MNA1_2 Y B0 N_21 VPW NCH W=0.32u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.49u L=0.06u
MNA2_2 N_21 B1 VSS VPW NCH W=0.32u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.49u L=0.06u
.ENDS AOI22X1P4MA10TR

****
.SUBCKT AOI22X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1
MNB2 VSS A1 N_23 VPW NCH W=0.455u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MNB1 Y A0 N_23 VPW NCH W=0.455u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MNB1_2 Y A0 N_25 VPW NCH W=0.455u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.7u L=0.06u
MNB2_2 N_25 A1 VSS VPW NCH W=0.455u L=0.06u
MNA2 VSS B1 N_27 VPW NCH W=0.455u L=0.06u
MPA2_2 Y B1 P1 VNW PCH W=0.7u L=0.06u
MNA1 Y B0 N_27 VPW NCH W=0.455u L=0.06u
MPA1_2 Y B0 P1 VNW PCH W=0.7u L=0.06u
MNA1_2 Y B0 N_21 VPW NCH W=0.455u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.7u L=0.06u
MNA2_2 N_21 B1 VSS VPW NCH W=0.455u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.7u L=0.06u
.ENDS AOI22X2MA10TR

****
.SUBCKT AOI2XB1X1P4MA10TR VDD VSS VPW VNW Y A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.22u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.295u L=0.06u
MNB2 VSS INT N_23 VPW NCH W=0.32u L=0.06u
MPB2_2 P1 INT VDD VNW PCH W=0.49u L=0.06u
MNB1 Y A0 N_23 VPW NCH W=0.32u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MNB1_2 Y A0 N_25 VPW NCH W=0.32u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.49u L=0.06u
MNB2_2 N_25 INT VSS VPW NCH W=0.32u L=0.06u
MPB2 P1 INT VDD VNW PCH W=0.49u L=0.06u
MNA106_2 Y B0 VSS VPW NCH W=0.2u L=0.06u
MPA108 Y B0 P1 VNW PCH W=0.49u L=0.06u
MNA106 Y B0 VSS VPW NCH W=0.2u L=0.06u
MPA108_2 Y B0 P1 VNW PCH W=0.49u L=0.06u
.ENDS AOI2XB1X1P4MA10TR

****
.SUBCKT AOI2XB1X2MA10TR VDD VSS VPW VNW Y A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.295u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.39u L=0.06u
MNB2 VSS INT N_23 VPW NCH W=0.455u L=0.06u
MPB2_2 P1 INT VDD VNW PCH W=0.7u L=0.06u
MNB1 Y A0 N_23 VPW NCH W=0.455u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MNB1_2 Y A0 N_25 VPW NCH W=0.455u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.7u L=0.06u
MNB2_2 N_25 INT VSS VPW NCH W=0.455u L=0.06u
MPB2 P1 INT VDD VNW PCH W=0.7u L=0.06u
MNA106_2 Y B0 VSS VPW NCH W=0.285u L=0.06u
MPA108 Y B0 P1 VNW PCH W=0.7u L=0.06u
MNA106 Y B0 VSS VPW NCH W=0.285u L=0.06u
MPA108_2 Y B0 P1 VNW PCH W=0.7u L=0.06u
.ENDS AOI2XB1X2MA10TR

****
.SUBCKT AOI32X1P4MA10TR VDD VSS VPW VNW Y A0 A1 A2 B0 B1
MPB3_2 P1 A2 VDD VNW PCH W=0.465u L=0.06u
MNB3 VSS A2 N_27 VPW NCH W=0.405u L=0.06u
MNB2 N_27 A1 N_28 VPW NCH W=0.405u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.465u L=0.06u
MNB1 Y A0 N_28 VPW NCH W=0.405u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.465u L=0.06u
MNB1_2 Y A0 N_30 VPW NCH W=0.405u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.465u L=0.06u
MNB2_2 N_30 A1 N_32 VPW NCH W=0.405u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.465u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=0.465u L=0.06u
MNB3_2 N_32 A2 VSS VPW NCH W=0.405u L=0.06u
MNA2_2 VSS B1 N_33 VPW NCH W=0.305u L=0.06u
MPA2_2 Y B1 P1 VNW PCH W=0.465u L=0.06u
MNA1_2 Y B0 N_33 VPW NCH W=0.305u L=0.06u
MPA1_2 Y B0 P1 VNW PCH W=0.465u L=0.06u
MNA1 Y B0 N_25 VPW NCH W=0.305u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.465u L=0.06u
MNA2 N_25 B1 VSS VPW NCH W=0.305u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.465u L=0.06u
.ENDS AOI32X1P4MA10TR

****
.SUBCKT AOI32X2MA10TR VDD VSS VPW VNW Y A0 A1 A2 B0 B1
MPB3_2 P1 A2 VDD VNW PCH W=0.665u L=0.06u
MNB3 VSS A2 N_27 VPW NCH W=0.58u L=0.06u
MNB2 N_27 A1 N_28 VPW NCH W=0.58u L=0.06u
MPB2_2 P1 A1 VDD VNW PCH W=0.665u L=0.06u
MNB1 Y A0 N_28 VPW NCH W=0.58u L=0.06u
MPB1_2 P1 A0 VDD VNW PCH W=0.665u L=0.06u
MNB1_2 Y A0 N_30 VPW NCH W=0.58u L=0.06u
MPB1 P1 A0 VDD VNW PCH W=0.665u L=0.06u
MNB2_2 N_30 A1 N_32 VPW NCH W=0.58u L=0.06u
MPB2 P1 A1 VDD VNW PCH W=0.665u L=0.06u
MPB3 P1 A2 VDD VNW PCH W=0.665u L=0.06u
MNB3_2 N_32 A2 VSS VPW NCH W=0.58u L=0.06u
MNA2_2 VSS B1 N_33 VPW NCH W=0.435u L=0.06u
MPA2_2 Y B1 P1 VNW PCH W=0.665u L=0.06u
MNA1_2 Y B0 N_33 VPW NCH W=0.435u L=0.06u
MPA1_2 Y B0 P1 VNW PCH W=0.665u L=0.06u
MNA1 Y B0 N_25 VPW NCH W=0.435u L=0.06u
MPA1 Y B0 P1 VNW PCH W=0.665u L=0.06u
MNA2 N_25 B1 VSS VPW NCH W=0.435u L=0.06u
MPA2 Y B1 P1 VNW PCH W=0.665u L=0.06u
.ENDS AOI32X2MA10TR

****
.SUBCKT FRICGX0P5BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 VSS HI N_3 VPW NCH W=0.15u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_3 CK NOUT VPW NCH W=0.15u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.18u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.18u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.35u L=0.06u
.ENDS FRICGX0P5BA10TR

****
.SUBCKT FRICGX0P6BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 VSS HI N_9 VPW NCH W=0.15u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_9 CK NOUT VPW NCH W=0.15u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.18u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.215u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.42u L=0.06u
.ENDS FRICGX0P6BA10TR

****
.SUBCKT FRICGX0P7BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 VSS HI N_9 VPW NCH W=0.15u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_9 CK NOUT VPW NCH W=0.15u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.18u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.255u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.49u L=0.06u
.ENDS FRICGX0P7BA10TR

****
.SUBCKT FRICGX0P8BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 VSS HI N_11 VPW NCH W=0.155u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_11 CK NOUT VPW NCH W=0.155u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.185u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.29u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.56u L=0.06u
.ENDS FRICGX0P8BA10TR

****
.SUBCKT FRICGX11BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.6u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1_2 N_148 HI VSS VPW NCH W=0.465u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0_2 NOUT CK N_148 VPW NCH W=0.465u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN0_4 N_150 CK NOUT VPW NCH W=0.465u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN1_4 VSS HI N_150 VPW NCH W=0.465u L=0.06u
MN1 VSS HI N_152 VPW NCH W=0.465u L=0.06u
MN0 NOUT CK N_152 VPW NCH W=0.465u L=0.06u
MP1_4 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN0_3 N_155 CK NOUT VPW NCH W=0.465u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN1_3 N_155 HI VSS VPW NCH W=0.465u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.23u L=0.06u
MNA1_3 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_10 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1_10 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1_9 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1_9 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1_7 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1_7 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1_5 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1_5 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1_6 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1_6 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1_4 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1_4 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1_8 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.36u L=0.06u
MPA1_8 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX11BA10TR

****
.SUBCKT FRICGX13BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.6u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_160 HI VSS VPW NCH W=0.555u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 NOUT CK N_160 VPW NCH W=0.555u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN0_3 N_162 CK NOUT VPW NCH W=0.555u L=0.06u
MP1_4 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN1_3 VSS HI N_162 VPW NCH W=0.555u L=0.06u
MN1_2 VSS HI N_164 VPW NCH W=0.555u L=0.06u
MN0_2 NOUT CK N_164 VPW NCH W=0.555u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN0_4 N_167 CK NOUT VPW NCH W=0.555u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN1_4 N_167 HI VSS VPW NCH W=0.555u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.27u L=0.06u
MNA1_8 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_11 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_5 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_8 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1_4 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_7 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_5 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1_11 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_4 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1_10 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1_7 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_10 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1_9 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1_6 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_9 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1_3 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1_6 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX13BA10TR

****
.SUBCKT FRICGX16BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.7u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_201 HI VSS VPW NCH W=0.54u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 NOUT CK N_201 VPW NCH W=0.54u L=0.06u
MP1_5 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN0_4 N_203 CK NOUT VPW NCH W=0.54u L=0.06u
MP1_4 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN1_4 VSS HI N_203 VPW NCH W=0.54u L=0.06u
MN1_5 VSS HI N_205 VPW NCH W=0.54u L=0.06u
MN0_5 NOUT CK N_205 VPW NCH W=0.54u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN0_3 N_207 CK NOUT VPW NCH W=0.54u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN1_3 VSS HI N_207 VPW NCH W=0.54u L=0.06u
MN1_2 VSS HI N_199 VPW NCH W=0.54u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.33u L=0.06u
MN0_2 N_199 CK NOUT VPW NCH W=0.54u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MPA1_11 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_8 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1_8 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_5 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1_5 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1_4 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1_13 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1_11 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1_14 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1_10 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1_13 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1_7 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1_10 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1_4 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1_7 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1_3 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1_6 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1_12 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1_9 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1_12 ECK NOUT VDD VNW PCH W=0.75u L=0.06u
MNA1_6 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1_9 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX16BA10TR

****
.SUBCKT FRICGX1BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 VSS HI N_11 VPW NCH W=0.18u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_11 CK NOUT VPW NCH W=0.18u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.22u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.36u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX1BA10TR

****
.SUBCKT FRICGX1P2BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN1 N_17 HI VSS VPW NCH W=0.235u L=0.06u
MN0 N_17 CK NOUT VPW NCH W=0.235u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.29u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.215u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.42u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.215u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.42u L=0.06u
.ENDS FRICGX1P2BA10TR

****
.SUBCKT FRICGX1P4BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_17 HI VSS VPW NCH W=0.26u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_17 CK NOUT VPW NCH W=0.26u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.32u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.255u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.49u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.255u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.49u L=0.06u
.ENDS FRICGX1P4BA10TR

****
.SUBCKT FRICGX1P7BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_17 HI VSS VPW NCH W=0.3u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_17 CK NOUT VPW NCH W=0.3u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.365u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.305u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.595u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.305u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.595u L=0.06u
.ENDS FRICGX1P7BA10TR

****
.SUBCKT FRICGX2BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_18 HI VSS VPW NCH W=0.34u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_18 CK NOUT VPW NCH W=0.34u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.41u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.36u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.36u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX2BA10TR

****
.SUBCKT FRICGX2P5BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_19 HI VSS VPW NCH W=0.455u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_19 CK NOUT VPW NCH W=0.455u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.55u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.58u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.58u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.58u L=0.06u
.ENDS FRICGX2P5BA10TR

****
.SUBCKT FRICGX3BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.15u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_16 HI VSS VPW NCH W=0.52u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MN0 N_16 CK NOUT VPW NCH W=0.52u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.63u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.54u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.54u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX3BA10TR

****
.SUBCKT FRICGX3P5BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.3u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1_2 N_26 HI VSS VPW NCH W=0.305u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MN0_2 NOUT CK N_26 VPW NCH W=0.305u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.375u L=0.06u
MN0 N_24 CK NOUT VPW NCH W=0.305u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.375u L=0.06u
MN1 VSS HI N_24 VPW NCH W=0.305u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.42u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.42u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
MNA1_3 ECK NOUT VSS VPW NCH W=0.42u L=0.06u
MPA1_4 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
.ENDS FRICGX3P5BA10TR

****
.SUBCKT FRICGX4BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.3u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_25 HI VSS VPW NCH W=0.34u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MN0 NOUT CK N_25 VPW NCH W=0.34u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.41u L=0.06u
MN0_2 N_23 CK NOUT VPW NCH W=0.34u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.41u L=0.06u
MN1_2 VSS HI N_23 VPW NCH W=0.34u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.48u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.48u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_3 ECK NOUT VSS VPW NCH W=0.48u L=0.06u
MPA1_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX4BA10TR

****
.SUBCKT FRICGX5BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.3u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_32 HI VSS VPW NCH W=0.43u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MN0 NOUT CK N_32 VPW NCH W=0.43u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN0_2 N_30 CK NOUT VPW NCH W=0.43u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN1_2 VSS HI N_30 VPW NCH W=0.43u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_3 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_4 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_5 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX5BA10TR

****
.SUBCKT FRICGX6BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.3u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_35 HI VSS VPW NCH W=0.51u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.15u L=0.06u
MN0 NOUT CK N_35 VPW NCH W=0.51u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.615u L=0.06u
MN0_2 N_33 CK NOUT VPW NCH W=0.51u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.615u L=0.06u
MN1_2 VSS HI N_33 VPW NCH W=0.51u L=0.06u
MPA1_5 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_3 ECK NOUT VSS VPW NCH W=0.435u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.435u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_5 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MPA1_6 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_4 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MPA1_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX6BA10TR

****
.SUBCKT FRICGX7P5BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.45u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1_2 N_116 HI VSS VPW NCH W=0.43u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0_2 NOUT CK N_116 VPW NCH W=0.43u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN0 N_118 CK NOUT VPW NCH W=0.43u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN1 VSS HI N_118 VPW NCH W=0.43u L=0.06u
MN1_3 VSS HI N_114 VPW NCH W=0.43u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.16u L=0.06u
MN0_3 N_114 CK NOUT VPW NCH W=0.43u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_6 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1_5 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_4 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1_3 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_7 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1_6 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_5 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1_4 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.69u L=0.06u
.ENDS FRICGX7P5BA10TR

****
.SUBCKT FRICGX9BA10TR VDD VSS VPW VNW ECK CK
MP4 HI LO VDD VNW PCH W=0.45u L=0.06u
MN4 LO HI VSS VPW NCH W=0.15u L=0.06u
MN1 N_133 HI VSS VPW NCH W=0.515u L=0.06u
MP5 HI HI VDD VNW PCH W=0.15u L=0.06u
MN0 NOUT CK N_133 VPW NCH W=0.515u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.62u L=0.06u
MN0_3 N_135 CK NOUT VPW NCH W=0.515u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.62u L=0.06u
MN1_3 VSS HI N_135 VPW NCH W=0.515u L=0.06u
MN1_2 VSS HI N_131 VPW NCH W=0.515u L=0.06u
MP0 NOUT HI VDD VNW PCH W=0.19u L=0.06u
MN0_2 N_131 CK NOUT VPW NCH W=0.515u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.62u L=0.06u
MNA1_8 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1_8 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1_5 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1_5 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1_7 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1_7 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1_4 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1_4 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1_2 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1_2 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1_6 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1_6 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1_3 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS FRICGX9BA10TR

****
.SUBCKT LATNSPQX3MA10TR VDD VSS VPW VNW Q GN D S
MPA1015 NCLK_ GN VDD VNW PCH W=0.2u L=0.06u
MNA1013 NCLK_ GN VSS VPW NCH W=0.15u L=0.06u
MP4 VDD S N_7 VNW PCH W=0.7u L=0.06u
MN0_2 NIN D VSS VPW NCH W=0.29u L=0.06u
MP0 NIN D N_7 VNW PCH W=0.7u L=0.06u
MP0_2 NIN D N_5 VNW PCH W=0.7u L=0.06u
MN0 NIN D VSS VPW NCH W=0.29u L=0.06u
MP4_2 N_5 S VDD VNW PCH W=0.7u L=0.06u
MNOE NM NCLK_ NIN VPW NCH W=0.58u L=0.06u
MN2 NM GN N_33 VPW NCH W=0.15u L=0.06u
MPOEN NM GN NIN VNW PCH W=0.58u L=0.06u
MP3 N_17 NCLK_ NM VNW PCH W=0.2u L=0.06u
MN3 VSS M N_33 VPW NCH W=0.15u L=0.06u
MP2 N_17 M N_14 VNW PCH W=0.2u L=0.06u
MN5 NM S VSS VPW NCH W=0.2u L=0.06u
MP5 N_14 S VDD VNW PCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.58u L=0.06u
MPA1019_3 Q NM VDD VNW PCH W=0.7u L=0.06u
MNA1017_3 Q NM VSS VPW NCH W=0.58u L=0.06u
MPA1019_2 Q NM VDD VNW PCH W=0.7u L=0.06u
MNA1017_2 Q NM VSS VPW NCH W=0.58u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.7u L=0.06u
.ENDS LATNSPQX3MA10TR

****
.SUBCKT LATSPQX3MA10TR VDD VSS VPW VNW Q G D S
MPA1015 NCLK G VDD VNW PCH W=0.23u L=0.06u
MNA1013 NCLK G VSS VPW NCH W=0.18u L=0.06u
MP4 VDD S N_7 VNW PCH W=0.7u L=0.06u
MN0 NIN D VSS VPW NCH W=0.29u L=0.06u
MP0 NIN D N_7 VNW PCH W=0.7u L=0.06u
MP0_2 NIN D N_5 VNW PCH W=0.7u L=0.06u
MN0_2 NIN D VSS VPW NCH W=0.29u L=0.06u
MP4_2 N_5 S VDD VNW PCH W=0.7u L=0.06u
MNOE NM G NIN VPW NCH W=0.58u L=0.06u
MN2 NM NCLK N_33 VPW NCH W=0.15u L=0.06u
MPOEN NM NCLK NIN VNW PCH W=0.58u L=0.06u
MP3 N_17 G NM VNW PCH W=0.2u L=0.06u
MN3 VSS M N_33 VPW NCH W=0.15u L=0.06u
MP2 N_17 M N_14 VNW PCH W=0.2u L=0.06u
MN5 NM S VSS VPW NCH W=0.2u L=0.06u
MP5 N_14 S VDD VNW PCH W=0.2u L=0.06u
MNA1 M NM VSS VPW NCH W=0.15u L=0.06u
MPA1 M NM VDD VNW PCH W=0.15u L=0.06u
MNA1017 Q NM VSS VPW NCH W=0.58u L=0.06u
MPA1019_3 Q NM VDD VNW PCH W=0.7u L=0.06u
MNA1017_3 Q NM VSS VPW NCH W=0.58u L=0.06u
MPA1019_2 Q NM VDD VNW PCH W=0.7u L=0.06u
MNA1017_2 Q NM VSS VPW NCH W=0.58u L=0.06u
MPA1019 Q NM VDD VNW PCH W=0.7u L=0.06u
.ENDS LATSPQX3MA10TR

****
.SUBCKT MX2X1P4BA10TR VDD VSS VPW VNW Y A B S0
MNA1016 INT0 A N_34 VPW NCH W=0.355u L=0.06u
MPA1020 INT0 A VDD VNW PCH W=0.43u L=0.06u
MNA2018 N_34 NSEL VSS VPW NCH W=0.355u L=0.06u
MPA2022 INT0 NSEL VDD VNW PCH W=0.43u L=0.06u
MNA1 NSEL S0 VSS VPW NCH W=0.45u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.595u L=0.06u
MNA2010 VSS S0 N_29 VPW NCH W=0.355u L=0.06u
MPA2014 INT1 S0 VDD VNW PCH W=0.43u L=0.06u
MNA108 INT1 B N_29 VPW NCH W=0.355u L=0.06u
MPA1012 INT1 B VDD VNW PCH W=0.43u L=0.06u
MNA2_2 N_26 INT1 VSS VPW NCH W=0.405u L=0.06u
MPA2_2 Y INT1 VDD VNW PCH W=0.49u L=0.06u
MNA102_2 Y INT0 N_26 VPW NCH W=0.405u L=0.06u
MPA105_2 Y INT0 VDD VNW PCH W=0.49u L=0.06u
MNA102 Y INT0 N_24 VPW NCH W=0.405u L=0.06u
MPA105 Y INT0 VDD VNW PCH W=0.49u L=0.06u
MNA2 N_24 INT1 VSS VPW NCH W=0.405u L=0.06u
MPA2 Y INT1 VDD VNW PCH W=0.49u L=0.06u
.ENDS MX2X1P4BA10TR

****
.SUBCKT MX2X1P4MA10TR VDD VSS VPW VNW Y A B S0
MPA1 NSEL S0 VDD VNW PCH W=0.7u L=0.06u
MNA1 NSEL S0 VSS VPW NCH W=0.53u L=0.06u
MNB2_2 N_30 S0 VSS VPW NCH W=0.28u L=0.06u
MPB2 P1 S0 VDD VNW PCH W=0.42u L=0.06u
MNB1_2 INT B N_30 VPW NCH W=0.28u L=0.06u
MPB1_2 P1 B VDD VNW PCH W=0.42u L=0.06u
MNB1 INT B N_32 VPW NCH W=0.28u L=0.06u
MPB1 P1 B VDD VNW PCH W=0.42u L=0.06u
MPB2_2 P1 S0 VDD VNW PCH W=0.42u L=0.06u
MNB2 N_32 S0 VSS VPW NCH W=0.28u L=0.06u
MNA2 VSS NSEL N_34 VPW NCH W=0.28u L=0.06u
MPA2_2 INT NSEL P1 VNW PCH W=0.42u L=0.06u
MNA1010 INT A N_34 VPW NCH W=0.28u L=0.06u
MPA1013_2 INT A P1 VNW PCH W=0.42u L=0.06u
MNA1010_2 INT A N_28 VPW NCH W=0.28u L=0.06u
MPA1013 INT A P1 VNW PCH W=0.42u L=0.06u
MNA2_2 N_28 NSEL VSS VPW NCH W=0.28u L=0.06u
MPA2 INT NSEL P1 VNW PCH W=0.42u L=0.06u
MNA102_2 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA104_2 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA102 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA104 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS MX2X1P4MA10TR

****
.SUBCKT MX2X2BA10TR VDD VSS VPW VNW Y A B S0
MNA1016 INT0 A N_30 VPW NCH W=0.47u L=0.06u
MPA1020 INT0 A VDD VNW PCH W=0.575u L=0.06u
MNA2018 N_30 NSEL VSS VPW NCH W=0.47u L=0.06u
MPA2022 INT0 NSEL VDD VNW PCH W=0.575u L=0.06u
MNA1 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.665u L=0.06u
MNA2010 VSS S0 N_25 VPW NCH W=0.47u L=0.06u
MPA2014 INT1 S0 VDD VNW PCH W=0.575u L=0.06u
MNA108 INT1 B N_25 VPW NCH W=0.47u L=0.06u
MPA1012 INT1 B VDD VNW PCH W=0.575u L=0.06u
MNA2_2 VSS INT1 N_34 VPW NCH W=0.58u L=0.06u
MPA2_2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_2 Y INT0 N_34 VPW NCH W=0.58u L=0.06u
MPA105_2 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102 Y INT0 N_32 VPW NCH W=0.58u L=0.06u
MPA105 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA2 N_32 INT1 VSS VPW NCH W=0.58u L=0.06u
MPA2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
.ENDS MX2X2BA10TR

****
.SUBCKT MX2X2MA10TR VDD VSS VPW VNW Y A B S0
MNA1 NSEL S0 VSS VPW NCH W=0.33u L=0.06u
MPA1_2 NSEL S0 VDD VNW PCH W=0.435u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.435u L=0.06u
MNA1_2 NSEL S0 VSS VPW NCH W=0.33u L=0.06u
MNB2 VSS S0 N_32 VPW NCH W=0.38u L=0.06u
MPB2_2 P1 S0 VDD VNW PCH W=0.575u L=0.06u
MNB1 INT B N_32 VPW NCH W=0.38u L=0.06u
MPB1_2 P1 B VDD VNW PCH W=0.575u L=0.06u
MNB1_2 INT B N_34 VPW NCH W=0.38u L=0.06u
MPB1 P1 B VDD VNW PCH W=0.575u L=0.06u
MPB2 P1 S0 VDD VNW PCH W=0.575u L=0.06u
MNB2_2 N_34 S0 VSS VPW NCH W=0.38u L=0.06u
MNA2_2 VSS NSEL N_36 VPW NCH W=0.38u L=0.06u
MPA2_2 INT NSEL P1 VNW PCH W=0.575u L=0.06u
MNA1010_2 INT A N_36 VPW NCH W=0.38u L=0.06u
MPA1013_2 INT A P1 VNW PCH W=0.575u L=0.06u
MNA1010 INT A N_30 VPW NCH W=0.38u L=0.06u
MPA1013 INT A P1 VNW PCH W=0.575u L=0.06u
MNA2 N_30 NSEL VSS VPW NCH W=0.38u L=0.06u
MPA2 INT NSEL P1 VNW PCH W=0.575u L=0.06u
MNA102_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA104_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA102 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA104 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS MX2X2MA10TR

****
.SUBCKT MX2X3BA10TR VDD VSS VPW VNW Y A B S0
MNA2018 VSS NSEL N_37 VPW NCH W=0.36u L=0.06u
MPA2022_2 INT0 NSEL VDD VNW PCH W=0.44u L=0.06u
MNA1016 INT0 A N_37 VPW NCH W=0.36u L=0.06u
MPA1020_2 INT0 A VDD VNW PCH W=0.44u L=0.06u
MNA1016_2 INT0 A N_39 VPW NCH W=0.36u L=0.06u
MPA1020 INT0 A VDD VNW PCH W=0.44u L=0.06u
MNA2018_2 N_39 NSEL VSS VPW NCH W=0.36u L=0.06u
MPA2022 INT0 NSEL VDD VNW PCH W=0.44u L=0.06u
MNA1 NSEL S0 VSS VPW NCH W=0.4u L=0.06u
MPA1_2 NSEL S0 VDD VNW PCH W=0.525u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.525u L=0.06u
MNA1_2 NSEL S0 VSS VPW NCH W=0.4u L=0.06u
MNA2010 N_43 S0 VSS VPW NCH W=0.36u L=0.06u
MPA2014_2 INT1 S0 VDD VNW PCH W=0.44u L=0.06u
MNA108 INT1 B N_43 VPW NCH W=0.36u L=0.06u
MPA1012_2 INT1 B VDD VNW PCH W=0.44u L=0.06u
MNA108_2 INT1 B N_45 VPW NCH W=0.36u L=0.06u
MPA1012 INT1 B VDD VNW PCH W=0.44u L=0.06u
MPA2014 INT1 S0 VDD VNW PCH W=0.44u L=0.06u
MNA2010_2 N_45 S0 VSS VPW NCH W=0.36u L=0.06u
MNA2_2 VSS INT1 N_47 VPW NCH W=0.58u L=0.06u
MPA2_3 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_2 Y INT0 N_47 VPW NCH W=0.58u L=0.06u
MPA105_3 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102_3 Y INT0 N_49 VPW NCH W=0.58u L=0.06u
MPA105_2 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA2_3 VSS INT1 N_49 VPW NCH W=0.58u L=0.06u
MPA2_2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA2 VSS INT1 N_35 VPW NCH W=0.58u L=0.06u
MPA2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102 N_35 INT0 Y VPW NCH W=0.58u L=0.06u
MPA105 Y INT0 VDD VNW PCH W=0.7u L=0.06u
.ENDS MX2X3BA10TR

****
.SUBCKT MX2X4BA10TR VDD VSS VPW VNW Y A B S0
MNA2018 VSS NSEL N_43 VPW NCH W=0.47u L=0.06u
MPA2022_2 INT0 NSEL VDD VNW PCH W=0.575u L=0.06u
MNA1016 INT0 A N_43 VPW NCH W=0.47u L=0.06u
MPA1020_2 INT0 A VDD VNW PCH W=0.575u L=0.06u
MNA1016_2 INT0 A N_45 VPW NCH W=0.47u L=0.06u
MPA1020 INT0 A VDD VNW PCH W=0.575u L=0.06u
MNA2018_2 N_45 NSEL VSS VPW NCH W=0.47u L=0.06u
MPA2022 INT0 NSEL VDD VNW PCH W=0.575u L=0.06u
MNA1 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MPA1_2 NSEL S0 VDD VNW PCH W=0.665u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.665u L=0.06u
MNA1_2 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MNA2010 N_49 S0 VSS VPW NCH W=0.47u L=0.06u
MPA2014_2 INT1 S0 VDD VNW PCH W=0.575u L=0.06u
MNA108 INT1 B N_49 VPW NCH W=0.47u L=0.06u
MPA1012_2 INT1 B VDD VNW PCH W=0.575u L=0.06u
MNA108_2 INT1 B N_51 VPW NCH W=0.47u L=0.06u
MPA1012 INT1 B VDD VNW PCH W=0.575u L=0.06u
MPA2014 INT1 S0 VDD VNW PCH W=0.575u L=0.06u
MNA2010_2 N_51 S0 VSS VPW NCH W=0.47u L=0.06u
MNA2_2 VSS INT1 N_53 VPW NCH W=0.58u L=0.06u
MPA2_4 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_2 Y INT0 N_53 VPW NCH W=0.58u L=0.06u
MPA105_4 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102_3 Y INT0 N_55 VPW NCH W=0.58u L=0.06u
MPA105_2 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MPA2_3 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA2_3 VSS INT1 N_55 VPW NCH W=0.58u L=0.06u
MNA2_4 VSS INT1 N_57 VPW NCH W=0.58u L=0.06u
MPA2_2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_4 Y INT0 N_57 VPW NCH W=0.58u L=0.06u
MPA105_3 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102 Y INT0 N_41 VPW NCH W=0.58u L=0.06u
MPA105 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA2 N_41 INT1 VSS VPW NCH W=0.58u L=0.06u
MPA2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
.ENDS MX2X4BA10TR

****
.SUBCKT MX2X6BA10TR VDD VSS VPW VNW Y A B S0
MNA2018 VSS NSEL N_63 VPW NCH W=0.47u L=0.06u
MPA2022 INT0 NSEL VDD VNW PCH W=0.57u L=0.06u
MNA1016 INT0 A N_63 VPW NCH W=0.47u L=0.06u
MPA1020_2 INT0 A VDD VNW PCH W=0.57u L=0.06u
MNA1016_2 INT0 A N_65 VPW NCH W=0.47u L=0.06u
MPA1020 INT0 A VDD VNW PCH W=0.57u L=0.06u
MNA2018_2 VSS NSEL N_65 VPW NCH W=0.47u L=0.06u
MPA2022_3 INT0 NSEL VDD VNW PCH W=0.57u L=0.06u
MNA2018_3 VSS NSEL N_61 VPW NCH W=0.47u L=0.06u
MPA2022_2 INT0 NSEL VDD VNW PCH W=0.57u L=0.06u
MNA1016_3 N_61 A INT0 VPW NCH W=0.47u L=0.06u
MPA1020_3 INT0 A VDD VNW PCH W=0.57u L=0.06u
MNA1_3 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MPA1_3 NSEL S0 VDD VNW PCH W=0.67u L=0.06u
MNA1_2 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MPA1_2 NSEL S0 VDD VNW PCH W=0.67u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.67u L=0.06u
MNA1 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MPA2014_3 INT1 S0 VDD VNW PCH W=0.57u L=0.06u
MNA2010 N_73 S0 VSS VPW NCH W=0.47u L=0.06u
MPA1012_2 INT1 B VDD VNW PCH W=0.57u L=0.06u
MNA108 INT1 B N_73 VPW NCH W=0.47u L=0.06u
MNA108_3 INT1 B N_75 VPW NCH W=0.47u L=0.06u
MPA1012 INT1 B VDD VNW PCH W=0.57u L=0.06u
MNA2010_3 VSS S0 N_75 VPW NCH W=0.47u L=0.06u
MPA2014_2 INT1 S0 VDD VNW PCH W=0.57u L=0.06u
MNA2010_2 VSS S0 N_68 VPW NCH W=0.47u L=0.06u
MPA2014 INT1 S0 VDD VNW PCH W=0.57u L=0.06u
MNA108_2 N_68 B INT1 VPW NCH W=0.47u L=0.06u
MPA1012_3 INT1 B VDD VNW PCH W=0.57u L=0.06u
MNA2_3 VSS INT1 N_80 VPW NCH W=0.58u L=0.06u
MPA2_4 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_3 Y INT0 N_80 VPW NCH W=0.58u L=0.06u
MPA105_6 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102 Y INT0 N_82 VPW NCH W=0.58u L=0.06u
MPA105_5 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MPA2_2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA2 VSS INT1 N_82 VPW NCH W=0.58u L=0.06u
MNA2_6 VSS INT1 N_84 VPW NCH W=0.58u L=0.06u
MPA2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_6 Y INT0 N_84 VPW NCH W=0.58u L=0.06u
MPA105_4 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102_5 Y INT0 N_86 VPW NCH W=0.58u L=0.06u
MPA105_3 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MPA2_5 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA2_5 N_86 INT1 VSS VPW NCH W=0.58u L=0.06u
MNA2_2 VSS INT1 N_88 VPW NCH W=0.58u L=0.06u
MPA2_6 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_2 Y INT0 N_88 VPW NCH W=0.58u L=0.06u
MPA105_2 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102_4 Y INT0 N_78 VPW NCH W=0.58u L=0.06u
MPA105 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA2_4 N_78 INT1 VSS VPW NCH W=0.58u L=0.06u
MPA2_3 Y INT1 VDD VNW PCH W=0.7u L=0.06u
.ENDS MX2X6BA10TR

****
.SUBCKT MX2X8BA10TR VDD VSS VPW VNW Y A B S0
MNA2018_3 VSS NSEL N_40 VPW NCH W=0.47u L=0.06u
MPA2022 INT0 NSEL VDD VNW PCH W=0.57u L=0.06u
MNA1016_3 INT0 A N_40 VPW NCH W=0.47u L=0.06u
MPA1020_2 INT0 A VDD VNW PCH W=0.57u L=0.06u
MNA1016 INT0 A N_42 VPW NCH W=0.47u L=0.06u
MPA1020 INT0 A VDD VNW PCH W=0.57u L=0.06u
MNA2018 VSS NSEL N_42 VPW NCH W=0.47u L=0.06u
MPA2022_4 INT0 NSEL VDD VNW PCH W=0.57u L=0.06u
MNA2018_2 VSS NSEL N_44 VPW NCH W=0.47u L=0.06u
MPA2022_3 INT0 NSEL VDD VNW PCH W=0.57u L=0.06u
MNA1016_2 INT0 A N_44 VPW NCH W=0.47u L=0.06u
MPA1020_4 INT0 A VDD VNW PCH W=0.57u L=0.06u
MNA1016_4 N_46 A INT0 VPW NCH W=0.47u L=0.06u
MPA1020_3 INT0 A VDD VNW PCH W=0.57u L=0.06u
MNA2018_4 VSS NSEL N_46 VPW NCH W=0.47u L=0.06u
MPA2022_2 INT0 NSEL VDD VNW PCH W=0.57u L=0.06u
MNA1_4 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MPA1_4 NSEL S0 VDD VNW PCH W=0.665u L=0.06u
MNA1_3 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MPA1_3 NSEL S0 VDD VNW PCH W=0.665u L=0.06u
MNA1_2 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MPA1_2 NSEL S0 VDD VNW PCH W=0.665u L=0.06u
MPA1 NSEL S0 VDD VNW PCH W=0.665u L=0.06u
MNA1 NSEL S0 VSS VPW NCH W=0.505u L=0.06u
MPA2014_2 INT1 S0 VDD VNW PCH W=0.57u L=0.06u
MNA2010_3 N_52 S0 VSS VPW NCH W=0.47u L=0.06u
MPA1012_2 INT1 B VDD VNW PCH W=0.57u L=0.06u
MNA108_3 INT1 B N_52 VPW NCH W=0.47u L=0.06u
MNA108_4 INT1 B N_54 VPW NCH W=0.47u L=0.06u
MPA1012 INT1 B VDD VNW PCH W=0.57u L=0.06u
MNA2010_4 VSS S0 N_54 VPW NCH W=0.47u L=0.06u
MPA2014_4 INT1 S0 VDD VNW PCH W=0.57u L=0.06u
MNA2010 VSS S0 N_56 VPW NCH W=0.47u L=0.06u
MPA2014_3 INT1 S0 VDD VNW PCH W=0.57u L=0.06u
MNA108 INT1 B N_56 VPW NCH W=0.47u L=0.06u
MPA1012_4 INT1 B VDD VNW PCH W=0.57u L=0.06u
MNA108_2 INT1 B N_58 VPW NCH W=0.47u L=0.06u
MPA1012_3 INT1 B VDD VNW PCH W=0.57u L=0.06u
MNA2010_2 N_58 S0 VSS VPW NCH W=0.47u L=0.06u
MPA2014 INT1 S0 VDD VNW PCH W=0.57u L=0.06u
MNA2_5 VSS INT1 N_61 VPW NCH W=0.58u L=0.06u
MPA2_8 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_5 Y INT0 N_61 VPW NCH W=0.58u L=0.06u
MPA105_6 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102_7 N_63 INT0 Y VPW NCH W=0.58u L=0.06u
MPA105_4 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MPA2_7 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA2_7 VSS INT1 N_63 VPW NCH W=0.58u L=0.06u
MNA2_3 VSS INT1 N_65 VPW NCH W=0.58u L=0.06u
MPA2_5 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_3 Y INT0 N_65 VPW NCH W=0.58u L=0.06u
MPA105_2 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102 Y INT0 N_67 VPW NCH W=0.58u L=0.06u
MPA105_8 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MPA2_3 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA2 VSS INT1 N_67 VPW NCH W=0.58u L=0.06u
MNA2_6 N_69 INT1 VSS VPW NCH W=0.58u L=0.06u
MPA2_2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_6 Y INT0 N_69 VPW NCH W=0.58u L=0.06u
MPA105_5 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102_8 Y INT0 N_73 VPW NCH W=0.58u L=0.06u
MPA105_3 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MPA2_6 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA2_8 VSS INT1 N_73 VPW NCH W=0.58u L=0.06u
MNA2_4 VSS INT1 N_75 VPW NCH W=0.58u L=0.06u
MPA2_4 Y INT1 VDD VNW PCH W=0.7u L=0.06u
MNA102_4 Y INT0 N_75 VPW NCH W=0.58u L=0.06u
MPA105 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA102_2 Y INT0 N_72 VPW NCH W=0.58u L=0.06u
MPA105_7 Y INT0 VDD VNW PCH W=0.7u L=0.06u
MNA2_2 N_72 INT1 VSS VPW NCH W=0.58u L=0.06u
MPA2 Y INT1 VDD VNW PCH W=0.7u L=0.06u
.ENDS MX2X8BA10TR

****
.SUBCKT NAND2BX1P4MA10TR VDD VSS VPW VNW Y AN B
MPA106 NET24 AN VDD VNW PCH W=0.28u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.21u L=0.06u
MNA2 N_17 B VSS VPW NCH W=0.41u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.34u L=0.06u
MNA1 Y NET24 N_17 VPW NCH W=0.41u L=0.06u
MPA1_2 Y NET24 VDD VNW PCH W=0.34u L=0.06u
MNA1_2 Y NET24 N_15 VPW NCH W=0.41u L=0.06u
MPA1 Y NET24 VDD VNW PCH W=0.34u L=0.06u
MNA2_2 N_15 B VSS VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.34u L=0.06u
.ENDS NAND2BX1P4MA10TR

****
.SUBCKT NAND2BX2MA10TR VDD VSS VPW VNW Y AN B
MPA106 NET24 AN VDD VNW PCH W=0.365u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.275u L=0.06u
MNA2 N_12 B VSS VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1 Y NET24 N_12 VPW NCH W=0.58u L=0.06u
MPA1_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y NET24 N_10 VPW NCH W=0.58u L=0.06u
MPA1 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_2 N_10 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2BX2MA10TR

****
.SUBCKT NAND2BX3MA10TR VDD VSS VPW VNW Y AN B
MPA106 NET24 AN VDD VNW PCH W=0.56u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.425u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_2 VSS B N_22 VPW NCH W=0.58u L=0.06u
MPA1_3 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y NET24 N_22 VPW NCH W=0.58u L=0.06u
MNA1 Y NET24 N_24 VPW NCH W=0.58u L=0.06u
MPA1_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS B N_24 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_3 VSS B N_19 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_3 N_19 NET24 Y VPW NCH W=0.58u L=0.06u
MPA1 Y NET24 VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2BX3MA10TR

****
.SUBCKT NAND2BX4MA10TR VDD VSS VPW VNW Y AN B
MPA106 NET24 AN VDD VNW PCH W=0.7u L=0.06u
MNA104 NET24 AN VSS VPW NCH W=0.53u L=0.06u
MPA2_4 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_4 VSS B N_26 VPW NCH W=0.58u L=0.06u
MPA1_4 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_4 Y NET24 N_26 VPW NCH W=0.58u L=0.06u
MNA1 Y NET24 N_28 VPW NCH W=0.58u L=0.06u
MPA1_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS B N_28 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_3 VSS B N_30 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y NET24 N_30 VPW NCH W=0.58u L=0.06u
MPA1_3 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y NET24 N_23 VPW NCH W=0.58u L=0.06u
MPA1 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_2 N_23 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2BX4MA10TR

****
.SUBCKT NAND2BX6MA10TR VDD VSS VPW VNW Y AN B
MNA104 NET24 AN VSS VPW NCH W=0.415u L=0.06u
MPA106_2 NET24 AN VDD VNW PCH W=0.55u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.55u L=0.06u
MNA104_2 NET24 AN VSS VPW NCH W=0.415u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_2 VSS B N_37 VPW NCH W=0.58u L=0.06u
MPA1_6 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y NET24 N_37 VPW NCH W=0.58u L=0.06u
MNA1_5 Y NET24 N_39 VPW NCH W=0.58u L=0.06u
MPA1_4 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MPA2_4 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_5 VSS B N_39 VPW NCH W=0.58u L=0.06u
MNA2_6 VSS B N_41 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_6 Y NET24 N_41 VPW NCH W=0.58u L=0.06u
MPA1_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1 Y NET24 N_43 VPW NCH W=0.58u L=0.06u
MPA1_5 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MPA2_6 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS B N_43 VPW NCH W=0.58u L=0.06u
MNA2_3 VSS B N_45 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y NET24 N_45 VPW NCH W=0.58u L=0.06u
MPA1_3 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_4 Y NET24 N_33 VPW NCH W=0.58u L=0.06u
MPA1 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_4 N_33 B VSS VPW NCH W=0.58u L=0.06u
MPA2_5 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2BX6MA10TR

****
.SUBCKT NAND2BX8MA10TR VDD VSS VPW VNW Y AN B
MNA104 NET24 AN VSS VPW NCH W=0.53u L=0.06u
MPA106_2 NET24 AN VDD VNW PCH W=0.7u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.7u L=0.06u
MNA104_2 NET24 AN VSS VPW NCH W=0.53u L=0.06u
MPA2_8 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS B N_45 VPW NCH W=0.58u L=0.06u
MPA1_8 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1 Y NET24 N_45 VPW NCH W=0.58u L=0.06u
MNA1_2 Y NET24 N_47 VPW NCH W=0.58u L=0.06u
MPA1_4 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MPA2_7 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_2 VSS B N_47 VPW NCH W=0.58u L=0.06u
MNA2_8 VSS B N_49 VPW NCH W=0.58u L=0.06u
MPA2_4 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_8 Y NET24 N_49 VPW NCH W=0.58u L=0.06u
MPA1_7 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_7 Y NET24 N_51 VPW NCH W=0.58u L=0.06u
MPA1_3 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MPA2_6 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_7 VSS B N_51 VPW NCH W=0.58u L=0.06u
MNA2_6 VSS B N_53 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_6 Y NET24 N_53 VPW NCH W=0.58u L=0.06u
MPA1_6 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_5 Y NET24 N_55 VPW NCH W=0.58u L=0.06u
MPA1_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MPA2_5 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2_5 VSS B N_55 VPW NCH W=0.58u L=0.06u
MNA2_4 VSS B N_57 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1_4 Y NET24 N_57 VPW NCH W=0.58u L=0.06u
MPA1_5 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y NET24 N_41 VPW NCH W=0.58u L=0.06u
MPA1 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_3 N_41 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2BX8MA10TR

****
.SUBCKT NAND2X1P4AA10TR VDD VSS VPW VNW Y A B
MPA2_2 Y B VDD VNW PCH W=0.415u L=0.06u
MNA2 VSS B N_15 VPW NCH W=0.405u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.415u L=0.06u
MNA1 Y A N_15 VPW NCH W=0.405u L=0.06u
MNA1_2 Y A N_13 VPW NCH W=0.405u L=0.06u
MPA1 Y A VDD VNW PCH W=0.415u L=0.06u
MNA2_2 N_13 B VSS VPW NCH W=0.405u L=0.06u
MPA2 Y B VDD VNW PCH W=0.415u L=0.06u
.ENDS NAND2X1P4AA10TR

****
.SUBCKT NAND2X1P4BA10TR VDD VSS VPW VNW Y A B
MPA2_2 Y B VDD VNW PCH W=0.49u L=0.06u
MNA2 VSS B N_15 VPW NCH W=0.405u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.49u L=0.06u
MNA1 Y A N_15 VPW NCH W=0.405u L=0.06u
MNA1_2 Y A N_13 VPW NCH W=0.405u L=0.06u
MPA1 Y A VDD VNW PCH W=0.49u L=0.06u
MNA2_2 N_13 B VSS VPW NCH W=0.405u L=0.06u
MPA2 Y B VDD VNW PCH W=0.49u L=0.06u
.ENDS NAND2X1P4BA10TR

****
.SUBCKT NAND2X1P4MA10TR VDD VSS VPW VNW Y A B
MPA2_2 Y B VDD VNW PCH W=0.34u L=0.06u
MNA2 VSS B N_5 VPW NCH W=0.41u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.34u L=0.06u
MNA1 Y A N_5 VPW NCH W=0.41u L=0.06u
MNA1_2 Y A N_3 VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.34u L=0.06u
MNA2_2 N_3 B VSS VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.34u L=0.06u
.ENDS NAND2X1P4MA10TR

****
.SUBCKT NAND2X2AA10TR VDD VSS VPW VNW Y A B
MPA2_2 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2 VSS B N_15 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1 Y A N_15 VPW NCH W=0.58u L=0.06u
MNA1_2 Y A N_13 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.59u L=0.06u
MNA2_2 N_13 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.59u L=0.06u
.ENDS NAND2X2AA10TR

****
.SUBCKT NAND2X2BA10TR VDD VSS VPW VNW Y A B
MNA2 VSS B N_15 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.7u L=0.06u
MNA1 Y A N_15 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y A N_13 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.7u L=0.06u
MNA2_2 N_13 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.7u L=0.06u
.ENDS NAND2X2BA10TR

****
.SUBCKT NAND2X2MA10TR VDD VSS VPW VNW Y A B
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS B N_15 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1 Y A N_15 VPW NCH W=0.58u L=0.06u
MNA1_2 Y A N_13 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_2 N_13 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2X2MA10TR

****
.SUBCKT NAND2X3AA10TR VDD VSS VPW VNW Y A B
MPA2_3 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2 VSS B N_19 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1 Y A N_19 VPW NCH W=0.58u L=0.06u
MNA1_3 Y A N_21 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.59u L=0.06u
MNA2_3 VSS B N_21 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2_2 VSS B N_17 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.59u L=0.06u
MNA1_2 N_17 A Y VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.59u L=0.06u
.ENDS NAND2X3AA10TR

****
.SUBCKT NAND2X3BA10TR VDD VSS VPW VNW Y A B
MNA2 VSS B N_19 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.7u L=0.06u
MNA1 Y A N_19 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1_3 Y A N_21 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.7u L=0.06u
MNA2_3 VSS B N_21 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2_2 VSS B N_17 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 N_17 A Y VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.7u L=0.06u
.ENDS NAND2X3BA10TR

****
.SUBCKT NAND2X4AA10TR VDD VSS VPW VNW Y A B
MPA2_4 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2 VSS B N_23 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1 Y A N_23 VPW NCH W=0.58u L=0.06u
MNA1_3 Y A N_25 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.59u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2_3 VSS B N_25 VPW NCH W=0.58u L=0.06u
MNA2_2 VSS B N_27 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.59u L=0.06u
MNA1_2 Y A N_27 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1_4 Y A N_21 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.59u L=0.06u
MNA2_4 N_21 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.59u L=0.06u
.ENDS NAND2X4AA10TR

****
.SUBCKT NAND2X4BA10TR VDD VSS VPW VNW Y A B
MPA2_4 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2 VSS B N_23 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1 Y A N_23 VPW NCH W=0.58u L=0.06u
MNA1_3 Y A N_25 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.7u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2_3 VSS B N_25 VPW NCH W=0.58u L=0.06u
MNA2_2 VSS B N_27 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y A N_27 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1_4 Y A N_21 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.7u L=0.06u
MNA2_4 N_21 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.7u L=0.06u
.ENDS NAND2X4BA10TR

****
.SUBCKT NAND2X6AA10TR VDD VSS VPW VNW Y A B
MPA2_2 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2_5 VSS B N_31 VPW NCH W=0.58u L=0.06u
MPA1_6 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1_5 Y A N_31 VPW NCH W=0.58u L=0.06u
MNA1_6 Y A N_33 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.59u L=0.06u
MPA2_4 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2_6 VSS B N_33 VPW NCH W=0.58u L=0.06u
MNA2 VSS B N_35 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.59u L=0.06u
MNA1 Y A N_35 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1_3 Y A N_37 VPW NCH W=0.58u L=0.06u
MPA1_5 Y A VDD VNW PCH W=0.59u L=0.06u
MPA2_6 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2_3 VSS B N_37 VPW NCH W=0.58u L=0.06u
MNA2_4 VSS B N_39 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.59u L=0.06u
MNA1_4 Y A N_39 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1_2 Y A N_29 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.59u L=0.06u
MNA2_2 N_29 B VSS VPW NCH W=0.58u L=0.06u
MPA2_5 Y B VDD VNW PCH W=0.59u L=0.06u
.ENDS NAND2X6AA10TR

****
.SUBCKT NAND2X6BA10TR VDD VSS VPW VNW Y A B
MPA2_2 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2_5 VSS B N_18 VPW NCH W=0.58u L=0.06u
MPA1_6 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1_5 Y A N_18 VPW NCH W=0.58u L=0.06u
MNA1_6 Y A N_20 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.7u L=0.06u
MPA2_4 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2_6 VSS B N_20 VPW NCH W=0.58u L=0.06u
MNA2 VSS B N_22 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.7u L=0.06u
MNA1 Y A N_22 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1_3 Y A N_24 VPW NCH W=0.58u L=0.06u
MPA1_5 Y A VDD VNW PCH W=0.7u L=0.06u
MPA2_6 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2_3 VSS B N_24 VPW NCH W=0.58u L=0.06u
MNA2_4 VSS B N_26 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.7u L=0.06u
MNA1_4 Y A N_26 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y A N_16 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.7u L=0.06u
MNA2_2 N_16 B VSS VPW NCH W=0.58u L=0.06u
MPA2_5 Y B VDD VNW PCH W=0.7u L=0.06u
.ENDS NAND2X6BA10TR

****
.SUBCKT NAND2X8AA10TR VDD VSS VPW VNW Y A B
MPA2_8 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2 VSS B N_22 VPW NCH W=0.58u L=0.06u
MPA1_8 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1 Y A N_22 VPW NCH W=0.58u L=0.06u
MNA1_8 Y A N_24 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.59u L=0.06u
MPA2_7 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2_8 VSS B N_24 VPW NCH W=0.58u L=0.06u
MNA2_2 VSS B N_26 VPW NCH W=0.58u L=0.06u
MPA2_4 Y B VDD VNW PCH W=0.59u L=0.06u
MNA1_2 Y A N_26 VPW NCH W=0.58u L=0.06u
MPA1_7 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1_6 Y A N_28 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.59u L=0.06u
MPA2_6 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2_6 VSS B N_28 VPW NCH W=0.58u L=0.06u
MNA2_7 VSS B N_30 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.59u L=0.06u
MNA1_7 Y A N_30 VPW NCH W=0.58u L=0.06u
MPA1_6 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1_4 Y A N_32 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.59u L=0.06u
MPA2_5 Y B VDD VNW PCH W=0.59u L=0.06u
MNA2_4 VSS B N_32 VPW NCH W=0.58u L=0.06u
MNA2_5 VSS B N_34 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.59u L=0.06u
MNA1_5 Y A N_34 VPW NCH W=0.58u L=0.06u
MPA1_5 Y A VDD VNW PCH W=0.59u L=0.06u
MNA1_3 Y A N_20 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.59u L=0.06u
MNA2_3 N_20 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.59u L=0.06u
.ENDS NAND2X8AA10TR

****
.SUBCKT NAND2X8BA10TR VDD VSS VPW VNW Y A B
MPA2_8 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2 VSS B N_39 VPW NCH W=0.58u L=0.06u
MPA1_8 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1 Y A N_39 VPW NCH W=0.58u L=0.06u
MNA1_8 Y A N_41 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.7u L=0.06u
MPA2_7 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2_8 VSS B N_41 VPW NCH W=0.58u L=0.06u
MNA2_2 VSS B N_43 VPW NCH W=0.58u L=0.06u
MPA2_4 Y B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y A N_43 VPW NCH W=0.58u L=0.06u
MPA1_7 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1_6 Y A N_45 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.7u L=0.06u
MPA2_6 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2_6 VSS B N_45 VPW NCH W=0.58u L=0.06u
MNA2_7 VSS B N_47 VPW NCH W=0.58u L=0.06u
MPA2_3 Y B VDD VNW PCH W=0.7u L=0.06u
MNA1_7 Y A N_47 VPW NCH W=0.58u L=0.06u
MPA1_6 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1_4 Y A N_49 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.7u L=0.06u
MPA2_5 Y B VDD VNW PCH W=0.7u L=0.06u
MNA2_4 VSS B N_49 VPW NCH W=0.58u L=0.06u
MNA2_5 VSS B N_51 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.7u L=0.06u
MNA1_5 Y A N_51 VPW NCH W=0.58u L=0.06u
MPA1_5 Y A VDD VNW PCH W=0.7u L=0.06u
MNA1_3 Y A N_37 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.7u L=0.06u
MNA2_3 N_37 B VSS VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.7u L=0.06u
.ENDS NAND2X8BA10TR

****
.SUBCKT NAND2XBX1P4MA10TR VDD VSS VPW VNW Y A BN
MPA106 NET24 BN VDD VNW PCH W=0.28u L=0.06u
MNA104 NET24 BN VSS VPW NCH W=0.21u L=0.06u
MNA2 N_17 NET24 VSS VPW NCH W=0.41u L=0.06u
MPA2_2 Y NET24 VDD VNW PCH W=0.34u L=0.06u
MNA1 Y A N_17 VPW NCH W=0.41u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.34u L=0.06u
MNA1_2 Y A N_15 VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.34u L=0.06u
MNA2_2 N_15 NET24 VSS VPW NCH W=0.41u L=0.06u
MPA2 Y NET24 VDD VNW PCH W=0.34u L=0.06u
.ENDS NAND2XBX1P4MA10TR

****
.SUBCKT NAND2XBX2MA10TR VDD VSS VPW VNW Y A BN
MPA106 NET24 BN VDD VNW PCH W=0.365u L=0.06u
MNA104 NET24 BN VSS VPW NCH W=0.275u L=0.06u
MNA2 N_18 NET24 VSS VPW NCH W=0.58u L=0.06u
MPA2_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1 Y A N_18 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y A N_16 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_2 N_16 NET24 VSS VPW NCH W=0.58u L=0.06u
MPA2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2XBX2MA10TR

****
.SUBCKT NAND2XBX3MA10TR VDD VSS VPW VNW Y A BN
MPA106 NET24 BN VDD VNW PCH W=0.56u L=0.06u
MNA104 NET24 BN VSS VPW NCH W=0.425u L=0.06u
MPA2_3 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_2 VSS NET24 N_22 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y A N_22 VPW NCH W=0.58u L=0.06u
MNA1 Y A N_24 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS NET24 N_24 VPW NCH W=0.58u L=0.06u
MPA2_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_3 VSS NET24 N_19 VPW NCH W=0.58u L=0.06u
MPA2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_3 N_19 A Y VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2XBX3MA10TR

****
.SUBCKT NAND2XBX4MA10TR VDD VSS VPW VNW Y A BN
MPA106 NET24 BN VDD VNW PCH W=0.7u L=0.06u
MNA104 NET24 BN VSS VPW NCH W=0.53u L=0.06u
MPA2_4 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_4 VSS NET24 N_26 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_4 Y A N_26 VPW NCH W=0.58u L=0.06u
MNA1 Y A N_28 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS NET24 N_28 VPW NCH W=0.58u L=0.06u
MPA2_3 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_3 VSS NET24 N_30 VPW NCH W=0.58u L=0.06u
MPA2_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y A N_30 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y A N_23 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_2 N_23 NET24 VSS VPW NCH W=0.58u L=0.06u
MPA2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2XBX4MA10TR

****
.SUBCKT NAND2XBX6MA10TR VDD VSS VPW VNW Y A BN
MNA104 NET24 BN VSS VPW NCH W=0.415u L=0.06u
MPA106_2 NET24 BN VDD VNW PCH W=0.55u L=0.06u
MPA106 NET24 BN VDD VNW PCH W=0.55u L=0.06u
MNA104_2 NET24 BN VSS VPW NCH W=0.415u L=0.06u
MPA2_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_2 VSS NET24 N_37 VPW NCH W=0.58u L=0.06u
MPA1_6 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y A N_37 VPW NCH W=0.58u L=0.06u
MNA1_5 Y A N_39 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_4 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_5 VSS NET24 N_39 VPW NCH W=0.58u L=0.06u
MNA2_6 VSS NET24 N_41 VPW NCH W=0.58u L=0.06u
MPA2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_6 Y A N_41 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1 Y A N_43 VPW NCH W=0.58u L=0.06u
MPA1_5 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_6 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS NET24 N_43 VPW NCH W=0.58u L=0.06u
MNA2_3 VSS NET24 N_45 VPW NCH W=0.58u L=0.06u
MPA2_3 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y A N_45 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_4 Y A N_33 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_4 N_33 NET24 VSS VPW NCH W=0.58u L=0.06u
MPA2_5 Y NET24 VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2XBX6MA10TR

****
.SUBCKT NAND2XBX8MA10TR VDD VSS VPW VNW Y A BN
MNA104 NET24 BN VSS VPW NCH W=0.53u L=0.06u
MPA106_2 NET24 BN VDD VNW PCH W=0.7u L=0.06u
MPA106 NET24 BN VDD VNW PCH W=0.7u L=0.06u
MNA104_2 NET24 BN VSS VPW NCH W=0.53u L=0.06u
MPA2_8 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2 VSS NET24 N_45 VPW NCH W=0.58u L=0.06u
MPA1_8 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1 Y A N_45 VPW NCH W=0.58u L=0.06u
MNA1_2 Y A N_47 VPW NCH W=0.58u L=0.06u
MPA1_4 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_7 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_2 VSS NET24 N_47 VPW NCH W=0.58u L=0.06u
MNA2_8 VSS NET24 N_49 VPW NCH W=0.58u L=0.06u
MPA2_4 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_8 Y A N_49 VPW NCH W=0.58u L=0.06u
MPA1_7 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_7 Y A N_51 VPW NCH W=0.58u L=0.06u
MPA1_3 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_6 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_7 VSS NET24 N_51 VPW NCH W=0.58u L=0.06u
MNA2_6 VSS NET24 N_53 VPW NCH W=0.58u L=0.06u
MPA2_3 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_6 Y A N_53 VPW NCH W=0.58u L=0.06u
MPA1_6 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_5 Y A N_55 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MPA2_5 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA2_5 VSS NET24 N_55 VPW NCH W=0.58u L=0.06u
MNA2_4 VSS NET24 N_57 VPW NCH W=0.58u L=0.06u
MPA2_2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
MNA1_4 Y A N_57 VPW NCH W=0.58u L=0.06u
MPA1_5 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y A N_41 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_3 N_41 NET24 VSS VPW NCH W=0.58u L=0.06u
MPA2 Y NET24 VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND2XBX8MA10TR

****
.SUBCKT NAND3BX1P4MA10TR VDD VSS VPW VNW Y AN B C
MPA1 NET14 AN VDD VNW PCH W=0.25u L=0.06u
MNA1 NET14 AN VSS VPW NCH W=0.19u L=0.06u
MPA3_2 Y C VDD VNW PCH W=0.25u L=0.06u
MNA3 N_22 C VSS VPW NCH W=0.41u L=0.06u
MNA2 N_22 B N_23 VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.25u L=0.06u
MNA102 Y NET14 N_23 VPW NCH W=0.41u L=0.06u
MPA105 Y NET14 VDD VNW PCH W=0.25u L=0.06u
MNA102_2 Y NET14 N_25 VPW NCH W=0.41u L=0.06u
MPA105_2 Y NET14 VDD VNW PCH W=0.25u L=0.06u
MNA2_2 N_25 B N_20 VPW NCH W=0.41u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.25u L=0.06u
MNA3_2 N_20 C VSS VPW NCH W=0.41u L=0.06u
MPA3 Y C VDD VNW PCH W=0.25u L=0.06u
.ENDS NAND3BX1P4MA10TR

****
.SUBCKT NAND3BX2MA10TR VDD VSS VPW VNW Y AN B C
MPA1 NET14 AN VDD VNW PCH W=0.33u L=0.06u
MNA1 NET14 AN VSS VPW NCH W=0.25u L=0.06u
MPA3_2 Y C VDD VNW PCH W=0.36u L=0.06u
MNA3 N_22 C VSS VPW NCH W=0.58u L=0.06u
MNA2 N_22 B N_23 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.36u L=0.06u
MNA102 Y NET14 N_23 VPW NCH W=0.58u L=0.06u
MPA105 Y NET14 VDD VNW PCH W=0.36u L=0.06u
MNA102_2 Y NET14 N_25 VPW NCH W=0.58u L=0.06u
MPA105_2 Y NET14 VDD VNW PCH W=0.36u L=0.06u
MNA2_2 N_25 B N_20 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.36u L=0.06u
MNA3_2 N_20 C VSS VPW NCH W=0.58u L=0.06u
MPA3 Y C VDD VNW PCH W=0.36u L=0.06u
.ENDS NAND3BX2MA10TR

****
.SUBCKT NAND3X1P4AA10TR VDD VSS VPW VNW Y A B C
MPA3_2 Y C VDD VNW PCH W=0.38u L=0.06u
MNA3 VSS C N_19 VPW NCH W=0.41u L=0.06u
MNA2 N_19 B N_20 VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.38u L=0.06u
MNA1 Y A N_20 VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.38u L=0.06u
MNA1_2 Y A N_22 VPW NCH W=0.41u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.38u L=0.06u
MNA2_2 N_22 B N_17 VPW NCH W=0.41u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.38u L=0.06u
MNA3_2 N_17 C VSS VPW NCH W=0.41u L=0.06u
MPA3 Y C VDD VNW PCH W=0.38u L=0.06u
.ENDS NAND3X1P4AA10TR

****
.SUBCKT NAND3X1P4MA10TR VDD VSS VPW VNW Y A B C
MNA3 VSS C N_13 VPW NCH W=0.41u L=0.06u
MNA2 N_13 B N_14 VPW NCH W=0.41u L=0.06u
MNA1 Y A N_14 VPW NCH W=0.41u L=0.06u
MNA1_2 Y A N_16 VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.5u L=0.06u
MNA2_2 N_16 B N_11 VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.5u L=0.06u
MNA3_2 N_11 C VSS VPW NCH W=0.41u L=0.06u
MPA3 Y C VDD VNW PCH W=0.5u L=0.06u
.ENDS NAND3X1P4MA10TR

****
.SUBCKT NAND3X2AA10TR VDD VSS VPW VNW Y A B C
MPA3_2 Y C VDD VNW PCH W=0.54u L=0.06u
MNA3 VSS C N_19 VPW NCH W=0.58u L=0.06u
MNA2 N_19 B N_20 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.54u L=0.06u
MNA1 Y A N_20 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.54u L=0.06u
MNA1_2 Y A N_22 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.54u L=0.06u
MNA2_2 N_22 B N_17 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.54u L=0.06u
MNA3_2 N_17 C VSS VPW NCH W=0.58u L=0.06u
MPA3 Y C VDD VNW PCH W=0.54u L=0.06u
.ENDS NAND3X2AA10TR

****
.SUBCKT NAND3XXBX1P4MA10TR VDD VSS VPW VNW Y A B CN
MPA1 NET14 CN VDD VNW PCH W=0.25u L=0.06u
MNA1 NET14 CN VSS VPW NCH W=0.19u L=0.06u
MPA3_2 Y NET14 VDD VNW PCH W=0.25u L=0.06u
MNA3 VSS NET14 N_22 VPW NCH W=0.41u L=0.06u
MNA2 N_22 B N_23 VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.25u L=0.06u
MNA102 Y A N_23 VPW NCH W=0.41u L=0.06u
MPA105 Y A VDD VNW PCH W=0.25u L=0.06u
MNA102_2 Y A N_25 VPW NCH W=0.41u L=0.06u
MPA105_2 Y A VDD VNW PCH W=0.25u L=0.06u
MNA2_2 N_25 B N_19 VPW NCH W=0.41u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.25u L=0.06u
MNA3_2 N_19 NET14 VSS VPW NCH W=0.41u L=0.06u
MPA3 Y NET14 VDD VNW PCH W=0.25u L=0.06u
.ENDS NAND3XXBX1P4MA10TR

****
.SUBCKT NAND3XXBX2MA10TR VDD VSS VPW VNW Y A B CN
MPA1 NET14 CN VDD VNW PCH W=0.33u L=0.06u
MNA1 NET14 CN VSS VPW NCH W=0.25u L=0.06u
MPA3_2 Y NET14 VDD VNW PCH W=0.36u L=0.06u
MNA3 N_22 NET14 VSS VPW NCH W=0.58u L=0.06u
MNA2 N_22 B N_23 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.36u L=0.06u
MNA102 Y A N_23 VPW NCH W=0.58u L=0.06u
MPA105 Y A VDD VNW PCH W=0.36u L=0.06u
MNA102_2 Y A N_25 VPW NCH W=0.58u L=0.06u
MPA105_2 Y A VDD VNW PCH W=0.36u L=0.06u
MNA2_2 N_25 B N_20 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.36u L=0.06u
MNA3_2 N_20 NET14 VSS VPW NCH W=0.58u L=0.06u
MPA3 Y NET14 VDD VNW PCH W=0.36u L=0.06u
.ENDS NAND3XXBX2MA10TR

****
.SUBCKT NAND4BX1P4MA10TR VDD VSS VPW VNW Y AN B C D
MPA1 NET32 AN VDD VNW PCH W=0.265u L=0.06u
MNA1 NET32 AN VSS VPW NCH W=0.2u L=0.06u
MNA4 N_20 D VSS VPW NCH W=0.41u L=0.06u
MNA3 N_21 C N_20 VPW NCH W=0.41u L=0.06u
MNA2 N_21 B N_22 VPW NCH W=0.41u L=0.06u
MNA102 Y NET32 N_22 VPW NCH W=0.41u L=0.06u
MPA105 Y NET32 VDD VNW PCH W=0.4u L=0.06u
MNA102_2 Y NET32 N_24 VPW NCH W=0.41u L=0.06u
MNA2_2 N_24 B N_25 VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.4u L=0.06u
MNA3_2 N_25 C N_17 VPW NCH W=0.41u L=0.06u
MPA3 Y C VDD VNW PCH W=0.4u L=0.06u
MNA4_2 N_17 D VSS VPW NCH W=0.41u L=0.06u
MPA4 Y D VDD VNW PCH W=0.4u L=0.06u
.ENDS NAND4BX1P4MA10TR

****
.SUBCKT NAND4BX2MA10TR VDD VSS VPW VNW Y AN B C D
MPA1 NET32 AN VDD VNW PCH W=0.34u L=0.06u
MNA1 NET32 AN VSS VPW NCH W=0.26u L=0.06u
MPA4_2 Y D VDD VNW PCH W=0.285u L=0.06u
MNA4 N_26 D VSS VPW NCH W=0.58u L=0.06u
MPA3 Y C VDD VNW PCH W=0.285u L=0.06u
MNA3 N_26 C N_27 VPW NCH W=0.58u L=0.06u
MNA2 N_27 B N_28 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.285u L=0.06u
MNA102 Y NET32 N_28 VPW NCH W=0.58u L=0.06u
MPA105_2 Y NET32 VDD VNW PCH W=0.285u L=0.06u
MNA102_2 Y NET32 N_30 VPW NCH W=0.58u L=0.06u
MPA105 Y NET32 VDD VNW PCH W=0.285u L=0.06u
MNA2_2 N_30 B N_31 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.285u L=0.06u
MNA3_2 N_31 C N_24 VPW NCH W=0.58u L=0.06u
MPA3_2 Y C VDD VNW PCH W=0.285u L=0.06u
MNA4_2 N_24 D VSS VPW NCH W=0.58u L=0.06u
MPA4 Y D VDD VNW PCH W=0.285u L=0.06u
.ENDS NAND4BX2MA10TR

****
.SUBCKT NAND4X1P4AA10TR VDD VSS VPW VNW Y A B C D
MPA4_2 Y D VDD VNW PCH W=0.335u L=0.06u
MNA4 VSS D N_23 VPW NCH W=0.41u L=0.06u
MPA3 Y C VDD VNW PCH W=0.335u L=0.06u
MNA3 N_23 C N_24 VPW NCH W=0.41u L=0.06u
MNA2 N_24 B N_25 VPW NCH W=0.41u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.335u L=0.06u
MNA1 Y A N_25 VPW NCH W=0.41u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.335u L=0.06u
MNA1_2 Y A N_27 VPW NCH W=0.41u L=0.06u
MPA1 Y A VDD VNW PCH W=0.335u L=0.06u
MNA2_2 N_27 B N_28 VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.335u L=0.06u
MNA3_2 N_28 C N_21 VPW NCH W=0.41u L=0.06u
MPA3_2 Y C VDD VNW PCH W=0.335u L=0.06u
MNA4_2 N_21 D VSS VPW NCH W=0.41u L=0.06u
MPA4 Y D VDD VNW PCH W=0.335u L=0.06u
.ENDS NAND4X1P4AA10TR

****
.SUBCKT NAND4X2AA10TR VDD VSS VPW VNW Y A B C D
MPA4_2 Y D VDD VNW PCH W=0.48u L=0.06u
MNA4 VSS D N_23 VPW NCH W=0.58u L=0.06u
MPA3 Y C VDD VNW PCH W=0.48u L=0.06u
MNA3 N_23 C N_24 VPW NCH W=0.58u L=0.06u
MNA2 N_24 B N_25 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA1 Y A N_25 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y A N_27 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.48u L=0.06u
MNA2_2 N_27 B N_28 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.48u L=0.06u
MNA3_2 N_28 C N_21 VPW NCH W=0.58u L=0.06u
MPA3_2 Y C VDD VNW PCH W=0.48u L=0.06u
MNA4_2 N_21 D VSS VPW NCH W=0.58u L=0.06u
MPA4 Y D VDD VNW PCH W=0.48u L=0.06u
.ENDS NAND4X2AA10TR

****
.SUBCKT NAND4X2MA10TR VDD VSS VPW VNW Y A B C D
MPA4_2 Y D VDD VNW PCH W=0.285u L=0.06u
MNA4 VSS D N_23 VPW NCH W=0.58u L=0.06u
MPA3 Y C VDD VNW PCH W=0.285u L=0.06u
MNA3 N_23 C N_24 VPW NCH W=0.58u L=0.06u
MNA2 N_24 B N_25 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.285u L=0.06u
MNA1 Y A N_25 VPW NCH W=0.58u L=0.06u
MPA1_2 Y A VDD VNW PCH W=0.285u L=0.06u
MNA1_2 Y A N_27 VPW NCH W=0.58u L=0.06u
MPA1 Y A VDD VNW PCH W=0.285u L=0.06u
MNA2_2 N_27 B N_28 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.285u L=0.06u
MNA3_2 N_28 C N_21 VPW NCH W=0.58u L=0.06u
MPA3_2 Y C VDD VNW PCH W=0.285u L=0.06u
MNA4_2 N_21 D VSS VPW NCH W=0.58u L=0.06u
MPA4 Y D VDD VNW PCH W=0.285u L=0.06u
.ENDS NAND4X2MA10TR

****
.SUBCKT NAND4XXXBX1P4MA10TR VDD VSS VPW VNW Y A B C DN
MPA1 NET32 DN VDD VNW PCH W=0.265u L=0.06u
MNA1 NET32 DN VSS VPW NCH W=0.2u L=0.06u
MNA4 N_20 NET32 VSS VPW NCH W=0.41u L=0.06u
MNA3 N_21 C N_20 VPW NCH W=0.41u L=0.06u
MNA2 N_21 B N_22 VPW NCH W=0.41u L=0.06u
MNA102 Y A N_22 VPW NCH W=0.41u L=0.06u
MPA105 Y A VDD VNW PCH W=0.4u L=0.06u
MNA102_2 Y A N_24 VPW NCH W=0.41u L=0.06u
MNA2_2 N_24 B N_25 VPW NCH W=0.41u L=0.06u
MPA2 Y B VDD VNW PCH W=0.4u L=0.06u
MNA3_2 N_25 C N_17 VPW NCH W=0.41u L=0.06u
MPA3 Y C VDD VNW PCH W=0.4u L=0.06u
MNA4_2 N_17 NET32 VSS VPW NCH W=0.41u L=0.06u
MPA4 Y NET32 VDD VNW PCH W=0.4u L=0.06u
.ENDS NAND4XXXBX1P4MA10TR

****
.SUBCKT NAND4XXXBX2MA10TR VDD VSS VPW VNW Y A B C DN
MPA1 NET32 DN VDD VNW PCH W=0.34u L=0.06u
MNA1 NET32 DN VSS VPW NCH W=0.26u L=0.06u
MPA4_2 Y NET32 VDD VNW PCH W=0.285u L=0.06u
MNA4 N_16 NET32 VSS VPW NCH W=0.58u L=0.06u
MPA3 Y C VDD VNW PCH W=0.285u L=0.06u
MNA3 N_16 C N_17 VPW NCH W=0.58u L=0.06u
MNA2 N_17 B N_18 VPW NCH W=0.58u L=0.06u
MPA2_2 Y B VDD VNW PCH W=0.285u L=0.06u
MNA102 Y A N_18 VPW NCH W=0.58u L=0.06u
MPA105_2 Y A VDD VNW PCH W=0.285u L=0.06u
MNA102_2 Y A N_20 VPW NCH W=0.58u L=0.06u
MPA105 Y A VDD VNW PCH W=0.285u L=0.06u
MNA2_2 N_20 B N_21 VPW NCH W=0.58u L=0.06u
MPA2 Y B VDD VNW PCH W=0.285u L=0.06u
MNA3_2 N_21 C N_14 VPW NCH W=0.58u L=0.06u
MPA3_2 Y C VDD VNW PCH W=0.285u L=0.06u
MNA4_2 N_14 NET32 VSS VPW NCH W=0.58u L=0.06u
MPA4 Y NET32 VDD VNW PCH W=0.285u L=0.06u
.ENDS NAND4XXXBX2MA10TR

****
.SUBCKT NOR2BX1P4MA10TR VDD VSS VPW VNW Y AN B
MNA104 NET24 AN VSS VPW NCH W=0.195u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.26u L=0.06u
MNA2 Y B VSS VPW NCH W=0.2u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.49u L=0.06u
MNA1 Y NET24 VSS VPW NCH W=0.2u L=0.06u
MPA1 Y NET24 N_5 VNW PCH W=0.49u L=0.06u
MPA1_2 Y NET24 N_3 VNW PCH W=0.49u L=0.06u
MNA1_2 Y NET24 VSS VPW NCH W=0.2u L=0.06u
MPA2_2 N_3 B VDD VNW PCH W=0.49u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.2u L=0.06u
.ENDS NOR2BX1P4MA10TR

****
.SUBCKT NOR2BX2MA10TR VDD VSS VPW VNW Y AN B
MNA104 NET24 AN VSS VPW NCH W=0.26u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.345u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1 Y NET24 N_5 VNW PCH W=0.7u L=0.06u
MPA1_2 Y NET24 N_3 VNW PCH W=0.7u L=0.06u
MNA1_2 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA2_2 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2BX2MA10TR

****
.SUBCKT NOR2BX3MA10TR VDD VSS VPW VNW Y AN B
MNA104 NET24 AN VSS VPW NCH W=0.4u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.53u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_6 VNW PCH W=0.7u L=0.06u
MNA1 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1 Y NET24 N_6 VNW PCH W=0.7u L=0.06u
MPA1_3 Y NET24 N_8 VNW PCH W=0.7u L=0.06u
MNA1_3 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA2_3 VDD B N_8 VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_2 VDD B N_3 VNW PCH W=0.7u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1_2 N_3 NET24 Y VNW PCH W=0.7u L=0.06u
MNA1_2 Y NET24 VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2BX3MA10TR

****
.SUBCKT NOR2BX4MA10TR VDD VSS VPW VNW Y AN B
MNA104 NET24 AN VSS VPW NCH W=0.52u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.69u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_6 VNW PCH W=0.7u L=0.06u
MNA1_2 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1 Y NET24 N_6 VNW PCH W=0.7u L=0.06u
MPA1_3 Y NET24 N_8 VNW PCH W=0.7u L=0.06u
MNA1_4 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_3 VDD B N_8 VNW PCH W=0.7u L=0.06u
MPA2_2 VDD B N_10 VNW PCH W=0.7u L=0.06u
MNA2_4 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y NET24 N_10 VNW PCH W=0.7u L=0.06u
MNA1 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1_4 Y NET24 N_3 VNW PCH W=0.7u L=0.06u
MNA1_3 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA2_4 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2BX4MA10TR

****
.SUBCKT NOR2BX6MA10TR VDD VSS VPW VNW Y AN B
MNA104 NET24 AN VSS VPW NCH W=0.39u L=0.06u
MPA106_2 NET24 AN VDD VNW PCH W=0.515u L=0.06u
MNA104_2 NET24 AN VSS VPW NCH W=0.39u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.515u L=0.06u
MNA2_4 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_5 VDD B N_7 VNW PCH W=0.7u L=0.06u
MNA1_2 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1_5 Y NET24 N_7 VNW PCH W=0.7u L=0.06u
MPA1_6 Y NET24 N_9 VNW PCH W=0.7u L=0.06u
MNA1_6 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MNA2_6 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_6 VDD B N_9 VNW PCH W=0.7u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_11 VNW PCH W=0.7u L=0.06u
MNA1_4 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1 Y NET24 N_11 VNW PCH W=0.7u L=0.06u
MPA1_3 Y NET24 N_13 VNW PCH W=0.7u L=0.06u
MNA1 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_3 VDD B N_13 VNW PCH W=0.7u L=0.06u
MPA2_4 VDD B N_15 VNW PCH W=0.7u L=0.06u
MNA2_5 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1_4 Y NET24 N_15 VNW PCH W=0.7u L=0.06u
MNA1_5 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y NET24 N_3 VNW PCH W=0.7u L=0.06u
MNA1_3 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA2_2 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2BX6MA10TR

****
.SUBCKT NOR2BX8MA10TR VDD VSS VPW VNW Y AN B
MNA104 NET24 AN VSS VPW NCH W=0.52u L=0.06u
MPA106_2 NET24 AN VDD VNW PCH W=0.69u L=0.06u
MNA104_2 NET24 AN VSS VPW NCH W=0.52u L=0.06u
MPA106 NET24 AN VDD VNW PCH W=0.69u L=0.06u
MNA2_8 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_7 VNW PCH W=0.7u L=0.06u
MNA1_8 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1 Y NET24 N_7 VNW PCH W=0.7u L=0.06u
MPA1_8 Y NET24 N_9 VNW PCH W=0.7u L=0.06u
MNA1_4 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MNA2_7 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_8 VDD B N_9 VNW PCH W=0.7u L=0.06u
MNA2_4 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_2 VDD B N_11 VNW PCH W=0.7u L=0.06u
MNA1_7 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y NET24 N_11 VNW PCH W=0.7u L=0.06u
MPA1_6 Y NET24 N_13 VNW PCH W=0.7u L=0.06u
MNA1_3 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MNA2_6 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_6 VDD B N_13 VNW PCH W=0.7u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_7 VDD B N_15 VNW PCH W=0.7u L=0.06u
MNA1_6 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1_7 Y NET24 N_15 VNW PCH W=0.7u L=0.06u
MPA1_4 Y NET24 N_17 VNW PCH W=0.7u L=0.06u
MNA1_2 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MNA2_5 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_4 VDD B N_17 VNW PCH W=0.7u L=0.06u
MPA2_5 VDD B N_19 VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1_5 Y NET24 N_19 VNW PCH W=0.7u L=0.06u
MNA1_5 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA1_3 Y NET24 N_3 VNW PCH W=0.7u L=0.06u
MNA1 Y NET24 VSS VPW NCH W=0.285u L=0.06u
MPA2_3 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2BX8MA10TR

****
.SUBCKT NOR2X1P4AA10TR VDD VSS VPW VNW Y A B
MNA2_2 Y B VSS VPW NCH W=0.345u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.49u L=0.06u
MNA1 Y A VSS VPW NCH W=0.345u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.49u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.345u L=0.06u
MPA1_2 Y A N_3 VNW PCH W=0.49u L=0.06u
MNA2 Y B VSS VPW NCH W=0.345u L=0.06u
MPA2_2 N_3 B VDD VNW PCH W=0.49u L=0.06u
.ENDS NOR2X1P4AA10TR

****
.SUBCKT NOR2X1P4MA10TR VDD VSS VPW VNW Y A B
MNA2_2 Y B VSS VPW NCH W=0.2u L=0.06u
MPA2 VDD B N_6 VNW PCH W=0.49u L=0.06u
MNA1 Y A VSS VPW NCH W=0.2u L=0.06u
MPA1 Y A N_6 VNW PCH W=0.49u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.2u L=0.06u
MPA1_2 Y A N_5 VNW PCH W=0.49u L=0.06u
MNA2 Y B VSS VPW NCH W=0.2u L=0.06u
MPA2_2 N_5 B VDD VNW PCH W=0.49u L=0.06u
.ENDS NOR2X1P4MA10TR

****
.SUBCKT XNOR2X1P4MA10TR VDD VSS VPW VNW Y A B
MNA108 NIN1 A VSS VPW NCH W=0.53u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.7u L=0.06u
MNA1_2 NIN2 B VSS VPW NCH W=0.33u L=0.06u
MPA1_2 NIN2 B VDD VNW PCH W=0.49u L=0.06u
MNA1 NIN2 B VSS VPW NCH W=0.33u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.49u L=0.06u
MNOE_2 Y NIN1 NIN2 VPW NCH W=0.33u L=0.06u
MPOEN Y A NIN2 VNW PCH W=0.33u L=0.06u
MNOE Y NIN1 NIN2 VPW NCH W=0.33u L=0.06u
MPOEN_2 Y A NIN2 VNW PCH W=0.33u L=0.06u
MNOE02_2 Y A BIN2 VPW NCH W=0.33u L=0.06u
MPOEN04 Y NIN1 BIN2 VNW PCH W=0.33u L=0.06u
MNOE02 Y A BIN2 VPW NCH W=0.33u L=0.06u
MPOEN04_2 Y NIN1 BIN2 VNW PCH W=0.33u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.33u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.66u L=0.06u
MNA1012_2 BIN2 NIN2 VSS VPW NCH W=0.33u L=0.06u
.ENDS XNOR2X1P4MA10TR

****
.SUBCKT NOR2X2AA10TR VDD VSS VPW VNW Y A B
MNA2_2 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MPA1_2 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.49u L=0.06u
MPA2_2 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.49u L=0.06u
.ENDS NOR2X2AA10TR

****
.SUBCKT NOR2X2MA10TR VDD VSS VPW VNW Y A B
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MPA1_2 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
MPA2_2 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2X2MA10TR

****
.SUBCKT XNOR2X2MA10TR VDD VSS VPW VNW Y A B
MNA108_2 NIN1 A VSS VPW NCH W=0.33u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.44u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.33u L=0.06u
MPA1010_2 NIN1 A VDD VNW PCH W=0.44u L=0.06u
MNA1_2 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_2 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNOE Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MPOEN Y A NIN2 VNW PCH W=0.47u L=0.06u
MNOE_2 Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_2 Y A NIN2 VNW PCH W=0.47u L=0.06u
MNOE02_2 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_2 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
MNOE02 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
MNA1012_2 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_2 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
.ENDS XNOR2X2MA10TR

****
.SUBCKT NOR2X3AA10TR VDD VSS VPW VNW Y A B
MNA2_3 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1_3 Y A N_7 VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_3 VDD B N_7 VNW PCH W=0.7u L=0.06u
MPA2_2 VDD B N_3 VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.49u L=0.06u
MPA1_2 N_3 A Y VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.49u L=0.06u
.ENDS NOR2X3AA10TR

****
.SUBCKT NOR2X3MA10TR VDD VSS VPW VNW Y A B
MNA2_3 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_3 Y A N_7 VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_3 VDD B N_7 VNW PCH W=0.7u L=0.06u
MPA2_2 VDD B N_3 VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1_2 N_3 A Y VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2X3MA10TR

****
.SUBCKT XNOR2X3MA10TR VDD VSS VPW VNW Y A B
MNA108 NIN1 A VSS VPW NCH W=0.485u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.645u L=0.06u
MNA108_2 NIN1 A VSS VPW NCH W=0.485u L=0.06u
MPA1010_2 NIN1 A VDD VNW PCH W=0.645u L=0.06u
MNA1 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_2 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_3 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_3 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNOE_2 Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MPOEN Y A NIN2 VNW PCH W=0.47u L=0.06u
MNOE Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_3 Y A NIN2 VNW PCH W=0.47u L=0.06u
MNOE_3 Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_2 Y A NIN2 VNW PCH W=0.47u L=0.06u
MNOE02_2 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
MNOE02 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_3 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
MNOE02_3 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_2 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
MNA1012_2 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_3 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MPA1014_2 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012_3 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
.ENDS XNOR2X3MA10TR

****
.SUBCKT NOR2X4AA10TR VDD VSS VPW VNW Y A B
MNA2_4 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1_4 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MPA1_3 Y A N_7 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.49u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_3 VDD B N_7 VNW PCH W=0.7u L=0.06u
MPA2_2 VDD B N_9 VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.49u L=0.06u
MPA1_2 Y A N_9 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1_4 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.49u L=0.06u
MPA2_4 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.49u L=0.06u
.ENDS NOR2X4AA10TR

****
.SUBCKT NOR2X4MA10TR VDD VSS VPW VNW Y A B
MNA2_4 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1_4 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_3 Y A N_7 VNW PCH W=0.7u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_3 VDD B N_7 VNW PCH W=0.7u L=0.06u
MPA2_2 VDD B N_9 VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y A N_9 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_4 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MPA2_4 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2X4MA10TR

****
.SUBCKT XNOR2X4MA10TR VDD VSS VPW VNW Y A B
MNA108_3 NIN1 A VSS VPW NCH W=0.415u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.55u L=0.06u
MNA108_2 NIN1 A VSS VPW NCH W=0.415u L=0.06u
MPA1010_3 NIN1 A VDD VNW PCH W=0.55u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.415u L=0.06u
MPA1010_2 NIN1 A VDD VNW PCH W=0.55u L=0.06u
MNA1_4 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_2 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_3 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_4 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_3 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNOE_4 Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_4 Y A NIN2 VNW PCH W=0.47u L=0.06u
MNOE_3 Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_3 Y A NIN2 VNW PCH W=0.47u L=0.06u
MNOE_2 Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_2 Y A NIN2 VNW PCH W=0.47u L=0.06u
MNOE Y NIN1 NIN2 VPW NCH W=0.47u L=0.06u
MPOEN Y A NIN2 VNW PCH W=0.47u L=0.06u
MNOE02_4 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_4 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
MNOE02_3 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_3 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
MNOE02_2 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_2 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
MNOE02 Y A BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04 Y NIN1 BIN2 VNW PCH W=0.47u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_3 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012_3 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_2 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012_2 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_4 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012_4 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
.ENDS XNOR2X4MA10TR

****
.SUBCKT NOR2X6AA10TR VDD VSS VPW VNW Y A B
MNA2_2 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_5 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1_6 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1_5 Y A N_5 VNW PCH W=0.7u L=0.06u
MPA1_6 Y A N_7 VNW PCH W=0.7u L=0.06u
MNA1_4 Y A VSS VPW NCH W=0.49u L=0.06u
MNA2_4 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_6 VDD B N_7 VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2 VDD B N_9 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1 Y A N_9 VNW PCH W=0.7u L=0.06u
MPA1_3 Y A N_11 VNW PCH W=0.7u L=0.06u
MNA1_5 Y A VSS VPW NCH W=0.49u L=0.06u
MNA2_6 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_3 VDD B N_11 VNW PCH W=0.7u L=0.06u
MPA2_4 VDD B N_13 VNW PCH W=0.7u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.49u L=0.06u
MPA1_4 Y A N_13 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1_2 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.49u L=0.06u
MPA2_2 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2_5 Y B VSS VPW NCH W=0.49u L=0.06u
.ENDS NOR2X6AA10TR

****
.SUBCKT NOR2X6MA10TR VDD VSS VPW VNW Y A B
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_5 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1_6 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_5 Y A N_5 VNW PCH W=0.7u L=0.06u
MPA1_6 Y A N_7 VNW PCH W=0.7u L=0.06u
MNA1_4 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_4 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_6 VDD B N_7 VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_9 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_9 VNW PCH W=0.7u L=0.06u
MPA1_3 Y A N_11 VNW PCH W=0.7u L=0.06u
MNA1_5 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_6 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_3 VDD B N_11 VNW PCH W=0.7u L=0.06u
MPA2_4 VDD B N_13 VNW PCH W=0.7u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1_4 Y A N_13 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MPA2_2 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2_5 Y B VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2X6MA10TR

****
.SUBCKT NOR2X8AA10TR VDD VSS VPW VNW Y A B
MNA2_8 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1_8 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MPA1_8 Y A N_7 VNW PCH W=0.7u L=0.06u
MNA1_4 Y A VSS VPW NCH W=0.49u L=0.06u
MNA2_7 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_8 VDD B N_7 VNW PCH W=0.7u L=0.06u
MNA2_4 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_2 VDD B N_9 VNW PCH W=0.7u L=0.06u
MNA1_7 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1_2 Y A N_9 VNW PCH W=0.7u L=0.06u
MPA1_6 Y A N_11 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.49u L=0.06u
MNA2_6 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_6 VDD B N_11 VNW PCH W=0.7u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_7 VDD B N_13 VNW PCH W=0.7u L=0.06u
MNA1_6 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1_7 Y A N_13 VNW PCH W=0.7u L=0.06u
MPA1_4 Y A N_15 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.49u L=0.06u
MNA2_5 Y B VSS VPW NCH W=0.49u L=0.06u
MPA2_4 VDD B N_15 VNW PCH W=0.7u L=0.06u
MPA2_5 VDD B N_17 VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.49u L=0.06u
MPA1_5 Y A N_17 VNW PCH W=0.7u L=0.06u
MNA1_5 Y A VSS VPW NCH W=0.49u L=0.06u
MPA1_3 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.49u L=0.06u
MPA2_3 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.49u L=0.06u
.ENDS NOR2X8AA10TR

****
.SUBCKT NOR2X8MA10TR VDD VSS VPW VNW Y A B
MNA2_8 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.7u L=0.06u
MNA1_8 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MPA1_8 Y A N_7 VNW PCH W=0.7u L=0.06u
MNA1_4 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_7 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_8 VDD B N_7 VNW PCH W=0.7u L=0.06u
MNA2_4 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_2 VDD B N_9 VNW PCH W=0.7u L=0.06u
MNA1_7 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y A N_9 VNW PCH W=0.7u L=0.06u
MPA1_6 Y A N_11 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_6 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_6 VDD B N_11 VNW PCH W=0.7u L=0.06u
MNA2_3 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_7 VDD B N_13 VNW PCH W=0.7u L=0.06u
MNA1_6 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_7 Y A N_13 VNW PCH W=0.7u L=0.06u
MPA1_4 Y A N_15 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_5 Y B VSS VPW NCH W=0.285u L=0.06u
MPA2_4 VDD B N_15 VNW PCH W=0.7u L=0.06u
MPA2_5 VDD B N_17 VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.285u L=0.06u
MPA1_5 Y A N_17 VNW PCH W=0.7u L=0.06u
MNA1_5 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_3 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MPA2_3 N_3 B VDD VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2X8MA10TR

****
.SUBCKT NOR2XBX1P4MA10TR VDD VSS VPW VNW Y A BN
MNA104 NET014 BN VSS VPW NCH W=0.195u L=0.06u
MPA106 NET014 BN VDD VNW PCH W=0.26u L=0.06u
MNA2 Y NET014 VSS VPW NCH W=0.2u L=0.06u
MPA2 VDD NET014 N_6 VNW PCH W=0.49u L=0.06u
MNA1 Y A VSS VPW NCH W=0.2u L=0.06u
MPA1 Y A N_6 VNW PCH W=0.49u L=0.06u
MPA1_2 Y A N_3 VNW PCH W=0.49u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.2u L=0.06u
MPA2_2 N_3 NET014 VDD VNW PCH W=0.49u L=0.06u
MNA2_2 Y NET014 VSS VPW NCH W=0.2u L=0.06u
.ENDS NOR2XBX1P4MA10TR

****
.SUBCKT NOR2XBX2MA10TR VDD VSS VPW VNW Y A BN
MNA104 NET014 BN VSS VPW NCH W=0.26u L=0.06u
MPA106 NET014 BN VDD VNW PCH W=0.345u L=0.06u
MNA2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD NET014 N_5 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MPA1_2 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
MPA2_2 N_3 NET014 VDD VNW PCH W=0.7u L=0.06u
MNA2_2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2XBX2MA10TR

****
.SUBCKT NOR2XBX3MA10TR VDD VSS VPW VNW Y A BN
MNA104 NET014 BN VSS VPW NCH W=0.4u L=0.06u
MPA106 NET014 BN VDD VNW PCH W=0.53u L=0.06u
MNA2_2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD NET014 N_5 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_5 VNW PCH W=0.7u L=0.06u
MPA1_3 Y A N_7 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.285u L=0.06u
MPA2_3 VDD NET014 N_7 VNW PCH W=0.7u L=0.06u
MNA2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_2 VDD NET014 N_3 VNW PCH W=0.7u L=0.06u
MNA2_3 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA1_2 N_3 A Y VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2XBX3MA10TR

****
.SUBCKT NOR2XBX4MA10TR VDD VSS VPW VNW Y A BN
MNA104 NET014 BN VSS VPW NCH W=0.52u L=0.06u
MPA106 NET014 BN VDD VNW PCH W=0.69u L=0.06u
MNA2_2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD NET014 N_6 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_6 VNW PCH W=0.7u L=0.06u
MPA1_3 Y A N_8 VNW PCH W=0.7u L=0.06u
MNA1_4 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_3 VDD NET014 N_8 VNW PCH W=0.7u L=0.06u
MPA2_2 VDD NET014 N_10 VNW PCH W=0.7u L=0.06u
MNA2_4 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y A N_10 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_4 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.285u L=0.06u
MPA2_4 N_3 NET014 VDD VNW PCH W=0.7u L=0.06u
MNA2_3 Y NET014 VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2XBX4MA10TR

****
.SUBCKT NOR2XBX6MA10TR VDD VSS VPW VNW Y A BN
MNA104 NET014 BN VSS VPW NCH W=0.39u L=0.06u
MPA106_2 NET014 BN VDD VNW PCH W=0.515u L=0.06u
MNA104_2 NET014 BN VSS VPW NCH W=0.39u L=0.06u
MPA106 NET014 BN VDD VNW PCH W=0.515u L=0.06u
MNA2_4 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_5 VDD NET014 N_7 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_5 Y A N_7 VNW PCH W=0.7u L=0.06u
MPA1_6 Y A N_9 VNW PCH W=0.7u L=0.06u
MNA1_6 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_6 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_6 VDD NET014 N_9 VNW PCH W=0.7u L=0.06u
MNA2_3 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD NET014 N_11 VNW PCH W=0.7u L=0.06u
MNA1_4 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_11 VNW PCH W=0.7u L=0.06u
MPA1_3 Y A N_13 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_3 VDD NET014 N_13 VNW PCH W=0.7u L=0.06u
MPA2_4 VDD NET014 N_15 VNW PCH W=0.7u L=0.06u
MNA2_5 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA1_4 Y A N_15 VNW PCH W=0.7u L=0.06u
MNA1_5 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y A N_3 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.285u L=0.06u
MPA2_2 N_3 NET014 VDD VNW PCH W=0.7u L=0.06u
MNA2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2XBX6MA10TR

****
.SUBCKT NOR2XBX8MA10TR VDD VSS VPW VNW Y A BN
MNA104 NET014 BN VSS VPW NCH W=0.52u L=0.06u
MPA106_2 NET014 BN VDD VNW PCH W=0.69u L=0.06u
MNA104_2 NET014 BN VSS VPW NCH W=0.52u L=0.06u
MPA106 NET014 BN VDD VNW PCH W=0.69u L=0.06u
MNA2_8 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD NET014 N_88 VNW PCH W=0.7u L=0.06u
MNA1_8 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1 Y A N_88 VNW PCH W=0.7u L=0.06u
MPA1_8 Y A N_90 VNW PCH W=0.7u L=0.06u
MNA1_4 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_7 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_8 VDD NET014 N_90 VNW PCH W=0.7u L=0.06u
MNA2_4 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_2 VDD NET014 N_92 VNW PCH W=0.7u L=0.06u
MNA1_7 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_2 Y A N_92 VNW PCH W=0.7u L=0.06u
MPA1_6 Y A N_94 VNW PCH W=0.7u L=0.06u
MNA1_3 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_6 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_6 VDD NET014 N_94 VNW PCH W=0.7u L=0.06u
MNA2_3 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_7 VDD NET014 N_96 VNW PCH W=0.7u L=0.06u
MNA1_6 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_7 Y A N_96 VNW PCH W=0.7u L=0.06u
MPA1_4 Y A N_98 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.285u L=0.06u
MNA2_5 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA2_4 VDD NET014 N_98 VNW PCH W=0.7u L=0.06u
MPA2_5 VDD NET014 N_100 VNW PCH W=0.7u L=0.06u
MNA2_2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
MPA1_5 Y A N_100 VNW PCH W=0.7u L=0.06u
MNA1_5 Y A VSS VPW NCH W=0.285u L=0.06u
MPA1_3 Y A N_84 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.285u L=0.06u
MPA2_3 N_84 NET014 VDD VNW PCH W=0.7u L=0.06u
MNA2 Y NET014 VSS VPW NCH W=0.285u L=0.06u
.ENDS NOR2XBX8MA10TR

****
.SUBCKT NOR3X1P4AA10TR VDD VSS VPW VNW Y A B C
MNA3_2 Y C VSS VPW NCH W=0.265u L=0.06u
MPA3 VDD C N_5 VNW PCH W=0.49u L=0.06u
MNA2 Y B VSS VPW NCH W=0.265u L=0.06u
MPA2 N_5 B N_6 VNW PCH W=0.49u L=0.06u
MNA1 Y A VSS VPW NCH W=0.265u L=0.06u
MPA1 Y A N_6 VNW PCH W=0.49u L=0.06u
MPA1_2 Y A N_8 VNW PCH W=0.49u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.265u L=0.06u
MPA2_2 N_8 B N_3 VNW PCH W=0.49u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.265u L=0.06u
MPA3_2 N_3 C VDD VNW PCH W=0.49u L=0.06u
MNA3 Y C VSS VPW NCH W=0.265u L=0.06u
.ENDS NOR3X1P4AA10TR

****
.SUBCKT XNOR3X1P4MA10TR VDD VSS VPW VNW Y A B C
MNA1020 NIN2 B VSS VPW NCH W=0.53u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 NIN3 C VSS VPW NCH W=0.33u L=0.06u
MPA1_2 NIN3 C VDD VNW PCH W=0.495u L=0.06u
MNA1 NIN3 C VSS VPW NCH W=0.33u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=0.495u L=0.06u
MNOE_2 XOR23 B NIN3 VPW NCH W=0.33u L=0.06u
MPOEN_2 XOR23 NIN2 NIN3 VNW PCH W=0.33u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.33u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.33u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.33u L=0.06u
MPOEN04_2 XOR23 B BIN3 VNW PCH W=0.33u L=0.06u
MNOE02_2 XOR23 NIN2 BIN3 VPW NCH W=0.33u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.33u L=0.06u
MNA1028_2 BIN3 NIN3 VSS VPW NCH W=0.33u L=0.06u
MPA1030_2 BIN3 NIN3 VDD VNW PCH W=0.495u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.33u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=0.495u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.395u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.525u L=0.06u
MNOE08 NOUT NIN1 XOR23 VPW NCH W=0.47u L=0.06u
MPOEN010 NOUT A XOR23 VNW PCH W=0.57u L=0.06u
MNOE012 NOUT A XNOR23 VPW NCH W=0.47u L=0.06u
MPOEN014 NOUT NIN1 XNOR23 VNW PCH W=0.57u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.47u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.7u L=0.06u
MNA1032_2 Y NOUT VSS VPW NCH W=0.37u L=0.06u
MPA1034_2 Y NOUT VDD VNW PCH W=0.49u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=0.37u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=0.49u L=0.06u
.ENDS XNOR3X1P4MA10TR

****
.SUBCKT NOR3X2AA10TR VDD VSS VPW VNW Y A B C
MNA3_2 Y C VSS VPW NCH W=0.38u L=0.06u
MPA3 VDD C N_5 VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.38u L=0.06u
MPA2 N_5 B N_6 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.38u L=0.06u
MPA1 Y A N_6 VNW PCH W=0.7u L=0.06u
MPA1_2 Y A N_8 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.38u L=0.06u
MPA2_2 N_8 B N_3 VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.38u L=0.06u
MPA3_2 N_3 C VDD VNW PCH W=0.7u L=0.06u
MNA3 Y C VSS VPW NCH W=0.38u L=0.06u
.ENDS NOR3X2AA10TR

****
.SUBCKT NOR3X2MA10TR VDD VSS VPW VNW Y A B C
MNA3_2 Y C VSS VPW NCH W=0.205u L=0.06u
MPA3 VDD C N_5 VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.205u L=0.06u
MPA2 N_5 B N_6 VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.205u L=0.06u
MPA1 Y A N_6 VNW PCH W=0.7u L=0.06u
MPA1_2 Y A N_8 VNW PCH W=0.7u L=0.06u
MNA1_2 Y A VSS VPW NCH W=0.205u L=0.06u
MPA2_2 N_8 B N_3 VNW PCH W=0.7u L=0.06u
MNA2_2 Y B VSS VPW NCH W=0.205u L=0.06u
MPA3_2 N_3 C VDD VNW PCH W=0.7u L=0.06u
MNA3 Y C VSS VPW NCH W=0.205u L=0.06u
.ENDS NOR3X2MA10TR

****
.SUBCKT XNOR3X2MA10TR VDD VSS VPW VNW Y A B C
MNA1020_2 NIN2 B VSS VPW NCH W=0.36u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.48u L=0.06u
MNA1020 NIN2 B VSS VPW NCH W=0.36u L=0.06u
MPA1022_2 NIN2 B VDD VNW PCH W=0.48u L=0.06u
MNA1 NIN3 C VSS VPW NCH W=0.445u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=0.665u L=0.06u
MNA1_2 NIN3 C VSS VPW NCH W=0.445u L=0.06u
MPA1_2 NIN3 C VDD VNW PCH W=0.665u L=0.06u
MNOE_2 XOR23 B NIN3 VPW NCH W=0.445u L=0.06u
MPOEN_2 XOR23 NIN2 NIN3 VNW PCH W=0.445u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.445u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.445u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.445u L=0.06u
MPOEN04_2 XOR23 B BIN3 VNW PCH W=0.445u L=0.06u
MNOE02_2 XOR23 NIN2 BIN3 VPW NCH W=0.445u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.445u L=0.06u
MNA1028_2 BIN3 NIN3 VSS VPW NCH W=0.445u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=0.665u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.445u L=0.06u
MPA1030_2 BIN3 NIN3 VDD VNW PCH W=0.665u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.47u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.63u L=0.06u
MNOE08_2 NOUT NIN1 XOR23 VPW NCH W=0.315u L=0.06u
MPOEN010_2 NOUT A XOR23 VNW PCH W=0.385u L=0.06u
MNOE08 NOUT NIN1 XOR23 VPW NCH W=0.315u L=0.06u
MPOEN010 NOUT A XOR23 VNW PCH W=0.385u L=0.06u
MNOE012 NOUT A XNOR23 VPW NCH W=0.315u L=0.06u
MPOEN014_2 NOUT NIN1 XNOR23 VNW PCH W=0.385u L=0.06u
MNOE012_2 NOUT A XNOR23 VPW NCH W=0.315u L=0.06u
MPOEN014 NOUT NIN1 XNOR23 VNW PCH W=0.385u L=0.06u
MNA1016_2 XNOR23 XOR23 VSS VPW NCH W=0.315u L=0.06u
MPA1018_2 XNOR23 XOR23 VDD VNW PCH W=0.47u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.315u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.47u L=0.06u
MNA1032_2 Y NOUT VSS VPW NCH W=0.53u L=0.06u
MPA1034_2 Y NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=0.53u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS XNOR3X2MA10TR

****
.SUBCKT OA211X1MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MPC2_2 VDD A1 N_5 VNW PCH W=0.41u L=0.06u
MPC1_2 INT A0 N_5 VNW PCH W=0.41u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.64u L=0.06u
MPC1 INT A0 N_7 VNW PCH W=0.41u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.64u L=0.06u
MPC2 N_7 A1 VDD VNW PCH W=0.41u L=0.06u
MNB1 N_23 B0 N1 VPW NCH W=0.64u L=0.06u
MPB1 INT B0 VDD VNW PCH W=0.38u L=0.06u
MNA1 N_23 C0 INT VPW NCH W=0.64u L=0.06u
MPA1 INT C0 VDD VNW PCH W=0.38u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OA211X1MA10TR

****
.SUBCKT OA211X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MNC2 N1 A1 VSS VPW NCH W=0.44u L=0.06u
MPC2 VDD A1 N_8 VNW PCH W=0.57u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.44u L=0.06u
MPC1 INT A0 N_8 VNW PCH W=0.57u L=0.06u
MPC1_2 INT A0 N_11 VNW PCH W=0.57u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.44u L=0.06u
MPC2_2 N_11 A1 VDD VNW PCH W=0.57u L=0.06u
MNC2_2 N1 A1 VSS VPW NCH W=0.44u L=0.06u
MNB1_2 N1 B0 N_32 VPW NCH W=0.44u L=0.06u
MPB1 INT B0 VDD VNW PCH W=0.53u L=0.06u
MPA1 INT C0 VDD VNW PCH W=0.53u L=0.06u
MNA1_2 INT C0 N_32 VPW NCH W=0.44u L=0.06u
MNA1 N_26 C0 INT VPW NCH W=0.44u L=0.06u
MNB1 N1 B0 N_26 VPW NCH W=0.44u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA108_2 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1010_2 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS OA211X1P4MA10TR

****
.SUBCKT OA211X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MNC2_2 N1 A1 VSS VPW NCH W=0.525u L=0.06u
MPC2 VDD A1 N_5 VNW PCH W=0.68u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.525u L=0.06u
MPC1 INT A0 N_5 VNW PCH W=0.68u L=0.06u
MPC1_2 INT A0 N_8 VNW PCH W=0.68u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.525u L=0.06u
MPC2_2 N_8 A1 VDD VNW PCH W=0.68u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.525u L=0.06u
MNB1 N_24 B0 N1 VPW NCH W=0.525u L=0.06u
MPB1_2 INT B0 VDD VNW PCH W=0.32u L=0.06u
MNA1 INT C0 N_24 VPW NCH W=0.525u L=0.06u
MPA1_2 INT C0 VDD VNW PCH W=0.32u L=0.06u
MNA1_2 INT C0 N_18 VPW NCH W=0.525u L=0.06u
MPA1 INT C0 VDD VNW PCH W=0.32u L=0.06u
MNB1_2 N_18 B0 N1 VPW NCH W=0.525u L=0.06u
MPB1 INT B0 VDD VNW PCH W=0.32u L=0.06u
MNA108_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OA211X2MA10TR

****
.SUBCKT OA211X3MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MNC1_2 N1 A0 VSS VPW NCH W=0.495u L=0.06u
MPC1_3 INT A0 N_5 VNW PCH W=0.64u L=0.06u
MNC2_3 N1 A1 VSS VPW NCH W=0.495u L=0.06u
MPC2_3 VDD A1 N_5 VNW PCH W=0.64u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.495u L=0.06u
MPC2_2 VDD A1 N_7 VNW PCH W=0.645u L=0.06u
MNC1_3 N1 A0 VSS VPW NCH W=0.495u L=0.06u
MPC1_2 INT A0 N_7 VNW PCH W=0.645u L=0.06u
MPC1 INT A0 N_9 VNW PCH W=0.645u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.495u L=0.06u
MPC2 N_9 A1 VDD VNW PCH W=0.645u L=0.06u
MNC2_2 N1 A1 VSS VPW NCH W=0.495u L=0.06u
MNB1_2 N1 B0 N_41 VPW NCH W=0.495u L=0.06u
MPB1_2 INT B0 VDD VNW PCH W=0.45u L=0.06u
MNA1_2 INT C0 N_41 VPW NCH W=0.495u L=0.06u
MPA1_2 INT C0 VDD VNW PCH W=0.45u L=0.06u
MNA1 INT C0 N_43 VPW NCH W=0.495u L=0.06u
MPA1 INT C0 VDD VNW PCH W=0.45u L=0.06u
MNB1 N1 B0 N_43 VPW NCH W=0.495u L=0.06u
MPB1 INT B0 VDD VNW PCH W=0.45u L=0.06u
MNB1_3 N_33 B0 N1 VPW NCH W=0.495u L=0.06u
MNA1_3 INT C0 N_33 VPW NCH W=0.495u L=0.06u
MNA108_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OA211X3MA10TR

****
.SUBCKT OA211X4MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MNC2_4 N1 A1 VSS VPW NCH W=0.495u L=0.06u
MPC2_3 VDD A1 N_5 VNW PCH W=0.64u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.495u L=0.06u
MPC1_3 INT A0 N_5 VNW PCH W=0.64u L=0.06u
MPC1_4 INT A0 N_7 VNW PCH W=0.64u L=0.06u
MNC1_4 N1 A0 VSS VPW NCH W=0.495u L=0.06u
MNC2_3 N1 A1 VSS VPW NCH W=0.495u L=0.06u
MPC2_4 VDD A1 N_7 VNW PCH W=0.64u L=0.06u
MNC2_2 N1 A1 VSS VPW NCH W=0.495u L=0.06u
MPC2 VDD A1 N_9 VNW PCH W=0.64u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.495u L=0.06u
MPC1 INT A0 N_9 VNW PCH W=0.64u L=0.06u
MPC1_2 INT A0 N_11 VNW PCH W=0.64u L=0.06u
MNC1_3 N1 A0 VSS VPW NCH W=0.495u L=0.06u
MPC2_2 N_11 A1 VDD VNW PCH W=0.64u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.495u L=0.06u
MPB1_3 INT B0 VDD VNW PCH W=0.4u L=0.06u
MNB1_3 N1 B0 N_53 VPW NCH W=0.495u L=0.06u
MPA1_3 INT C0 VDD VNW PCH W=0.4u L=0.06u
MNA1_3 INT C0 N_53 VPW NCH W=0.495u L=0.06u
MNA1_4 INT C0 N_55 VPW NCH W=0.495u L=0.06u
MPA1_2 INT C0 VDD VNW PCH W=0.4u L=0.06u
MNB1_4 N1 B0 N_55 VPW NCH W=0.495u L=0.06u
MPB1_2 INT B0 VDD VNW PCH W=0.4u L=0.06u
MNB1 N1 B0 N_57 VPW NCH W=0.495u L=0.06u
MPB1 INT B0 VDD VNW PCH W=0.4u L=0.06u
MNA1 INT C0 N_57 VPW NCH W=0.495u L=0.06u
MPA1 INT C0 VDD VNW PCH W=0.4u L=0.06u
MNA1_2 N_43 C0 INT VPW NCH W=0.495u L=0.06u
MNB1_2 N1 B0 N_43 VPW NCH W=0.495u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_4 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OA211X4MA10TR

****
.SUBCKT OA211X6MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MNC2_5 N1 A1 VSS VPW NCH W=0.49u L=0.06u
MPC2_6 VDD A1 N_5 VNW PCH W=0.63u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.49u L=0.06u
MPC1_6 INT A0 N_5 VNW PCH W=0.63u L=0.06u
MPC1_5 INT A0 N_7 VNW PCH W=0.63u L=0.06u
MNC1_6 N1 A0 VSS VPW NCH W=0.49u L=0.06u
MNC2_3 N1 A1 VSS VPW NCH W=0.49u L=0.06u
MPC2_5 VDD A1 N_7 VNW PCH W=0.63u L=0.06u
MNC2_2 N1 A1 VSS VPW NCH W=0.49u L=0.06u
MPC2_2 VDD A1 N_9 VNW PCH W=0.63u L=0.06u
MNC1_5 N1 A0 VSS VPW NCH W=0.49u L=0.06u
MPC1_2 INT A0 N_9 VNW PCH W=0.63u L=0.06u
MPC1_4 INT A0 N_11 VNW PCH W=0.63u L=0.06u
MNC1_4 N1 A0 VSS VPW NCH W=0.49u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.49u L=0.06u
MPC2_4 VDD A1 N_11 VNW PCH W=0.63u L=0.06u
MNC2_6 N1 A1 VSS VPW NCH W=0.49u L=0.06u
MPC2_3 VDD A1 N_13 VNW PCH W=0.63u L=0.06u
MNC1_3 N1 A0 VSS VPW NCH W=0.49u L=0.06u
MPC1_3 INT A0 N_13 VNW PCH W=0.63u L=0.06u
MPC1 INT A0 N_15 VNW PCH W=0.63u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.49u L=0.06u
MPC2 N_15 A1 VDD VNW PCH W=0.63u L=0.06u
MNC2_4 N1 A1 VSS VPW NCH W=0.49u L=0.06u
MPB1 INT B0 VDD VNW PCH W=0.435u L=0.06u
MNB1_5 N_71 B0 N1 VPW NCH W=0.49u L=0.06u
MPA1_4 INT C0 VDD VNW PCH W=0.435u L=0.06u
MNA1_5 INT C0 N_71 VPW NCH W=0.49u L=0.06u
MNA1_3 INT C0 N_73 VPW NCH W=0.49u L=0.06u
MPA1_3 INT C0 VDD VNW PCH W=0.435u L=0.06u
MNB1_3 N1 B0 N_73 VPW NCH W=0.49u L=0.06u
MPB1_4 INT B0 VDD VNW PCH W=0.435u L=0.06u
MNB1_4 N1 B0 N_75 VPW NCH W=0.49u L=0.06u
MPB1_3 INT B0 VDD VNW PCH W=0.435u L=0.06u
MNA1_4 INT C0 N_75 VPW NCH W=0.49u L=0.06u
MPA1_2 INT C0 VDD VNW PCH W=0.435u L=0.06u
MNA1_2 INT C0 N_77 VPW NCH W=0.49u L=0.06u
MPA1 INT C0 VDD VNW PCH W=0.435u L=0.06u
MNB1_2 N1 B0 N_77 VPW NCH W=0.49u L=0.06u
MPB1_2 INT B0 VDD VNW PCH W=0.435u L=0.06u
MNB1 N_81 B0 N1 VPW NCH W=0.49u L=0.06u
MNA1 INT C0 N_81 VPW NCH W=0.49u L=0.06u
MNA1_6 N_79 C0 INT VPW NCH W=0.49u L=0.06u
MNB1_6 N1 B0 N_79 VPW NCH W=0.49u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108_6 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108_5 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_6 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_5 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_4 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OA211X6MA10TR

****
.SUBCKT OA21X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0
MNB2 N1 A1 VSS VPW NCH W=0.24u L=0.06u
MPB2_2 VDD A1 N_5 VNW PCH W=0.395u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.24u L=0.06u
MPB1_2 INT A0 N_5 VNW PCH W=0.395u L=0.06u
MPB1 INT A0 N_7 VNW PCH W=0.395u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.24u L=0.06u
MPB2 N_7 A1 VDD VNW PCH W=0.395u L=0.06u
MNB2_2 N1 A1 VSS VPW NCH W=0.24u L=0.06u
MPA108 INT B0 VDD VNW PCH W=0.39u L=0.06u
MNA106_2 INT B0 N1 VPW NCH W=0.24u L=0.06u
MNA106 INT B0 N1 VPW NCH W=0.24u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS OA21X1P4MA10TR

****
.SUBCKT OA21X2MA10TR VDD VSS VPW VNW Y A0 A1 B0
MNB2 N1 A1 VSS VPW NCH W=0.335u L=0.06u
MPB2_2 VDD A1 N_5 VNW PCH W=0.555u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.335u L=0.06u
MPB1_2 INT A0 N_5 VNW PCH W=0.555u L=0.06u
MPB1 INT A0 N_7 VNW PCH W=0.555u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.335u L=0.06u
MPB2 N_7 A1 VDD VNW PCH W=0.555u L=0.06u
MNB2_2 N1 A1 VSS VPW NCH W=0.335u L=0.06u
MPA108 INT B0 VDD VNW PCH W=0.55u L=0.06u
MNA106_2 INT B0 N1 VPW NCH W=0.335u L=0.06u
MNA106 INT B0 N1 VPW NCH W=0.335u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OA21X2MA10TR

****
.SUBCKT OA21X3MA10TR VDD VSS VPW VNW Y A0 A1 B0
MPB1_2 INT A0 N_5 VNW PCH W=0.54u L=0.06u
MPB2_2 VDD A1 N_5 VNW PCH W=0.54u L=0.06u
MNB2_2 N1 A1 VSS VPW NCH W=0.495u L=0.06u
MPB2_3 VDD A1 N_7 VNW PCH W=0.54u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.495u L=0.06u
MPB1_3 INT A0 N_7 VNW PCH W=0.54u L=0.06u
MPB1 INT A0 N_9 VNW PCH W=0.54u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.495u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.495u L=0.06u
MPB2 N_9 A1 VDD VNW PCH W=0.54u L=0.06u
MNA106 INT B0 N1 VPW NCH W=0.495u L=0.06u
MPA108_2 INT B0 VDD VNW PCH W=0.405u L=0.06u
MNA106_2 INT B0 N1 VPW NCH W=0.495u L=0.06u
MPA108 INT B0 VDD VNW PCH W=0.405u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OA21X3MA10TR

****
.SUBCKT OA21X4MA10TR VDD VSS VPW VNW Y A0 A1 B0
MNB1_3 N1 A0 VSS VPW NCH W=0.425u L=0.06u
MPB1_3 INT A0 N_5 VNW PCH W=0.7u L=0.06u
MNB2_3 N1 A1 VSS VPW NCH W=0.425u L=0.06u
MPB2_3 VDD A1 N_5 VNW PCH W=0.7u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.425u L=0.06u
MPB2 VDD A1 N_7 VNW PCH W=0.7u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.425u L=0.06u
MPB1 INT A0 N_7 VNW PCH W=0.7u L=0.06u
MPB1_2 INT A0 N_3 VNW PCH W=0.7u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.425u L=0.06u
MNB2_2 N1 A1 VSS VPW NCH W=0.425u L=0.06u
MPB2_2 N_3 A1 VDD VNW PCH W=0.7u L=0.06u
MNA106_2 INT B0 N1 VPW NCH W=0.425u L=0.06u
MPA108_2 INT B0 VDD VNW PCH W=0.52u L=0.06u
MPA108 INT B0 VDD VNW PCH W=0.52u L=0.06u
MNA106 INT B0 N1 VPW NCH W=0.425u L=0.06u
MNA106_3 INT B0 N1 VPW NCH W=0.425u L=0.06u
MNA1_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA1_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1_4 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OA21X4MA10TR

****
.SUBCKT OA22X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1
MNB2_2 N1 A1 VSS VPW NCH W=0.27u L=0.06u
MPB2_2 VDD A1 N_8 VNW PCH W=0.4u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.27u L=0.06u
MPB1_2 INT A0 N_8 VNW PCH W=0.4u L=0.06u
MPB1 INT A0 N_10 VNW PCH W=0.4u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.27u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.27u L=0.06u
MPB2 N_10 A1 VDD VNW PCH W=0.4u L=0.06u
MNA2_2 INT B1 N1 VPW NCH W=0.27u L=0.06u
MPA2 VDD B1 N_12 VNW PCH W=0.4u L=0.06u
MNA1_2 INT B0 N1 VPW NCH W=0.27u L=0.06u
MPA1 INT B0 N_12 VNW PCH W=0.4u L=0.06u
MPA1_2 INT B0 N_6 VNW PCH W=0.4u L=0.06u
MNA1 INT B0 N1 VPW NCH W=0.27u L=0.06u
MPA2_2 N_6 B1 VDD VNW PCH W=0.4u L=0.06u
MNA2 INT B1 N1 VPW NCH W=0.27u L=0.06u
MNA108_2 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1010_2 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS OA22X1P4MA10TR

****
.SUBCKT OA22X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1
MNB2_2 N1 A1 VSS VPW NCH W=0.37u L=0.06u
MPB2_2 VDD A1 N_5 VNW PCH W=0.55u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.37u L=0.06u
MPB1_2 INT A0 N_5 VNW PCH W=0.55u L=0.06u
MPB1 INT A0 N_7 VNW PCH W=0.55u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.37u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.37u L=0.06u
MPB2 N_7 A1 VDD VNW PCH W=0.55u L=0.06u
MNA2_2 INT B1 N1 VPW NCH W=0.37u L=0.06u
MPA2_2 VDD B1 N_9 VNW PCH W=0.55u L=0.06u
MNA1_2 INT B0 N1 VPW NCH W=0.37u L=0.06u
MPA1_2 INT B0 N_9 VNW PCH W=0.55u L=0.06u
MPA1 INT B0 N_3 VNW PCH W=0.55u L=0.06u
MNA1 INT B0 N1 VPW NCH W=0.37u L=0.06u
MPA2 N_3 B1 VDD VNW PCH W=0.55u L=0.06u
MNA2 INT B1 N1 VPW NCH W=0.37u L=0.06u
MNA108_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA108 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1010 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OA22X2MA10TR

****
.SUBCKT OAI211X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MNC2 N1 A1 VSS VPW NCH W=0.405u L=0.06u
MPC2 VDD A1 N_5 VNW PCH W=0.465u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.405u L=0.06u
MPC1 Y A0 N_5 VNW PCH W=0.465u L=0.06u
MPC1_2 Y A0 N_7 VNW PCH W=0.465u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.405u L=0.06u
MPC2_2 N_7 A1 VDD VNW PCH W=0.465u L=0.06u
MNC2_2 N1 A1 VSS VPW NCH W=0.405u L=0.06u
MNB1_2 N1 B0 N_23 VPW NCH W=0.405u L=0.06u
MPB1 Y B0 VDD VNW PCH W=0.5u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.5u L=0.06u
MNA1_2 Y C0 N_23 VPW NCH W=0.405u L=0.06u
MNA1 N_17 C0 Y VPW NCH W=0.405u L=0.06u
MNB1 N1 B0 N_17 VPW NCH W=0.405u L=0.06u
.ENDS OAI211X1P4MA10TR

****
.SUBCKT OAI211X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MNC2_2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2 VDD A1 N_5 VNW PCH W=0.665u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1 Y A0 N_5 VNW PCH W=0.665u L=0.06u
MPC1_2 Y A0 N_8 VNW PCH W=0.665u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC2_2 N_8 A1 VDD VNW PCH W=0.665u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MNB1 N_27 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1_2 Y B0 VDD VNW PCH W=0.36u L=0.06u
MNA1 Y C0 N_27 VPW NCH W=0.58u L=0.06u
MPA1_2 Y C0 VDD VNW PCH W=0.36u L=0.06u
MNA1_2 Y C0 N_21 VPW NCH W=0.58u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.36u L=0.06u
MNB1_2 N_21 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1 Y B0 VDD VNW PCH W=0.36u L=0.06u
.ENDS OAI211X2MA10TR

****
.SUBCKT OAI211X3MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MNC1_2 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_3 Y A0 N_5 VNW PCH W=0.665u L=0.06u
MNC2_3 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_3 VDD A1 N_5 VNW PCH W=0.665u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_2 VDD A1 N_7 VNW PCH W=0.665u L=0.06u
MNC1_3 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_2 Y A0 N_7 VNW PCH W=0.665u L=0.06u
MPC1 Y A0 N_9 VNW PCH W=0.665u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC2 N_9 A1 VDD VNW PCH W=0.665u L=0.06u
MNC2_2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MNB1_2 N1 B0 N_33 VPW NCH W=0.58u L=0.06u
MPB1_2 Y B0 VDD VNW PCH W=0.54u L=0.06u
MNA1_2 Y C0 N_33 VPW NCH W=0.58u L=0.06u
MPA1_2 Y C0 VDD VNW PCH W=0.54u L=0.06u
MNA1 Y C0 N_35 VPW NCH W=0.58u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.54u L=0.06u
MNB1 N1 B0 N_35 VPW NCH W=0.58u L=0.06u
MPB1 Y B0 VDD VNW PCH W=0.54u L=0.06u
MNB1_3 N_25 B0 N1 VPW NCH W=0.58u L=0.06u
MNA1_3 Y C0 N_25 VPW NCH W=0.58u L=0.06u
.ENDS OAI211X3MA10TR

****
.SUBCKT OAI211X4MA10TR VDD VSS VPW VNW Y A0 A1 B0 C0
MNC2_4 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_3 VDD A1 N_5 VNW PCH W=0.665u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_3 Y A0 N_5 VNW PCH W=0.665u L=0.06u
MPC1_4 Y A0 N_7 VNW PCH W=0.665u L=0.06u
MNC1_4 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2_3 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_4 VDD A1 N_7 VNW PCH W=0.665u L=0.06u
MNC2_2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2 VDD A1 N_9 VNW PCH W=0.665u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1 Y A0 N_9 VNW PCH W=0.665u L=0.06u
MPC1_2 Y A0 N_12 VNW PCH W=0.665u L=0.06u
MNC1_3 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC2_2 N_12 A1 VDD VNW PCH W=0.665u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPB1_3 Y B0 VDD VNW PCH W=0.48u L=0.06u
MNB1_3 N1 B0 N_43 VPW NCH W=0.58u L=0.06u
MPA1_3 Y C0 VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y C0 N_43 VPW NCH W=0.58u L=0.06u
MNA1_4 Y C0 N_45 VPW NCH W=0.58u L=0.06u
MPA1_2 Y C0 VDD VNW PCH W=0.48u L=0.06u
MNB1_4 N1 B0 N_45 VPW NCH W=0.58u L=0.06u
MPB1_2 Y B0 VDD VNW PCH W=0.48u L=0.06u
MNB1 N1 B0 N_47 VPW NCH W=0.58u L=0.06u
MPB1 Y B0 VDD VNW PCH W=0.48u L=0.06u
MNA1 Y C0 N_47 VPW NCH W=0.58u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.48u L=0.06u
MNA1_2 N_33 C0 Y VPW NCH W=0.58u L=0.06u
MNB1_2 N1 B0 N_33 VPW NCH W=0.58u L=0.06u
.ENDS OAI211X4MA10TR

****
.SUBCKT OAI21X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0
MNB2_2 N1 A1 VSS VPW NCH W=0.32u L=0.06u
MPB2 VDD A1 N_5 VNW PCH W=0.49u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MPB1 Y A0 N_5 VNW PCH W=0.49u L=0.06u
MPB1_2 Y A0 N_8 VNW PCH W=0.49u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.32u L=0.06u
MPB2_2 N_8 A1 VDD VNW PCH W=0.49u L=0.06u
MNA1 Y B0 N1 VPW NCH W=0.32u L=0.06u
MPA1 Y B0 VDD VNW PCH W=0.265u L=0.06u
MNA1_2 Y B0 N1 VPW NCH W=0.32u L=0.06u
MPA1_2 Y B0 VDD VNW PCH W=0.265u L=0.06u
.ENDS OAI21X1P4MA10TR

****
.SUBCKT OAI21X2MA10TR VDD VSS VPW VNW Y A0 A1 B0
MNB2_2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPB2 VDD A1 N_5 VNW PCH W=0.7u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MPB1 Y A0 N_5 VNW PCH W=0.7u L=0.06u
MPB1_2 Y A0 N_3 VNW PCH W=0.7u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPB2_2 N_3 A1 VDD VNW PCH W=0.7u L=0.06u
MNA1 Y B0 N1 VPW NCH W=0.455u L=0.06u
MPA1_2 Y B0 VDD VNW PCH W=0.38u L=0.06u
MNA1_2 Y B0 N1 VPW NCH W=0.455u L=0.06u
MPA1 Y B0 VDD VNW PCH W=0.38u L=0.06u
.ENDS OAI21X2MA10TR

****
.SUBCKT OAI21X3MA10TR VDD VSS VPW VNW Y A0 A1 B0
MNB1_3 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MPB1 Y A0 N_5 VNW PCH W=0.7u L=0.06u
MNB2_3 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPB2 VDD A1 N_5 VNW PCH W=0.7u L=0.06u
MNB2_2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPB2_3 VDD A1 N_7 VNW PCH W=0.7u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MPB1_3 Y A0 N_7 VNW PCH W=0.7u L=0.06u
MPB1_2 Y A0 N_10 VNW PCH W=0.7u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPB2_2 N_10 A1 VDD VNW PCH W=0.7u L=0.06u
MNA1 Y B0 N1 VPW NCH W=0.455u L=0.06u
MPA1 Y B0 VDD VNW PCH W=0.57u L=0.06u
MPA1_2 Y B0 VDD VNW PCH W=0.57u L=0.06u
MNA1_3 Y B0 N1 VPW NCH W=0.455u L=0.06u
MNA1_2 Y B0 N1 VPW NCH W=0.455u L=0.06u
.ENDS OAI21X3MA10TR

****
.SUBCKT OAI221X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0
MNC2_2 N1 A1 VSS VPW NCH W=0.405u L=0.06u
MPC2_2 VDD A1 N_5 VNW PCH W=0.465u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.405u L=0.06u
MPC1_2 Y A0 N_5 VNW PCH W=0.465u L=0.06u
MPC1 Y A0 N_3 VNW PCH W=0.465u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.405u L=0.06u
MPC2 N_3 A1 VDD VNW PCH W=0.465u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.405u L=0.06u
MPB2 VDD B1 N_10 VNW PCH W=0.465u L=0.06u
MNB2_2 N2 B1 N1 VPW NCH W=0.405u L=0.06u
MPB1 Y B0 N_10 VNW PCH W=0.465u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.405u L=0.06u
MPB1_2 Y B0 N_13 VNW PCH W=0.465u L=0.06u
MNB1_2 N2 B0 N1 VPW NCH W=0.405u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.405u L=0.06u
MPB2_2 N_13 B1 VDD VNW PCH W=0.465u L=0.06u
MNA1 Y C0 N2 VPW NCH W=0.405u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.25u L=0.06u
MNA1_2 Y C0 N2 VPW NCH W=0.405u L=0.06u
MPA1_2 Y C0 VDD VNW PCH W=0.25u L=0.06u
.ENDS OAI221X1P4MA10TR

****
.SUBCKT OAI221X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0
MNC2_2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_2 VDD A1 N_5 VNW PCH W=0.665u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_2 Y A0 N_5 VNW PCH W=0.665u L=0.06u
MPC1 Y A0 N_3 VNW PCH W=0.665u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC2 N_3 A1 VDD VNW PCH W=0.665u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPB2 VDD B1 N_10 VNW PCH W=0.665u L=0.06u
MNB2_2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB1 Y B0 N_10 VNW PCH W=0.665u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1_2 Y B0 N_8 VNW PCH W=0.665u L=0.06u
MNB1_2 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2_2 N_8 B1 VDD VNW PCH W=0.665u L=0.06u
MNA1 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.36u L=0.06u
MNA1_2 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA1_2 Y C0 VDD VNW PCH W=0.36u L=0.06u
.ENDS OAI221X2MA10TR

****
.SUBCKT OAI221X3MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0
MNC2_2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_3 VDD A1 N_8 VNW PCH W=0.665u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_3 Y A0 N_8 VNW PCH W=0.665u L=0.06u
MPC1 Y A0 N_10 VNW PCH W=0.665u L=0.06u
MNC1_3 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2_3 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2 VDD A1 N_10 VNW PCH W=0.665u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_2 VDD A1 N_12 VNW PCH W=0.665u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_2 N_12 A0 Y VNW PCH W=0.665u L=0.06u
MPB1_3 Y B0 N_14 VNW PCH W=0.665u L=0.06u
MNB1_2 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MNB2_2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2_3 VDD B1 N_14 VNW PCH W=0.665u L=0.06u
MNB2_3 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2_2 VDD B1 N_16 VNW PCH W=0.665u L=0.06u
MNB1_3 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1_2 Y B0 N_16 VNW PCH W=0.665u L=0.06u
MPB1 Y B0 N_6 VNW PCH W=0.665u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB2 N_6 B1 VDD VNW PCH W=0.665u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MNA1 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA1_2 Y C0 VDD VNW PCH W=0.54u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.54u L=0.06u
MNA1_3 Y C0 N2 VPW NCH W=0.58u L=0.06u
MNA1_2 Y C0 N2 VPW NCH W=0.58u L=0.06u
.ENDS OAI221X3MA10TR

****
.SUBCKT OAI221X4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0
MNC2_2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_4 VDD A1 N_5 VNW PCH W=0.665u L=0.06u
MNC1_4 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_4 Y A0 N_5 VNW PCH W=0.665u L=0.06u
MPC1_2 Y A0 N_7 VNW PCH W=0.665u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_2 VDD A1 N_7 VNW PCH W=0.665u L=0.06u
MNC2_4 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_3 VDD A1 N_9 VNW PCH W=0.665u L=0.06u
MNC1_3 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_3 Y A0 N_9 VNW PCH W=0.665u L=0.06u
MPC1 Y A0 N_3 VNW PCH W=0.665u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC2 N_3 A1 VDD VNW PCH W=0.665u L=0.06u
MNC2_3 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPB2_4 VDD B1 N_14 VNW PCH W=0.665u L=0.06u
MNB2_2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB1_4 Y B0 N_14 VNW PCH W=0.665u L=0.06u
MNB1_4 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1_2 Y B0 N_16 VNW PCH W=0.665u L=0.06u
MNB1_2 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2_2 VDD B1 N_16 VNW PCH W=0.665u L=0.06u
MPB2_3 VDD B1 N_18 VNW PCH W=0.665u L=0.06u
MNB2_4 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB1_3 Y B0 N_18 VNW PCH W=0.665u L=0.06u
MNB1_3 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1 Y B0 N_12 VNW PCH W=0.665u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MNB2_3 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2 N_12 B1 VDD VNW PCH W=0.665u L=0.06u
MNA1_4 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA1_3 Y C0 VDD VNW PCH W=0.48u L=0.06u
MNA1_3 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA1_2 Y C0 VDD VNW PCH W=0.48u L=0.06u
MPA1 Y C0 VDD VNW PCH W=0.48u L=0.06u
MNA1_2 Y C0 N2 VPW NCH W=0.58u L=0.06u
MNA1 Y C0 N2 VPW NCH W=0.58u L=0.06u
.ENDS OAI221X4MA10TR

****
.SUBCKT OAI222X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0 C1
MNC2_2 N1 A1 VSS VPW NCH W=0.405u L=0.06u
MPC2 VDD A1 N_5 VNW PCH W=0.465u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.405u L=0.06u
MPC1 Y A0 N_5 VNW PCH W=0.465u L=0.06u
MPC1_2 Y A0 N_7 VNW PCH W=0.465u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.405u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.405u L=0.06u
MPC2_2 N_7 A1 VDD VNW PCH W=0.465u L=0.06u
MNB2_2 N2 B1 N1 VPW NCH W=0.405u L=0.06u
MPB2 VDD B1 N_9 VNW PCH W=0.465u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.405u L=0.06u
MPB1 Y B0 N_9 VNW PCH W=0.465u L=0.06u
MPB1_2 Y B0 N_3 VNW PCH W=0.465u L=0.06u
MNB1_2 N2 B0 N1 VPW NCH W=0.405u L=0.06u
MPB2_2 N_3 B1 VDD VNW PCH W=0.465u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.405u L=0.06u
MNA2_2 Y C1 N2 VPW NCH W=0.405u L=0.06u
MPA2_2 VDD C1 N_14 VNW PCH W=0.465u L=0.06u
MNA1_2 Y C0 N2 VPW NCH W=0.405u L=0.06u
MPA1_2 Y C0 N_14 VNW PCH W=0.465u L=0.06u
MPA1 Y C0 N_12 VNW PCH W=0.465u L=0.06u
MNA1 Y C0 N2 VPW NCH W=0.405u L=0.06u
MPA2 N_12 C1 VDD VNW PCH W=0.465u L=0.06u
MNA2 Y C1 N2 VPW NCH W=0.405u L=0.06u
.ENDS OAI222X1P4MA10TR

****
.SUBCKT OAI222X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0 C1
MNC2_2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2 VDD A1 N_5 VNW PCH W=0.665u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1 Y A0 N_5 VNW PCH W=0.665u L=0.06u
MPC1_2 Y A0 N_7 VNW PCH W=0.665u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_2 N_7 A1 VDD VNW PCH W=0.665u L=0.06u
MNB2_2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2 VDD B1 N_9 VNW PCH W=0.665u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1 Y B0 N_9 VNW PCH W=0.665u L=0.06u
MPB1_2 Y B0 N_3 VNW PCH W=0.665u L=0.06u
MNB1_2 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB2_2 N_3 B1 VDD VNW PCH W=0.665u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MNA2_2 Y C1 N2 VPW NCH W=0.58u L=0.06u
MPA2_2 VDD C1 N_14 VNW PCH W=0.665u L=0.06u
MNA1_2 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA1_2 Y C0 N_14 VNW PCH W=0.665u L=0.06u
MPA1 Y C0 N_12 VNW PCH W=0.665u L=0.06u
MNA1 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA2 N_12 C1 VDD VNW PCH W=0.665u L=0.06u
MNA2 Y C1 N2 VPW NCH W=0.58u L=0.06u
.ENDS OAI222X2MA10TR

****
.SUBCKT OAI222X3MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0 C1
MNC2_3 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_3 VDD A1 N_5 VNW PCH W=0.665u L=0.06u
MNC1_3 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_3 Y A0 N_5 VNW PCH W=0.665u L=0.06u
MPC1_2 Y A0 N_7 VNW PCH W=0.665u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2_2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_2 VDD A1 N_7 VNW PCH W=0.665u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2 VDD A1 N_9 VNW PCH W=0.665u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1 N_9 A0 Y VNW PCH W=0.665u L=0.06u
MPB1_3 Y B0 N_11 VNW PCH W=0.665u L=0.06u
MNB1_3 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MNB2_3 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2_3 VDD B1 N_11 VNW PCH W=0.665u L=0.06u
MNB2_2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2_2 VDD B1 N_13 VNW PCH W=0.665u L=0.06u
MNB1_2 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1_2 Y B0 N_13 VNW PCH W=0.665u L=0.06u
MPB1 Y B0 N_3 VNW PCH W=0.665u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB2 N_3 B1 VDD VNW PCH W=0.665u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPA1_3 Y C0 N_18 VNW PCH W=0.665u L=0.06u
MNA1_3 Y C0 N2 VPW NCH W=0.58u L=0.06u
MNA2_3 Y C1 N2 VPW NCH W=0.58u L=0.06u
MPA2_3 VDD C1 N_18 VNW PCH W=0.665u L=0.06u
MNA2_2 Y C1 N2 VPW NCH W=0.58u L=0.06u
MPA2_2 VDD C1 N_20 VNW PCH W=0.665u L=0.06u
MNA1_2 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA1_2 Y C0 N_20 VNW PCH W=0.665u L=0.06u
MPA1 Y C0 N_16 VNW PCH W=0.665u L=0.06u
MNA1 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA2 N_16 C1 VDD VNW PCH W=0.665u L=0.06u
MNA2 Y C1 N2 VPW NCH W=0.58u L=0.06u
.ENDS OAI222X3MA10TR

****
.SUBCKT OAI222X4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1 C0 C1
MNC2_4 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_4 VDD A1 N_113 VNW PCH W=0.665u L=0.06u
MNC1_3 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1_4 Y A0 N_113 VNW PCH W=0.665u L=0.06u
MPC1_3 Y A0 N_115 VNW PCH W=0.665u L=0.06u
MNC1_2 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2_3 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_3 VDD A1 N_115 VNW PCH W=0.665u L=0.06u
MNC2_2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2 VDD A1 N_117 VNW PCH W=0.665u L=0.06u
MNC1 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MPC1 Y A0 N_117 VNW PCH W=0.665u L=0.06u
MPC1_2 Y A0 N_119 VNW PCH W=0.665u L=0.06u
MNC1_4 N1 A0 VSS VPW NCH W=0.58u L=0.06u
MNC2 N1 A1 VSS VPW NCH W=0.58u L=0.06u
MPC2_2 N_119 A1 VDD VNW PCH W=0.665u L=0.06u
MNB2_3 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2_3 VDD B1 N_121 VNW PCH W=0.665u L=0.06u
MNB1_4 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1_3 Y B0 N_121 VNW PCH W=0.665u L=0.06u
MPB1_4 Y B0 N_123 VNW PCH W=0.665u L=0.06u
MNB1_3 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MNB2_2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2_4 VDD B1 N_123 VNW PCH W=0.665u L=0.06u
MNB2 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MPB2 VDD B1 N_125 VNW PCH W=0.665u L=0.06u
MNB1_2 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB1 Y B0 N_125 VNW PCH W=0.665u L=0.06u
MPB1_2 Y B0 N_111 VNW PCH W=0.665u L=0.06u
MNB1 N2 B0 N1 VPW NCH W=0.58u L=0.06u
MPB2_2 N_111 B1 VDD VNW PCH W=0.665u L=0.06u
MNB2_4 N2 B1 N1 VPW NCH W=0.58u L=0.06u
MNA2 Y C1 N2 VPW NCH W=0.58u L=0.06u
MPA2_4 VDD C1 N_130 VNW PCH W=0.665u L=0.06u
MNA1_4 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA1_4 Y C0 N_130 VNW PCH W=0.665u L=0.06u
MPA1 Y C0 N_132 VNW PCH W=0.665u L=0.06u
MNA1_3 Y C0 N2 VPW NCH W=0.58u L=0.06u
MNA2_4 Y C1 N2 VPW NCH W=0.58u L=0.06u
MPA2 VDD C1 N_132 VNW PCH W=0.665u L=0.06u
MNA2_3 Y C1 N2 VPW NCH W=0.58u L=0.06u
MPA2_3 VDD C1 N_134 VNW PCH W=0.665u L=0.06u
MNA1_2 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA1_3 Y C0 N_134 VNW PCH W=0.665u L=0.06u
MPA1_2 Y C0 N_128 VNW PCH W=0.665u L=0.06u
MNA1 Y C0 N2 VPW NCH W=0.58u L=0.06u
MPA2_2 N_128 C1 VDD VNW PCH W=0.665u L=0.06u
MNA2_2 Y C1 N2 VPW NCH W=0.58u L=0.06u
.ENDS OAI222X4MA10TR

****
.SUBCKT OAI22X1P4MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1
MNB2_2 N1 A1 VSS VPW NCH W=0.32u L=0.06u
MPB2 VDD A1 N_5 VNW PCH W=0.49u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MPB1 Y A0 N_5 VNW PCH W=0.49u L=0.06u
MPB1_2 Y A0 N_7 VNW PCH W=0.49u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.32u L=0.06u
MPB2_2 N_7 A1 VDD VNW PCH W=0.49u L=0.06u
MNA2_2 Y B1 N1 VPW NCH W=0.32u L=0.06u
MPA2 VDD B1 N_9 VNW PCH W=0.49u L=0.06u
MNA1_2 Y B0 N1 VPW NCH W=0.32u L=0.06u
MPA1 Y B0 N_9 VNW PCH W=0.49u L=0.06u
MPA1_2 Y B0 N_3 VNW PCH W=0.49u L=0.06u
MNA1 Y B0 N1 VPW NCH W=0.32u L=0.06u
MPA2_2 N_3 B1 VDD VNW PCH W=0.49u L=0.06u
MNA2 Y B1 N1 VPW NCH W=0.32u L=0.06u
.ENDS OAI22X1P4MA10TR

****
.SUBCKT OAI22X2MA10TR VDD VSS VPW VNW Y A0 A1 B0 B1
MNB2_2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPB2 VDD A1 N_5 VNW PCH W=0.7u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MPB1 Y A0 N_5 VNW PCH W=0.7u L=0.06u
MPB1_2 Y A0 N_7 VNW PCH W=0.7u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MNB2 N1 A1 VSS VPW NCH W=0.455u L=0.06u
MPB2_2 N_7 A1 VDD VNW PCH W=0.7u L=0.06u
MNA2_2 Y B1 N1 VPW NCH W=0.455u L=0.06u
MPA2 VDD B1 N_9 VNW PCH W=0.7u L=0.06u
MNA1_2 Y B0 N1 VPW NCH W=0.455u L=0.06u
MPA1 Y B0 N_9 VNW PCH W=0.7u L=0.06u
MPA1_2 Y B0 N_3 VNW PCH W=0.7u L=0.06u
MNA1 Y B0 N1 VPW NCH W=0.455u L=0.06u
MPA2_2 N_3 B1 VDD VNW PCH W=0.7u L=0.06u
MNA2 Y B1 N1 VPW NCH W=0.455u L=0.06u
.ENDS OAI22X2MA10TR

****
.SUBCKT OAI2XB1X1P4MA10TR VDD VSS VPW VNW Y A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.22u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.295u L=0.06u
MNB2_2 N1 INT VSS VPW NCH W=0.32u L=0.06u
MPB2 VDD INT N_7 VNW PCH W=0.49u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MPB1 Y A0 N_7 VNW PCH W=0.49u L=0.06u
MPB1_2 Y A0 N_10 VNW PCH W=0.49u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.32u L=0.06u
MNB2 N1 INT VSS VPW NCH W=0.32u L=0.06u
MPB2_2 N_10 INT VDD VNW PCH W=0.49u L=0.06u
MNA106 Y B0 N1 VPW NCH W=0.32u L=0.06u
MPA108 Y B0 VDD VNW PCH W=0.265u L=0.06u
MNA106_2 Y B0 N1 VPW NCH W=0.32u L=0.06u
MPA108_2 Y B0 VDD VNW PCH W=0.265u L=0.06u
.ENDS OAI2XB1X1P4MA10TR

****
.SUBCKT OAI2XB1X2MA10TR VDD VSS VPW VNW Y A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.295u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.39u L=0.06u
MNB2_2 N1 INT VSS VPW NCH W=0.455u L=0.06u
MPB2 VDD INT N_5 VNW PCH W=0.7u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MPB1 Y A0 N_5 VNW PCH W=0.7u L=0.06u
MPB1_2 Y A0 N_3 VNW PCH W=0.7u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MNB2 N1 INT VSS VPW NCH W=0.455u L=0.06u
MPB2_2 N_3 INT VDD VNW PCH W=0.7u L=0.06u
MNA106 Y B0 N1 VPW NCH W=0.455u L=0.06u
MPA108_2 Y B0 VDD VNW PCH W=0.38u L=0.06u
MNA106_2 Y B0 N1 VPW NCH W=0.455u L=0.06u
MPA108 Y B0 VDD VNW PCH W=0.38u L=0.06u
.ENDS OAI2XB1X2MA10TR

****
.SUBCKT OAI2XB1X3MA10TR VDD VSS VPW VNW Y A0 A1N B0
MNA1 INT A1N VSS VPW NCH W=0.455u L=0.06u
MPA1 INT A1N VDD VNW PCH W=0.6u L=0.06u
MNB1_3 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MPB1 Y A0 N_7 VNW PCH W=0.7u L=0.06u
MNB2_3 N1 INT VSS VPW NCH W=0.455u L=0.06u
MPB2 VDD INT N_7 VNW PCH W=0.7u L=0.06u
MNB2_2 N1 INT VSS VPW NCH W=0.455u L=0.06u
MPB2_3 VDD INT N_9 VNW PCH W=0.7u L=0.06u
MNB1_2 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MPB1_3 Y A0 N_9 VNW PCH W=0.7u L=0.06u
MPB1_2 Y A0 N_12 VNW PCH W=0.7u L=0.06u
MNB1 N1 A0 VSS VPW NCH W=0.455u L=0.06u
MNB2 N1 INT VSS VPW NCH W=0.455u L=0.06u
MPB2_2 N_12 INT VDD VNW PCH W=0.7u L=0.06u
MNA106 Y B0 N1 VPW NCH W=0.455u L=0.06u
MPA108 Y B0 VDD VNW PCH W=0.57u L=0.06u
MPA108_2 Y B0 VDD VNW PCH W=0.57u L=0.06u
MNA106_3 Y B0 N1 VPW NCH W=0.455u L=0.06u
MNA106_2 Y B0 N1 VPW NCH W=0.455u L=0.06u
.ENDS OAI2XB1X3MA10TR

****
.SUBCKT OR2X11MA10TR VDD VSS VPW VNW Y A B
MNA2_6 INT B VSS VPW NCH W=0.27u L=0.06u
MPA2_2 VDD B N_5 VNW PCH W=0.685u L=0.06u
MNA1_8 INT A VSS VPW NCH W=0.27u L=0.06u
MPA1_2 INT A N_5 VNW PCH W=0.685u L=0.06u
MPA1 INT A N_7 VNW PCH W=0.685u L=0.06u
MNA1_6 INT A VSS VPW NCH W=0.27u L=0.06u
MNA2_3 INT B VSS VPW NCH W=0.27u L=0.06u
MPA2 VDD B N_7 VNW PCH W=0.685u L=0.06u
MNA2_2 INT B VSS VPW NCH W=0.27u L=0.06u
MPA2_7 VDD B N_9 VNW PCH W=0.685u L=0.06u
MNA1_4 INT A VSS VPW NCH W=0.27u L=0.06u
MPA1_7 INT A N_9 VNW PCH W=0.685u L=0.06u
MPA1_5 INT A N_11 VNW PCH W=0.685u L=0.06u
MNA1_3 INT A VSS VPW NCH W=0.27u L=0.06u
MNA2_8 INT B VSS VPW NCH W=0.27u L=0.06u
MPA2_5 VDD B N_11 VNW PCH W=0.685u L=0.06u
MNA2_7 INT B VSS VPW NCH W=0.27u L=0.06u
MPA2_8 VDD B N_13 VNW PCH W=0.685u L=0.06u
MNA1_2 INT A VSS VPW NCH W=0.27u L=0.06u
MPA1_8 INT A N_13 VNW PCH W=0.685u L=0.06u
MPA1_6 INT A N_15 VNW PCH W=0.685u L=0.06u
MNA1 INT A VSS VPW NCH W=0.27u L=0.06u
MNA2_5 INT B VSS VPW NCH W=0.27u L=0.06u
MPA2_6 VDD B N_15 VNW PCH W=0.685u L=0.06u
MPA2_3 VDD B N_17 VNW PCH W=0.685u L=0.06u
MNA2_4 INT B VSS VPW NCH W=0.27u L=0.06u
MPA1_3 INT A N_17 VNW PCH W=0.685u L=0.06u
MNA1_7 INT A VSS VPW NCH W=0.27u L=0.06u
MPA1_4 INT A N_19 VNW PCH W=0.685u L=0.06u
MNA1_5 INT A VSS VPW NCH W=0.27u L=0.06u
MNA2 INT B VSS VPW NCH W=0.27u L=0.06u
MPA2_4 N_19 B VDD VNW PCH W=0.685u L=0.06u
MNA104_10 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_5 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_8 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_6 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_10 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_8 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_7 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_11 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_6 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_9 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_7 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_5 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_11 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_9 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OR2X11MA10TR

****
.SUBCKT OR2X1P4MA10TR VDD VSS VPW VNW Y A B
MNA2_2 INT B VSS VPW NCH W=0.15u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.38u L=0.06u
MNA1_2 INT A VSS VPW NCH W=0.15u L=0.06u
MPA1 INT A N_5 VNW PCH W=0.38u L=0.06u
MNA1 INT A VSS VPW NCH W=0.15u L=0.06u
MPA1_2 INT A N_7 VNW PCH W=0.38u L=0.06u
MNA2 INT B VSS VPW NCH W=0.15u L=0.06u
MPA2_2 N_7 B VDD VNW PCH W=0.38u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS OR2X1P4MA10TR

****
.SUBCKT XOR2X1P4MA10TR VDD VSS VPW VNW Y A B
MNA108 NIN1 A VSS VPW NCH W=0.53u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.7u L=0.06u
MNA1_2 NIN2 B VSS VPW NCH W=0.33u L=0.06u
MPA1_2 NIN2 B VDD VNW PCH W=0.49u L=0.06u
MNA1 NIN2 B VSS VPW NCH W=0.33u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.49u L=0.06u
MNOE_2 Y A NIN2 VPW NCH W=0.33u L=0.06u
MPOEN Y NIN1 NIN2 VNW PCH W=0.33u L=0.06u
MNOE Y A NIN2 VPW NCH W=0.33u L=0.06u
MPOEN_2 Y NIN1 NIN2 VNW PCH W=0.33u L=0.06u
MNOE02_2 Y NIN1 BIN2 VPW NCH W=0.33u L=0.06u
MPOEN04 Y A BIN2 VNW PCH W=0.33u L=0.06u
MNOE02 Y NIN1 BIN2 VPW NCH W=0.33u L=0.06u
MPOEN04_2 Y A BIN2 VNW PCH W=0.33u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.33u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.66u L=0.06u
MNA1012_2 BIN2 NIN2 VSS VPW NCH W=0.33u L=0.06u
.ENDS XOR2X1P4MA10TR

****
.SUBCKT OR2X2MA10TR VDD VSS VPW VNW Y A B
MNA2_2 INT B VSS VPW NCH W=0.195u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.495u L=0.06u
MNA1_2 INT A VSS VPW NCH W=0.195u L=0.06u
MPA1 INT A N_5 VNW PCH W=0.495u L=0.06u
MNA1 INT A VSS VPW NCH W=0.195u L=0.06u
MPA1_2 INT A N_7 VNW PCH W=0.495u L=0.06u
MNA2 INT B VSS VPW NCH W=0.195u L=0.06u
MPA2_2 N_7 B VDD VNW PCH W=0.495u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OR2X2MA10TR

****
.SUBCKT XOR2X2MA10TR VDD VSS VPW VNW Y A B
MNA108_2 NIN1 A VSS VPW NCH W=0.33u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.44u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.33u L=0.06u
MPA1010_2 NIN1 A VDD VNW PCH W=0.44u L=0.06u
MNA1_2 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_2 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNOE Y A NIN2 VPW NCH W=0.47u L=0.06u
MPOEN Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MNOE_2 Y A NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_2 Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MNOE02_2 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_2 Y A BIN2 VNW PCH W=0.47u L=0.06u
MNOE02 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04 Y A BIN2 VNW PCH W=0.47u L=0.06u
MNA1012_2 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_2 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
.ENDS XOR2X2MA10TR

****
.SUBCKT OR2X3MA10TR VDD VSS VPW VNW Y A B
MNA1_3 INT A VSS VPW NCH W=0.195u L=0.06u
MPA1_2 INT A N_5 VNW PCH W=0.5u L=0.06u
MNA2_3 INT B VSS VPW NCH W=0.195u L=0.06u
MPA2_2 VDD B N_5 VNW PCH W=0.5u L=0.06u
MNA2_2 INT B VSS VPW NCH W=0.195u L=0.06u
MPA2 VDD B N_7 VNW PCH W=0.5u L=0.06u
MNA1_2 INT A VSS VPW NCH W=0.195u L=0.06u
MPA1 INT A N_7 VNW PCH W=0.5u L=0.06u
MPA1_3 INT A N_9 VNW PCH W=0.5u L=0.06u
MNA1 INT A VSS VPW NCH W=0.195u L=0.06u
MNA2 INT B VSS VPW NCH W=0.195u L=0.06u
MPA2_3 N_9 B VDD VNW PCH W=0.5u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OR2X3MA10TR

****
.SUBCKT XOR2X3MA10TR VDD VSS VPW VNW Y A B
MNA108 NIN1 A VSS VPW NCH W=0.485u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.645u L=0.06u
MNA108_2 NIN1 A VSS VPW NCH W=0.485u L=0.06u
MPA1010_2 NIN1 A VDD VNW PCH W=0.645u L=0.06u
MNA1 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_2 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_3 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_3 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNOE_2 Y A NIN2 VPW NCH W=0.47u L=0.06u
MPOEN Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MNOE Y A NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_3 Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MNOE_3 Y A NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_2 Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MNOE02_2 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04 Y A BIN2 VNW PCH W=0.47u L=0.06u
MNOE02 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_3 Y A BIN2 VNW PCH W=0.47u L=0.06u
MNOE02_3 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_2 Y A BIN2 VNW PCH W=0.47u L=0.06u
MNA1012_2 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_3 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MPA1014_2 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012_3 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
.ENDS XOR2X3MA10TR

****
.SUBCKT OR2X4MA10TR VDD VSS VPW VNW Y A B
MNA1_2 INT A VSS VPW NCH W=0.26u L=0.06u
MPA1_3 INT A N_5 VNW PCH W=0.66u L=0.06u
MNA2_2 INT B VSS VPW NCH W=0.26u L=0.06u
MPA2_3 VDD B N_5 VNW PCH W=0.66u L=0.06u
MNA2_3 INT B VSS VPW NCH W=0.26u L=0.06u
MPA2 VDD B N_7 VNW PCH W=0.66u L=0.06u
MNA1_3 INT A VSS VPW NCH W=0.26u L=0.06u
MPA1 INT A N_7 VNW PCH W=0.66u L=0.06u
MPA1_2 INT A N_9 VNW PCH W=0.66u L=0.06u
MNA1 INT A VSS VPW NCH W=0.26u L=0.06u
MNA2 INT B VSS VPW NCH W=0.26u L=0.06u
MPA2_2 N_9 B VDD VNW PCH W=0.66u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_4 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OR2X4MA10TR

****
.SUBCKT XOR2X4MA10TR VDD VSS VPW VNW Y A B
MNA108_3 NIN1 A VSS VPW NCH W=0.415u L=0.06u
MPA1010 NIN1 A VDD VNW PCH W=0.55u L=0.06u
MNA108_2 NIN1 A VSS VPW NCH W=0.415u L=0.06u
MPA1010_3 NIN1 A VDD VNW PCH W=0.55u L=0.06u
MNA108 NIN1 A VSS VPW NCH W=0.415u L=0.06u
MPA1010_2 NIN1 A VDD VNW PCH W=0.55u L=0.06u
MNA1_4 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_2 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_3 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_4 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1 NIN2 B VSS VPW NCH W=0.47u L=0.06u
MPA1_3 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNOE_4 Y A NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_3 Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MNOE_3 Y A NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_2 Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MNOE_2 Y A NIN2 VPW NCH W=0.47u L=0.06u
MPOEN Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MNOE Y A NIN2 VPW NCH W=0.47u L=0.06u
MPOEN_4 Y NIN1 NIN2 VNW PCH W=0.47u L=0.06u
MNOE02_4 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_4 Y A BIN2 VNW PCH W=0.47u L=0.06u
MNOE02_3 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_3 Y A BIN2 VNW PCH W=0.47u L=0.06u
MNOE02_2 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04_2 Y A BIN2 VNW PCH W=0.47u L=0.06u
MNOE02 Y NIN1 BIN2 VPW NCH W=0.47u L=0.06u
MPOEN04 Y A BIN2 VNW PCH W=0.47u L=0.06u
MNA1012 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_3 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012_3 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_2 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MPA1014 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012_2 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
MPA1014_4 BIN2 NIN2 VDD VNW PCH W=0.7u L=0.06u
MNA1012_4 BIN2 NIN2 VSS VPW NCH W=0.47u L=0.06u
.ENDS XOR2X4MA10TR

****
.SUBCKT OR2X6MA10TR VDD VSS VPW VNW Y A B
MPA1 INT A N_5 VNW PCH W=0.595u L=0.06u
MNA1_5 INT A VSS VPW NCH W=0.235u L=0.06u
MNA2_5 INT B VSS VPW NCH W=0.235u L=0.06u
MPA2 VDD B N_5 VNW PCH W=0.595u L=0.06u
MNA2_3 INT B VSS VPW NCH W=0.235u L=0.06u
MPA2_5 VDD B N_7 VNW PCH W=0.595u L=0.06u
MNA1_4 INT A VSS VPW NCH W=0.235u L=0.06u
MPA1_5 INT A N_7 VNW PCH W=0.595u L=0.06u
MPA1_3 INT A N_9 VNW PCH W=0.595u L=0.06u
MNA1_2 INT A VSS VPW NCH W=0.235u L=0.06u
MNA2_4 INT B VSS VPW NCH W=0.235u L=0.06u
MPA2_3 VDD B N_9 VNW PCH W=0.595u L=0.06u
MPA2_4 VDD B N_11 VNW PCH W=0.595u L=0.06u
MNA2_2 INT B VSS VPW NCH W=0.235u L=0.06u
MPA1_4 INT A N_11 VNW PCH W=0.595u L=0.06u
MNA1_3 INT A VSS VPW NCH W=0.235u L=0.06u
MPA1_2 INT A N_13 VNW PCH W=0.595u L=0.06u
MNA1 INT A VSS VPW NCH W=0.235u L=0.06u
MNA2 INT B VSS VPW NCH W=0.235u L=0.06u
MPA2_2 N_13 B VDD VNW PCH W=0.595u L=0.06u
MNA104_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_6 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_6 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_5 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_5 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OR2X6MA10TR

****
.SUBCKT OR2X8MA10TR VDD VSS VPW VNW Y A B
MNA2_4 INT B VSS VPW NCH W=0.26u L=0.06u
MPA2_6 VDD B N_96 VNW PCH W=0.66u L=0.06u
MNA1_6 INT A VSS VPW NCH W=0.26u L=0.06u
MPA1_6 INT A N_96 VNW PCH W=0.66u L=0.06u
MPA1_3 INT A N_98 VNW PCH W=0.66u L=0.06u
MNA1_5 INT A VSS VPW NCH W=0.26u L=0.06u
MNA2_3 INT B VSS VPW NCH W=0.26u L=0.06u
MPA2_3 VDD B N_98 VNW PCH W=0.66u L=0.06u
MNA2_2 INT B VSS VPW NCH W=0.26u L=0.06u
MPA2_2 VDD B N_100 VNW PCH W=0.66u L=0.06u
MNA1_4 INT A VSS VPW NCH W=0.26u L=0.06u
MPA1_2 INT A N_100 VNW PCH W=0.66u L=0.06u
MPA1_5 INT A N_102 VNW PCH W=0.66u L=0.06u
MNA1_3 INT A VSS VPW NCH W=0.26u L=0.06u
MNA2 INT B VSS VPW NCH W=0.26u L=0.06u
MPA2_5 VDD B N_102 VNW PCH W=0.66u L=0.06u
MPA2_4 VDD B N_104 VNW PCH W=0.66u L=0.06u
MNA2_6 INT B VSS VPW NCH W=0.26u L=0.06u
MPA1_4 INT A N_104 VNW PCH W=0.66u L=0.06u
MNA1_2 INT A VSS VPW NCH W=0.26u L=0.06u
MPA1 INT A N_106 VNW PCH W=0.66u L=0.06u
MNA1 INT A VSS VPW NCH W=0.26u L=0.06u
MNA2_5 INT B VSS VPW NCH W=0.26u L=0.06u
MPA2 N_106 B VDD VNW PCH W=0.66u L=0.06u
MNA104_3 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_3 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_7 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_7 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_6 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_6 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_5 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_5 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_4 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_4 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_2 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_2 Y INT VDD VNW PCH W=0.7u L=0.06u
MNA104_8 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA106_8 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OR2X8MA10TR

****
.SUBCKT NOR3X0P7MA10TR VDD VSS VPW VNW Y A B C
MPA3 VDD C N_5 VNW PCH W=0.49u L=0.06u
MNA3 Y C VSS VPW NCH W=0.15u L=0.06u
MPA2 N_5 B N_3 VNW PCH W=0.49u L=0.06u
MNA2 Y B VSS VPW NCH W=0.15u L=0.06u
MPA1 N_3 A Y VNW PCH W=0.49u L=0.06u
MNA1 Y A VSS VPW NCH W=0.15u L=0.06u
.ENDS NOR3X0P7MA10TR

****
.SUBCKT OR3X0P7MA10TR VDD VSS VPW VNW Y A B C
MPA3 VDD C N_5 VNW PCH W=0.395u L=0.06u
MPA2 N_5 B N_6 VNW PCH W=0.395u L=0.06u
MPA106 INT A N_6 VNW PCH W=0.395u L=0.06u
MNA102 INT A VSS VPW NCH W=0.26u L=0.06u
MPA106_2 INT A N_8 VNW PCH W=0.395u L=0.06u
MNA2 INT B VSS VPW NCH W=0.26u L=0.06u
MPA2_2 N_8 B N_9 VNW PCH W=0.395u L=0.06u
MNA3 INT C VSS VPW NCH W=0.26u L=0.06u
MPA3_2 N_9 C VDD VNW PCH W=0.395u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS OR3X0P7MA10TR

****
.SUBCKT XNOR3X0P7MA10TR VDD VSS VPW VNW Y A B C
MNA1020 NIN2 B VSS VPW NCH W=0.32u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.42u L=0.06u
MNA1 NIN3 C VSS VPW NCH W=0.37u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.37u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=0.555u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.455u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.37u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.455u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.37u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=0.555u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.24u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.32u L=0.06u
MNOE08 NOUT NIN1 XOR23 VPW NCH W=0.28u L=0.06u
MPOEN010 NOUT A XOR23 VNW PCH W=0.34u L=0.06u
MNOE012 NOUT A XNOR23 VPW NCH W=0.28u L=0.06u
MPOEN014 NOUT NIN1 XNOR23 VNW PCH W=0.34u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.28u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.42u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=0.37u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=0.49u L=0.06u
.ENDS XNOR3X0P7MA10TR

****
.SUBCKT XOR3X0P7MA10TR VDD VSS VPW VNW Y A B C
MNA1020 NIN2 B VSS VPW NCH W=0.32u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.42u L=0.06u
MNA1 NIN3 C VSS VPW NCH W=0.37u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=0.555u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.37u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.455u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.37u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.455u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.37u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=0.555u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.24u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.32u L=0.06u
MNOE08 NOUT A XOR23 VPW NCH W=0.28u L=0.06u
MPOEN010 NOUT NIN1 XOR23 VNW PCH W=0.34u L=0.06u
MNOE012 NOUT NIN1 XNOR23 VPW NCH W=0.28u L=0.06u
MPOEN014 NOUT A XNOR23 VNW PCH W=0.34u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.28u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.42u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=0.37u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=0.49u L=0.06u
.ENDS XOR3X0P7MA10TR

****
.SUBCKT NOR3X1MA10TR VDD VSS VPW VNW Y A B C
MPA3 VDD C N_5 VNW PCH W=0.7u L=0.06u
MNA3 Y C VSS VPW NCH W=0.205u L=0.06u
MPA2 N_5 B N_3 VNW PCH W=0.7u L=0.06u
MNA2 Y B VSS VPW NCH W=0.205u L=0.06u
MPA1 N_3 A Y VNW PCH W=0.7u L=0.06u
MNA1 Y A VSS VPW NCH W=0.205u L=0.06u
.ENDS NOR3X1MA10TR

****
.SUBCKT OR3X1MA10TR VDD VSS VPW VNW Y A B C
MPA3 VDD C N_5 VNW PCH W=0.5u L=0.06u
MPA2 N_5 B N_6 VNW PCH W=0.5u L=0.06u
MPA106 INT A N_6 VNW PCH W=0.5u L=0.06u
MNA102 INT A VSS VPW NCH W=0.33u L=0.06u
MPA106_2 INT A N_8 VNW PCH W=0.5u L=0.06u
MNA2 INT B VSS VPW NCH W=0.33u L=0.06u
MPA2_2 N_8 B N_9 VNW PCH W=0.5u L=0.06u
MNA3 INT C VSS VPW NCH W=0.33u L=0.06u
MPA3_2 N_9 C VDD VNW PCH W=0.5u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.53u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.7u L=0.06u
.ENDS OR3X1MA10TR

****
.SUBCKT XNOR3X1MA10TR VDD VSS VPW VNW Y A B C
MNA1020 NIN2 B VSS VPW NCH W=0.37u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.47u L=0.06u
MNA1 NIN3 C VSS VPW NCH W=0.47u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.47u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=0.7u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.47u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.47u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.47u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.47u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=0.7u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.28u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.36u L=0.06u
MNOE08 NOUT NIN1 XOR23 VPW NCH W=0.36u L=0.06u
MPOEN010 NOUT A XOR23 VNW PCH W=0.43u L=0.06u
MNOE012 NOUT A XNOR23 VPW NCH W=0.36u L=0.06u
MPOEN014 NOUT NIN1 XNOR23 VNW PCH W=0.43u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.36u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.54u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=0.53u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS XNOR3X1MA10TR

****
.SUBCKT XOR3X1MA10TR VDD VSS VPW VNW Y A B C
MNA1020 NIN2 B VSS VPW NCH W=0.37u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.47u L=0.06u
MNA1 NIN3 C VSS VPW NCH W=0.47u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.47u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=0.7u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.47u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.47u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.47u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.47u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=0.7u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.28u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.36u L=0.06u
MNOE08 NOUT A XOR23 VPW NCH W=0.36u L=0.06u
MPOEN010 NOUT NIN1 XOR23 VNW PCH W=0.43u L=0.06u
MNOE012 NOUT NIN1 XNOR23 VPW NCH W=0.36u L=0.06u
MPOEN014 NOUT A XNOR23 VNW PCH W=0.43u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.36u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.54u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=0.53u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS XOR3X1MA10TR

****
.SUBCKT NOR3X1P4MA10TR VDD VSS VPW VNW Y A B C
MPA3 VDD C N_18 VNW PCH W=0.49u L=0.06u
MPA2 N_18 B N_19 VNW PCH W=0.49u L=0.06u
MPA1 Y A N_19 VNW PCH W=0.49u L=0.06u
MPA1_2 Y A N_21 VNW PCH W=0.49u L=0.06u
MNA1 Y A VSS VPW NCH W=0.29u L=0.06u
MPA2_2 N_21 B N_16 VNW PCH W=0.49u L=0.06u
MNA2 Y B VSS VPW NCH W=0.29u L=0.06u
MPA3_2 N_16 C VDD VNW PCH W=0.49u L=0.06u
MNA3 Y C VSS VPW NCH W=0.29u L=0.06u
.ENDS NOR3X1P4MA10TR

****
.SUBCKT OR3X1P4MA10TR VDD VSS VPW VNW Y A B C
MNA3_2 INT C VSS VPW NCH W=0.23u L=0.06u
MPA3 VDD C N_5 VNW PCH W=0.7u L=0.06u
MNA2 INT B VSS VPW NCH W=0.23u L=0.06u
MPA2 N_5 B N_6 VNW PCH W=0.7u L=0.06u
MNA102 INT A VSS VPW NCH W=0.23u L=0.06u
MPA106 INT A N_6 VNW PCH W=0.7u L=0.06u
MPA106_2 INT A N_8 VNW PCH W=0.7u L=0.06u
MNA102_2 INT A VSS VPW NCH W=0.23u L=0.06u
MPA2_2 N_8 B N_10 VNW PCH W=0.7u L=0.06u
MNA2_2 INT B VSS VPW NCH W=0.23u L=0.06u
MNA3 INT C VSS VPW NCH W=0.23u L=0.06u
MPA3_2 N_10 C VDD VNW PCH W=0.7u L=0.06u
MNA1 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1 Y INT VDD VNW PCH W=0.49u L=0.06u
MNA1_2 Y INT VSS VPW NCH W=0.37u L=0.06u
MPA1_2 Y INT VDD VNW PCH W=0.49u L=0.06u
.ENDS OR3X1P4MA10TR

****
.SUBCKT XOR3X1P4MA10TR VDD VSS VPW VNW Y A B C
MNA1020 NIN2 B VSS VPW NCH W=0.53u L=0.06u
MPA1022 NIN2 B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 NIN3 C VSS VPW NCH W=0.33u L=0.06u
MPA1_2 NIN3 C VDD VNW PCH W=0.495u L=0.06u
MNA1 NIN3 C VSS VPW NCH W=0.33u L=0.06u
MPA1 NIN3 C VDD VNW PCH W=0.495u L=0.06u
MNOE_2 XOR23 B NIN3 VPW NCH W=0.33u L=0.06u
MPOEN_2 XOR23 NIN2 NIN3 VNW PCH W=0.33u L=0.06u
MNOE XOR23 B NIN3 VPW NCH W=0.33u L=0.06u
MPOEN XOR23 NIN2 NIN3 VNW PCH W=0.33u L=0.06u
MNOE02 XOR23 NIN2 BIN3 VPW NCH W=0.33u L=0.06u
MPOEN04_2 XOR23 B BIN3 VNW PCH W=0.33u L=0.06u
MNOE02_2 XOR23 NIN2 BIN3 VPW NCH W=0.33u L=0.06u
MPOEN04 XOR23 B BIN3 VNW PCH W=0.33u L=0.06u
MNA1028_2 BIN3 NIN3 VSS VPW NCH W=0.33u L=0.06u
MPA1030_2 BIN3 NIN3 VDD VNW PCH W=0.495u L=0.06u
MNA1028 BIN3 NIN3 VSS VPW NCH W=0.33u L=0.06u
MPA1030 BIN3 NIN3 VDD VNW PCH W=0.495u L=0.06u
MNA1024 NIN1 A VSS VPW NCH W=0.395u L=0.06u
MPA1026 NIN1 A VDD VNW PCH W=0.525u L=0.06u
MNOE08 NOUT A XOR23 VPW NCH W=0.47u L=0.06u
MPOEN010 NOUT NIN1 XOR23 VNW PCH W=0.57u L=0.06u
MNOE012 NOUT NIN1 XNOR23 VPW NCH W=0.47u L=0.06u
MPOEN014 NOUT A XNOR23 VNW PCH W=0.57u L=0.06u
MNA1016 XNOR23 XOR23 VSS VPW NCH W=0.47u L=0.06u
MPA1018 XNOR23 XOR23 VDD VNW PCH W=0.7u L=0.06u
MNA1032_2 Y NOUT VSS VPW NCH W=0.37u L=0.06u
MPA1034_2 Y NOUT VDD VNW PCH W=0.49u L=0.06u
MNA1032 Y NOUT VSS VPW NCH W=0.37u L=0.06u
MPA1034 Y NOUT VDD VNW PCH W=0.49u L=0.06u
.ENDS XOR3X1P4MA10TR

****
.SUBCKT OR4X2MA10TR VDD VSS VPW VNW Y A B C D
MPA2010_2 VDD D N_5 VNW PCH W=0.44u L=0.06u
MNA206 INT2 D VSS VPW NCH W=0.36u L=0.06u
MPA108_2 INT2 C N_5 VNW PCH W=0.44u L=0.06u
MNA104 INT2 C VSS VPW NCH W=0.36u L=0.06u
MPA108 INT2 C N_7 VNW PCH W=0.44u L=0.06u
MPA2010 N_7 D VDD VNW PCH W=0.44u L=0.06u
MNA2014 VSS INT2 N_34 VPW NCH W=0.58u L=0.06u
MPA2018_2 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_2 VSS INT2 N_34 VPW NCH W=0.58u L=0.06u
MPA2018 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA1012_2 N_34 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016_2 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012 N_34 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MPA2_2 VDD B N_13 VNW PCH W=0.44u L=0.06u
MPA1_2 INT1 A N_13 VNW PCH W=0.44u L=0.06u
MNA1 INT1 A VSS VPW NCH W=0.36u L=0.06u
MPA1 INT1 A N_3 VNW PCH W=0.44u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.36u L=0.06u
MPA2 N_3 B VDD VNW PCH W=0.44u L=0.06u
.ENDS OR4X2MA10TR

****
.SUBCKT OR4X3MA10TR VDD VSS VPW VNW Y A B C D
MPA2010 VDD D N_5 VNW PCH W=0.66u L=0.06u
MNA206 INT2 D VSS VPW NCH W=0.54u L=0.06u
MPA108 INT2 C N_5 VNW PCH W=0.66u L=0.06u
MNA104 INT2 C VSS VPW NCH W=0.54u L=0.06u
MPA108_2 INT2 C N_7 VNW PCH W=0.66u L=0.06u
MPA2010_2 N_7 D VDD VNW PCH W=0.66u L=0.06u
MNA2014 N_39 INT2 VSS VPW NCH W=0.58u L=0.06u
MPA2018_2 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_3 VSS INT2 N_39 VPW NCH W=0.58u L=0.06u
MPA2018 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_2 VSS INT2 N_39 VPW NCH W=0.58u L=0.06u
MPA2018_3 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA1012 Y INT1 N_39 VPW NCH W=0.58u L=0.06u
MPA1016_2 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_3 N_39 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_2 Y INT1 N_39 VPW NCH W=0.58u L=0.06u
MPA1016_3 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MPA2_2 VDD B N_15 VNW PCH W=0.66u L=0.06u
MPA1_2 INT1 A N_15 VNW PCH W=0.66u L=0.06u
MNA1 INT1 A VSS VPW NCH W=0.54u L=0.06u
MPA1 INT1 A N_3 VNW PCH W=0.66u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.54u L=0.06u
MPA2 N_3 B VDD VNW PCH W=0.66u L=0.06u
.ENDS OR4X3MA10TR

****
.SUBCKT OR4X4MA10TR VDD VSS VPW VNW Y A B C D
MPA108_2 INT2 C N_5 VNW PCH W=0.59u L=0.06u
MNA206 INT2 D VSS VPW NCH W=0.36u L=0.06u
MPA2010_2 VDD D N_5 VNW PCH W=0.59u L=0.06u
MPA2010 VDD D N_7 VNW PCH W=0.59u L=0.06u
MNA206_2 INT2 D VSS VPW NCH W=0.36u L=0.06u
MPA108 INT2 C N_7 VNW PCH W=0.59u L=0.06u
MNA104_2 INT2 C VSS VPW NCH W=0.36u L=0.06u
MPA108_3 INT2 C N_10 VNW PCH W=0.59u L=0.06u
MNA104 INT2 C VSS VPW NCH W=0.36u L=0.06u
MPA2010_3 N_10 D VDD VNW PCH W=0.59u L=0.06u
MNA2014_3 VSS INT2 N_54 VPW NCH W=0.58u L=0.06u
MPA2018 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_2 N_54 INT2 VSS VPW NCH W=0.58u L=0.06u
MPA2018_4 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014 VSS INT2 N_54 VPW NCH W=0.58u L=0.06u
MPA2018_3 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_4 VSS INT2 N_54 VPW NCH W=0.58u L=0.06u
MPA2018_2 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA1012_3 Y INT1 N_54 VPW NCH W=0.58u L=0.06u
MPA1016 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_2 N_54 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016_4 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012 Y INT1 N_54 VPW NCH W=0.58u L=0.06u
MPA1016_3 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_4 N_54 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016_2 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MPA2 VDD B N_19 VNW PCH W=0.59u L=0.06u
MNA1 INT1 A VSS VPW NCH W=0.36u L=0.06u
MPA1 INT1 A N_19 VNW PCH W=0.59u L=0.06u
MPA1_3 INT1 A N_21 VNW PCH W=0.59u L=0.06u
MNA1_2 INT1 A VSS VPW NCH W=0.36u L=0.06u
MPA2_3 VDD B N_21 VNW PCH W=0.59u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.36u L=0.06u
MPA2_2 VDD B N_3 VNW PCH W=0.59u L=0.06u
MNA2_2 INT1 B VSS VPW NCH W=0.36u L=0.06u
MPA1_2 N_3 A INT1 VNW PCH W=0.59u L=0.06u
.ENDS OR4X4MA10TR

****
.SUBCKT OR4X6MA10TR VDD VSS VPW VNW Y A B C D
MPA2010_2 VDD D N_5 VNW PCH W=0.66u L=0.06u
MNA206_3 INT2 D VSS VPW NCH W=0.36u L=0.06u
MPA108_2 INT2 C N_5 VNW PCH W=0.66u L=0.06u
MNA104_2 INT2 C VSS VPW NCH W=0.36u L=0.06u
MPA108 INT2 C N_7 VNW PCH W=0.66u L=0.06u
MNA104 INT2 C VSS VPW NCH W=0.36u L=0.06u
MPA2010 VDD D N_7 VNW PCH W=0.66u L=0.06u
MNA206_2 INT2 D VSS VPW NCH W=0.36u L=0.06u
MPA2010_4 VDD D N_9 VNW PCH W=0.66u L=0.06u
MNA206 INT2 D VSS VPW NCH W=0.36u L=0.06u
MPA108_4 INT2 C N_9 VNW PCH W=0.66u L=0.06u
MNA104_3 INT2 C VSS VPW NCH W=0.36u L=0.06u
MPA108_3 INT2 C N_11 VNW PCH W=0.66u L=0.06u
MPA2010_3 N_11 D VDD VNW PCH W=0.66u L=0.06u
MNA2014_5 VSS INT2 N_74 VPW NCH W=0.58u L=0.06u
MPA2018 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_4 N_74 INT2 VSS VPW NCH W=0.58u L=0.06u
MPA2018_6 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_3 VSS INT2 N_74 VPW NCH W=0.58u L=0.06u
MPA2018_5 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_2 N_74 INT2 VSS VPW NCH W=0.58u L=0.06u
MPA2018_4 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014 VSS INT2 N_74 VPW NCH W=0.58u L=0.06u
MPA2018_3 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_6 VSS INT2 N_74 VPW NCH W=0.58u L=0.06u
MPA2018_2 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA1012_5 Y INT1 N_74 VPW NCH W=0.58u L=0.06u
MPA1016 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_4 N_74 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016_6 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_3 Y INT1 N_74 VPW NCH W=0.58u L=0.06u
MPA1016_5 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_2 N_74 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016_4 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012 Y INT1 N_74 VPW NCH W=0.58u L=0.06u
MPA1016_3 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_6 N_74 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016_2 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MPA2 VDD B N_25 VNW PCH W=0.66u L=0.06u
MPA1 INT1 A N_25 VNW PCH W=0.66u L=0.06u
MNA1_3 INT1 A VSS VPW NCH W=0.36u L=0.06u
MPA1_3 INT1 A N_27 VNW PCH W=0.66u L=0.06u
MNA2_2 INT1 B VSS VPW NCH W=0.36u L=0.06u
MPA2_3 VDD B N_27 VNW PCH W=0.66u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.36u L=0.06u
MPA2_2 VDD B N_29 VNW PCH W=0.66u L=0.06u
MNA1_2 INT1 A VSS VPW NCH W=0.36u L=0.06u
MPA1_2 INT1 A N_29 VNW PCH W=0.66u L=0.06u
MNA1 INT1 A VSS VPW NCH W=0.36u L=0.06u
MPA1_4 INT1 A N_3 VNW PCH W=0.66u L=0.06u
MNA2_3 INT1 B VSS VPW NCH W=0.36u L=0.06u
MPA2_4 N_3 B VDD VNW PCH W=0.66u L=0.06u
.ENDS OR4X6MA10TR

****
.SUBCKT OR4X8MA10TR VDD VSS VPW VNW Y A B C D
MPA108_4 INT2 C N_5 VNW PCH W=0.7u L=0.06u
MNA104_3 INT2 C VSS VPW NCH W=0.355u L=0.06u
MPA2010_4 VDD D N_5 VNW PCH W=0.7u L=0.06u
MNA206_3 INT2 D VSS VPW NCH W=0.355u L=0.06u
MPA2010 VDD D N_7 VNW PCH W=0.7u L=0.06u
MNA206 INT2 D VSS VPW NCH W=0.355u L=0.06u
MPA108 INT2 C N_7 VNW PCH W=0.7u L=0.06u
MNA104 INT2 C VSS VPW NCH W=0.355u L=0.06u
MPA108_5 INT2 C N_9 VNW PCH W=0.7u L=0.06u
MNA104_4 INT2 C VSS VPW NCH W=0.355u L=0.06u
MPA2010_5 VDD D N_9 VNW PCH W=0.7u L=0.06u
MNA206_2 INT2 D VSS VPW NCH W=0.355u L=0.06u
MPA2010_3 VDD D N_11 VNW PCH W=0.7u L=0.06u
MNA206_4 INT2 D VSS VPW NCH W=0.36u L=0.06u
MPA108_3 INT2 C N_11 VNW PCH W=0.7u L=0.06u
MPA108_2 INT2 C N_14 VNW PCH W=0.7u L=0.06u
MNA104_2 INT2 C VSS VPW NCH W=0.36u L=0.06u
MPA2010_2 N_14 D VDD VNW PCH W=0.7u L=0.06u
MNA2014_5 VSS INT2 N_85 VPW NCH W=0.58u L=0.06u
MPA2018_7 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_4 N_85 INT2 VSS VPW NCH W=0.58u L=0.06u
MPA2018_6 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_2 VSS INT2 N_85 VPW NCH W=0.58u L=0.06u
MPA2018_5 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_6 N_85 INT2 VSS VPW NCH W=0.58u L=0.06u
MPA2018_4 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_3 VSS INT2 N_85 VPW NCH W=0.58u L=0.06u
MPA2018_3 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014 N_85 INT2 VSS VPW NCH W=0.58u L=0.06u
MPA2018_2 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_8 VSS INT2 N_85 VPW NCH W=0.58u L=0.06u
MPA2018 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2014_7 N_85 INT2 VSS VPW NCH W=0.58u L=0.06u
MPA2018_8 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA1012_5 Y INT1 N_85 VPW NCH W=0.58u L=0.06u
MPA1016_5 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_3 N_85 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016_3 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_8 Y INT1 N_85 VPW NCH W=0.58u L=0.06u
MPA1016_2 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_7 Y INT1 N_85 VPW NCH W=0.58u L=0.06u
MPA1016 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_6 Y INT1 N_85 VPW NCH W=0.58u L=0.06u
MPA1016_8 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_4 N_85 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016_7 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012_2 Y INT1 N_85 VPW NCH W=0.58u L=0.06u
MPA1016_6 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1012 N_85 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1016_4 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MPA2 VDD B N_31 VNW PCH W=0.7u L=0.06u
MPA1 INT1 A N_31 VNW PCH W=0.7u L=0.06u
MNA1_4 INT1 A VSS VPW NCH W=0.36u L=0.06u
MPA1_3 INT1 A N_33 VNW PCH W=0.7u L=0.06u
MNA2_4 INT1 B VSS VPW NCH W=0.36u L=0.06u
MPA2_3 VDD B N_33 VNW PCH W=0.7u L=0.06u
MNA2_3 INT1 B VSS VPW NCH W=0.355u L=0.06u
MPA2_2 N_35 B VDD VNW PCH W=0.7u L=0.06u
MNA1_2 INT1 A VSS VPW NCH W=0.355u L=0.06u
MPA1_2 INT1 A N_35 VNW PCH W=0.7u L=0.06u
MNA1 INT1 A VSS VPW NCH W=0.355u L=0.06u
MPA1_4 INT1 A N_37 VNW PCH W=0.7u L=0.06u
MNA2_2 INT1 B VSS VPW NCH W=0.355u L=0.06u
MPA2_4 VDD B N_37 VNW PCH W=0.7u L=0.06u
MPA2_5 VDD B N_3 VNW PCH W=0.7u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.355u L=0.06u
MPA1_5 N_3 A INT1 VNW PCH W=0.7u L=0.06u
MNA1_3 INT1 A VSS VPW NCH W=0.355u L=0.06u
.ENDS OR4X8MA10TR

****
.SUBCKT OR6X1P4MA10TR VDD VSS VPW VNW Y A B C D E F
MPA3016_2 VDD F N_5 VNW PCH W=0.51u L=0.06u
MNA3010 INT2 F VSS VPW NCH W=0.3u L=0.06u
MPA2014_2 N_5 E N_6 VNW PCH W=0.51u L=0.06u
MNA208 INT2 E VSS VPW NCH W=0.3u L=0.06u
MPA1012_2 INT2 D N_6 VNW PCH W=0.51u L=0.06u
MNA106 INT2 D VSS VPW NCH W=0.3u L=0.06u
MPA1012 INT2 D N_8 VNW PCH W=0.51u L=0.06u
MPA2014 N_8 E N_10 VNW PCH W=0.51u L=0.06u
MPA3016 N_10 F VDD VNW PCH W=0.51u L=0.06u
MNA2020_2 VSS INT2 N_44 VPW NCH W=0.41u L=0.06u
MPA2024 Y INT2 VDD VNW PCH W=0.34u L=0.06u
MNA2020 VSS INT2 N_44 VPW NCH W=0.41u L=0.06u
MPA2024_2 Y INT2 VDD VNW PCH W=0.34u L=0.06u
MNA1018_2 N_44 INT1 Y VPW NCH W=0.41u L=0.06u
MPA1022_2 Y INT1 VDD VNW PCH W=0.34u L=0.06u
MNA1018 N_44 INT1 Y VPW NCH W=0.41u L=0.06u
MPA1022 Y INT1 VDD VNW PCH W=0.34u L=0.06u
MPA3_2 VDD C N_15 VNW PCH W=0.51u L=0.06u
MPA2_2 N_15 B N_16 VNW PCH W=0.51u L=0.06u
MPA1_2 INT1 A N_16 VNW PCH W=0.51u L=0.06u
MNA1 INT1 A VSS VPW NCH W=0.3u L=0.06u
MPA1 INT1 A N_18 VNW PCH W=0.51u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.3u L=0.06u
MPA2 N_18 B N_3 VNW PCH W=0.51u L=0.06u
MNA3 INT1 C VSS VPW NCH W=0.3u L=0.06u
MPA3 N_3 C VDD VNW PCH W=0.51u L=0.06u
.ENDS OR6X1P4MA10TR

****
.SUBCKT OR6X2MA10TR VDD VSS VPW VNW Y A B C D E F
MPA3016_2 VDD F N_5 VNW PCH W=0.665u L=0.06u
MNA3010 INT2 F VSS VPW NCH W=0.39u L=0.06u
MPA2014_2 N_5 E N_6 VNW PCH W=0.665u L=0.06u
MNA208 INT2 E VSS VPW NCH W=0.39u L=0.06u
MPA1012_2 INT2 D N_6 VNW PCH W=0.665u L=0.06u
MNA106 INT2 D VSS VPW NCH W=0.39u L=0.06u
MPA1012 INT2 D N_8 VNW PCH W=0.665u L=0.06u
MPA2014 N_8 E N_9 VNW PCH W=0.665u L=0.06u
MPA3016 N_9 F VDD VNW PCH W=0.665u L=0.06u
MNA2020_2 VSS INT2 N_44 VPW NCH W=0.58u L=0.06u
MPA2024 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA2020 VSS INT2 N_44 VPW NCH W=0.58u L=0.06u
MPA2024_2 Y INT2 VDD VNW PCH W=0.48u L=0.06u
MNA1018_2 N_44 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1022_2 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MNA1018 N_44 INT1 Y VPW NCH W=0.58u L=0.06u
MPA1022 Y INT1 VDD VNW PCH W=0.48u L=0.06u
MPA3_2 VDD C N_15 VNW PCH W=0.665u L=0.06u
MPA2_2 N_15 B N_16 VNW PCH W=0.665u L=0.06u
MPA1_2 INT1 A N_16 VNW PCH W=0.665u L=0.06u
MNA1 INT1 A VSS VPW NCH W=0.39u L=0.06u
MPA1 INT1 A N_18 VNW PCH W=0.665u L=0.06u
MNA2 INT1 B VSS VPW NCH W=0.39u L=0.06u
MPA2 N_18 B N_3 VNW PCH W=0.665u L=0.06u
MNA3 INT1 C VSS VPW NCH W=0.39u L=0.06u
MPA3 N_3 C VDD VNW PCH W=0.665u L=0.06u
.ENDS OR6X2MA10TR

****
.SUBCKT POSTICGX11BA10TR VDD VSS VPW VNW ECK CK E SEN
MNA1012 NCLK_ CK VSS VPW NCH W=0.2u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.26u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.51u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.38u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.38u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.38u L=0.06u
MPOEN07 N_177 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_197 CK NM VPW NCH W=0.15u L=0.06u
MPA1 N_177 M VDD VNW PCH W=0.15u L=0.06u
MNA1 N_197 M VSS VPW NCH W=0.15u L=0.06u
MNA2 VSS SEN N_199 VPW NCH W=0.435u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.32u L=0.06u
MNA1020 M NM N_199 VPW NCH W=0.435u L=0.06u
MPA1023_2 M NM VDD VNW PCH W=0.32u L=0.06u
MNA1020_2 M NM N_202 VPW NCH W=0.435u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.32u L=0.06u
MNA2_2 N_202 SEN VSS VPW NCH W=0.435u L=0.06u
MN1_4 VSS M N_203 VPW NCH W=0.465u L=0.06u
MPA2_2 M SEN VDD VNW PCH W=0.32u L=0.06u
MN0_4 NOUT CK N_203 VPW NCH W=0.465u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN0_2 N_205 CK NOUT VPW NCH W=0.465u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN1_2 VSS M N_205 VPW NCH W=0.465u L=0.06u
MN1 VSS M N_207 VPW NCH W=0.465u L=0.06u
MN0 NOUT CK N_207 VPW NCH W=0.465u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN0_3 N_210 CK NOUT VPW NCH W=0.465u L=0.06u
MP1_4 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN1_3 N_210 M VSS VPW NCH W=0.465u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.23u L=0.06u
MNA1026_10 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_8 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_10 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_9 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_9 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_7 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_8 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.36u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS POSTICGX11BA10TR

****
.SUBCKT POSTICGX13BA10TR VDD VSS VPW VNW ECK CK E SEN
MNA1012 NCLK_ CK VSS VPW NCH W=0.21u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.28u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.555u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.42u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.42u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.42u L=0.06u
MPOEN07 N_187 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_209 CK NM VPW NCH W=0.15u L=0.06u
MPA1 N_187 M VDD VNW PCH W=0.15u L=0.06u
MNA1 N_209 M VSS VPW NCH W=0.15u L=0.06u
MNA2_2 VSS SEN N_211 VPW NCH W=0.48u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.35u L=0.06u
MNA1020_2 M NM N_211 VPW NCH W=0.48u L=0.06u
MPA1023_2 M NM VDD VNW PCH W=0.35u L=0.06u
MNA1020 M NM N_213 VPW NCH W=0.48u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.35u L=0.06u
MNA2 VSS SEN N_213 VPW NCH W=0.48u L=0.06u
MN1_4 VSS M N_215 VPW NCH W=0.555u L=0.06u
MPA2_2 M SEN VDD VNW PCH W=0.35u L=0.06u
MN0_4 NOUT CK N_215 VPW NCH W=0.555u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN0_2 N_217 CK NOUT VPW NCH W=0.555u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN1_2 VSS M N_217 VPW NCH W=0.555u L=0.06u
MN1_3 VSS M N_219 VPW NCH W=0.555u L=0.06u
MN0_3 NOUT CK N_219 VPW NCH W=0.555u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN0 N_222 CK NOUT VPW NCH W=0.555u L=0.06u
MP1_4 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN1 N_222 M VSS VPW NCH W=0.555u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.27u L=0.06u
MNA1026_7 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_10 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_11 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_8 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_9 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_11 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_9 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_10 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_8 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS POSTICGX13BA10TR

****
.SUBCKT POSTICGX16BA10TR VDD VSS VPW VNW ECK CK E SEN
MNA1012 NCLK_ CK VSS VPW NCH W=0.24u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.32u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.66u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.5u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.5u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.5u L=0.06u
MPOEN07 N_218 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_225 CK NM VPW NCH W=0.15u L=0.06u
MPA1 N_218 M VDD VNW PCH W=0.15u L=0.06u
MNA1 N_225 M VSS VPW NCH W=0.15u L=0.06u
MNA2_2 VSS SEN N_227 VPW NCH W=0.58u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.425u L=0.06u
MNA1020_2 M NM N_227 VPW NCH W=0.58u L=0.06u
MPA1023_2 M NM VDD VNW PCH W=0.425u L=0.06u
MNA1020 N_229 NM M VPW NCH W=0.58u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.425u L=0.06u
MPA2_2 M SEN VDD VNW PCH W=0.425u L=0.06u
MNA2 VSS SEN N_229 VPW NCH W=0.58u L=0.06u
MN1_5 VSS M N_231 VPW NCH W=0.54u L=0.06u
MN0_5 NOUT CK N_231 VPW NCH W=0.54u L=0.06u
MP1_5 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN0 N_233 CK NOUT VPW NCH W=0.54u L=0.06u
MP1_4 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN1 VSS M N_233 VPW NCH W=0.54u L=0.06u
MN1_3 VSS M N_235 VPW NCH W=0.54u L=0.06u
MN0_3 NOUT CK N_235 VPW NCH W=0.54u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN0_4 N_241 CK NOUT VPW NCH W=0.54u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN1_4 VSS M N_241 VPW NCH W=0.54u L=0.06u
MN1_2 N_239 M VSS VPW NCH W=0.54u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.33u L=0.06u
MN0_2 NOUT CK N_239 VPW NCH W=0.54u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MPA1028_10 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_11 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_8 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_9 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_14 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_13 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_12 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_8 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_7 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_13 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_12 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_11 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_10 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_9 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.75u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS POSTICGX16BA10TR

****
.SUBCKT POSTICGX3P5BA10TR VDD VSS VPW VNW ECK CK E SEN
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.32u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.18u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.18u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.18u L=0.06u
MPOEN07 N_16 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_30 CK NM VPW NCH W=0.15u L=0.06u
MPA1 N_16 M VDD VNW PCH W=0.15u L=0.06u
MNA1 VSS M N_30 VPW NCH W=0.15u L=0.06u
MNA2 N_41 SEN VSS VPW NCH W=0.415u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.305u L=0.06u
MNA1020 N_41 NM M VPW NCH W=0.415u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.305u L=0.06u
MN1_2 VSS M N_38 VPW NCH W=0.305u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.375u L=0.06u
MN0_2 NOUT CK N_38 VPW NCH W=0.305u L=0.06u
MN0 N_36 CK NOUT VPW NCH W=0.305u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.375u L=0.06u
MN1 VSS M N_36 VPW NCH W=0.305u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.42u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.42u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.42u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
.ENDS POSTICGX3P5BA10TR

****
.SUBCKT POSTICGX4BA10TR VDD VSS VPW VNW ECK CK E SEN
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.325u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.185u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.185u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.185u L=0.06u
MPOEN07 N_25 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_30 CK NM VPW NCH W=0.15u L=0.06u
MPA1 N_25 M VDD VNW PCH W=0.15u L=0.06u
MNA1 VSS M N_30 VPW NCH W=0.15u L=0.06u
MNA2 N_41 SEN VSS VPW NCH W=0.425u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.31u L=0.06u
MNA1020 N_41 NM M VPW NCH W=0.425u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.31u L=0.06u
MN1_2 VSS M N_34 VPW NCH W=0.34u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.41u L=0.06u
MN0_2 NOUT CK N_34 VPW NCH W=0.34u L=0.06u
MN0 N_32 CK NOUT VPW NCH W=0.34u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.41u L=0.06u
MN1 VSS M N_32 VPW NCH W=0.34u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.48u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.48u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.48u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS POSTICGX4BA10TR

****
.SUBCKT POSTICGX5BA10TR VDD VSS VPW VNW ECK CK E SEN
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.36u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.22u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.22u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.22u L=0.06u
MPOEN07 N_30 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_48 CK NM VPW NCH W=0.15u L=0.06u
MPA1 N_30 M VDD VNW PCH W=0.15u L=0.06u
MNA1 N_48 M VSS VPW NCH W=0.15u L=0.06u
MNA2 VSS SEN N_44 VPW NCH W=0.505u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.37u L=0.06u
MNA1020 N_44 NM M VPW NCH W=0.505u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.37u L=0.06u
MN1 VSS M N_36 VPW NCH W=0.43u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN0 NOUT CK N_36 VPW NCH W=0.43u L=0.06u
MN0_2 N_34 CK NOUT VPW NCH W=0.43u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN1_2 VSS M N_34 VPW NCH W=0.43u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS POSTICGX5BA10TR

****
.SUBCKT POSTICGX6BA10TR VDD VSS VPW VNW ECK CK E SEN
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.385u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.24u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.24u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.24u L=0.06u
MPOEN07 N_32 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_51 CK NM VPW NCH W=0.15u L=0.06u
MPA1 N_32 M VDD VNW PCH W=0.15u L=0.06u
MNA1 N_51 M VSS VPW NCH W=0.15u L=0.06u
MNA2 VSS SEN N_47 VPW NCH W=0.56u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.41u L=0.06u
MNA1020 N_47 NM M VPW NCH W=0.56u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.41u L=0.06u
MN1_2 VSS M N_44 VPW NCH W=0.51u L=0.06u
MN0_2 NOUT CK N_44 VPW NCH W=0.51u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.615u L=0.06u
MN0 N_42 CK NOUT VPW NCH W=0.51u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.615u L=0.06u
MN1 VSS M N_42 VPW NCH W=0.51u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.435u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.435u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS POSTICGX6BA10TR

****
.SUBCKT POSTICGX7P5BA10TR VDD VSS VPW VNW ECK CK E SEN
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.4u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.285u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.285u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.285u L=0.06u
MPOEN07 N_139 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_174 CK NM VPW NCH W=0.15u L=0.06u
MPA1 N_139 M VDD VNW PCH W=0.15u L=0.06u
MNA1 N_174 M VSS VPW NCH W=0.15u L=0.06u
MNA2 VSS SEN N_176 VPW NCH W=0.33u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.24u L=0.06u
MNA1020 M NM N_176 VPW NCH W=0.33u L=0.06u
MPA1023_2 M NM VDD VNW PCH W=0.24u L=0.06u
MNA1020_2 M NM N_179 VPW NCH W=0.33u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.24u L=0.06u
MNA2_2 N_179 SEN VSS VPW NCH W=0.33u L=0.06u
MN1_3 VSS M N_180 VPW NCH W=0.43u L=0.06u
MPA2_2 M SEN VDD VNW PCH W=0.24u L=0.06u
MN0_3 NOUT CK N_180 VPW NCH W=0.43u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN0_2 N_182 CK NOUT VPW NCH W=0.43u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN1_2 VSS M N_182 VPW NCH W=0.43u L=0.06u
MN1 VSS M N_170 VPW NCH W=0.43u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.16u L=0.06u
MN0 N_170 CK NOUT VPW NCH W=0.43u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.69u L=0.06u
.ENDS POSTICGX7P5BA10TR

****
.SUBCKT POSTICGX9BA10TR VDD VSS VPW VNW ECK CK E SEN
MNA1012 NCLK_ CK VSS VPW NCH W=0.17u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.225u L=0.06u
MPA1018 NEN E VDD VNW PCH W=0.45u L=0.06u
MNA1016 NEN E VSS VPW NCH W=0.33u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.33u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.33u L=0.06u
MPOEN07 N_135 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_183 CK NM VPW NCH W=0.15u L=0.06u
MPA1 N_135 M VDD VNW PCH W=0.15u L=0.06u
MNA1 N_183 M VSS VPW NCH W=0.15u L=0.06u
MNA2 VSS SEN N_185 VPW NCH W=0.38u L=0.06u
MPA2 M SEN VDD VNW PCH W=0.28u L=0.06u
MNA1020 M NM N_185 VPW NCH W=0.38u L=0.06u
MPA1023_2 M NM VDD VNW PCH W=0.28u L=0.06u
MNA1020_2 M NM N_188 VPW NCH W=0.38u L=0.06u
MPA1023 M NM VDD VNW PCH W=0.28u L=0.06u
MNA2_2 N_188 SEN VSS VPW NCH W=0.38u L=0.06u
MN1_2 VSS M N_189 VPW NCH W=0.515u L=0.06u
MPA2_2 M SEN VDD VNW PCH W=0.28u L=0.06u
MN0_2 NOUT CK N_189 VPW NCH W=0.515u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.62u L=0.06u
MN0 N_191 CK NOUT VPW NCH W=0.515u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.62u L=0.06u
MN1 VSS M N_191 VPW NCH W=0.515u L=0.06u
MN1_3 VSS M N_179 VPW NCH W=0.515u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.19u L=0.06u
MN0_3 N_179 CK NOUT VPW NCH W=0.515u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.62u L=0.06u
MNA1026_8 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_8 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026_7 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS POSTICGX9BA10TR

****
.SUBCKT PREICGX11BA10TR VDD VSS VPW VNW ECK CK E SE
MPA2_2 VDD SE N_18 VNW PCH W=0.54u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.38u L=0.06u
MPA2 VDD SE N_18 VNW PCH W=0.54u L=0.06u
MPA1023 N_18 E NEN VNW PCH W=0.48u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.38u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.38u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.38u L=0.06u
MPOEN07 N_171 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 NM CK N_220 VPW NCH W=0.15u L=0.06u
MNA1 VSS M N_220 VPW NCH W=0.15u L=0.06u
MPA1 N_171 M VDD VNW PCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.515u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.645u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.2u L=0.06u
MN1 N_189 M VSS VPW NCH W=0.465u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.26u L=0.06u
MN0 NOUT CK N_189 VPW NCH W=0.465u L=0.06u
MP1_4 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN0_4 N_191 CK NOUT VPW NCH W=0.465u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN1_4 VSS M N_191 VPW NCH W=0.465u L=0.06u
MN1_2 VSS M N_193 VPW NCH W=0.465u L=0.06u
MN0_2 NOUT CK N_193 VPW NCH W=0.465u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN0_3 N_196 CK NOUT VPW NCH W=0.465u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.57u L=0.06u
MN1_3 N_196 M VSS VPW NCH W=0.465u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.23u L=0.06u
MNA1026_8 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_10 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_8 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_10 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_9 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_7 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.8u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.4u L=0.06u
MPA1028_9 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.36u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS PREICGX11BA10TR

****
.SUBCKT PREICGX13BA10TR VDD VSS VPW VNW ECK CK E SE
MPA2_2 VDD SE N_5 VNW PCH W=0.6u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.42u L=0.06u
MPA2 VDD SE N_5 VNW PCH W=0.6u L=0.06u
MPA1023 N_5 E NEN VNW PCH W=0.52u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.42u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.42u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.42u L=0.06u
MPOEN07 N_176 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 NM CK N_207 VPW NCH W=0.15u L=0.06u
MNA1 VSS M N_207 VPW NCH W=0.15u L=0.06u
MPA1 N_176 M VDD VNW PCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.58u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.7u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.21u L=0.06u
MN1 N_211 M VSS VPW NCH W=0.555u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.28u L=0.06u
MN0 NOUT CK N_211 VPW NCH W=0.555u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN0_4 N_213 CK NOUT VPW NCH W=0.555u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN1_4 VSS M N_213 VPW NCH W=0.555u L=0.06u
MN1_2 VSS M N_215 VPW NCH W=0.555u L=0.06u
MN0_2 NOUT CK N_215 VPW NCH W=0.555u L=0.06u
MP1_4 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN0_3 N_218 CK NOUT VPW NCH W=0.555u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.67u L=0.06u
MN1_3 N_218 M VSS VPW NCH W=0.555u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.27u L=0.06u
MNA1026_9 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_7 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_11 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_11 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_9 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_8 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_10 ECK NOUT VDD VNW PCH W=0.855u L=0.06u
MNA1026_10 ECK NOUT VSS VPW NCH W=0.425u L=0.06u
MPA1028_8 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS PREICGX13BA10TR

****
.SUBCKT PREICGX16BA10TR VDD VSS VPW VNW ECK CK E SE
MPA2_2 VDD SE N_5 VNW PCH W=0.7u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.5u L=0.06u
MPA2 VDD SE N_5 VNW PCH W=0.7u L=0.06u
MPA1023 N_5 E NEN VNW PCH W=0.62u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.5u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.5u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.5u L=0.06u
MPOEN07 N_206 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 NM CK N_242 VPW NCH W=0.15u L=0.06u
MNA1 VSS M N_242 VPW NCH W=0.15u L=0.06u
MPA1 N_206 M VDD VNW PCH W=0.15u L=0.06u
MNA1016_2 M NM VSS VPW NCH W=0.34u L=0.06u
MPA1018_2 M NM VDD VNW PCH W=0.425u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.34u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.425u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.24u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.32u L=0.06u
MN1_3 VSS M N_251 VPW NCH W=0.54u L=0.06u
MN0_3 NOUT CK N_251 VPW NCH W=0.54u L=0.06u
MP1_4 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN0 N_253 CK NOUT VPW NCH W=0.54u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN1 VSS M N_253 VPW NCH W=0.54u L=0.06u
MN1_4 VSS M N_255 VPW NCH W=0.54u L=0.06u
MN0_4 NOUT CK N_255 VPW NCH W=0.54u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN0_2 N_261 CK NOUT VPW NCH W=0.54u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MN1_2 VSS M N_261 VPW NCH W=0.54u L=0.06u
MN1_5 VSS M N_259 VPW NCH W=0.54u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.33u L=0.06u
MN0_5 N_259 CK NOUT VPW NCH W=0.54u L=0.06u
MP1_5 NOUT CK VDD VNW PCH W=0.66u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_13 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_11 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_12 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_10 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.44u L=0.06u
MPA1028_8 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_10 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_9 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_8 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_14 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_9 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_12 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.835u L=0.06u
MNA1026_7 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_13 ECK NOUT VDD VNW PCH W=0.75u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.445u L=0.06u
MPA1028_11 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS PREICGX16BA10TR

****
.SUBCKT PREICGX3P5BA10TR VDD VSS VPW VNW ECK CK E SE
MNA2 NEN SE VSS VPW NCH W=0.18u L=0.06u
MPA2 VDD SE N_7 VNW PCH W=0.63u L=0.06u
MPA1023 NEN E N_7 VNW PCH W=0.225u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.18u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.18u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.18u L=0.06u
MPOEN07 N_26 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_32 CK NM VPW NCH W=0.15u L=0.06u
MNA1 VSS M N_32 VPW NCH W=0.15u L=0.06u
MPA1 N_26 M VDD VNW PCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.24u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.305u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MN1_2 N_42 M VSS VPW NCH W=0.305u L=0.06u
MN0_2 NOUT CK N_42 VPW NCH W=0.305u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.375u L=0.06u
MN0 N_40 CK NOUT VPW NCH W=0.305u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.375u L=0.06u
MN1 VSS M N_40 VPW NCH W=0.305u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.42u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.42u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.42u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.61u L=0.06u
.ENDS PREICGX3P5BA10TR

****
.SUBCKT PREICGX4BA10TR VDD VSS VPW VNW ECK CK E SE
MNA2 NEN SE VSS VPW NCH W=0.185u L=0.06u
MPA2 VDD SE N_2 VNW PCH W=0.645u L=0.06u
MPA1023 NEN E N_2 VNW PCH W=0.23u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.185u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.185u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.185u L=0.06u
MPOEN07 N_18 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_33 CK NM VPW NCH W=0.15u L=0.06u
MNA1 VSS M N_33 VPW NCH W=0.15u L=0.06u
MPA1 N_18 M VDD VNW PCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.25u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.31u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MN1_2 N_41 M VSS VPW NCH W=0.34u L=0.06u
MN0_2 NOUT CK N_41 VPW NCH W=0.34u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.41u L=0.06u
MN0 N_39 CK NOUT VPW NCH W=0.34u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.41u L=0.06u
MN1 VSS M N_39 VPW NCH W=0.34u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.48u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.48u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.48u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS PREICGX4BA10TR

****
.SUBCKT PREICGX5BA10TR VDD VSS VPW VNW ECK CK E SE
MNA2 NEN SE VSS VPW NCH W=0.22u L=0.06u
MPA2 VDD SE N_2 VNW PCH W=0.7u L=0.06u
MPA1023 NEN E N_2 VNW PCH W=0.275u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.22u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.22u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.22u L=0.06u
MPOEN07 N_22 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_49 CK NM VPW NCH W=0.15u L=0.06u
MNA1 N_49 M VSS VPW NCH W=0.15u L=0.06u
MPA1 N_22 M VDD VNW PCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.3u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.37u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MN1_2 N_42 M VSS VPW NCH W=0.43u L=0.06u
MN0_2 NOUT CK N_42 VPW NCH W=0.43u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN0 N_40 CK NOUT VPW NCH W=0.43u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN1 VSS M N_40 VPW NCH W=0.43u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS PREICGX5BA10TR

****
.SUBCKT PREICGX6BA10TR VDD VSS VPW VNW ECK CK E SE
MNA2 NEN SE VSS VPW NCH W=0.24u L=0.06u
MPA2 VDD SE N_6 VNW PCH W=0.7u L=0.06u
MPA1023 NEN E N_6 VNW PCH W=0.3u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.24u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.24u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.24u L=0.06u
MPOEN07 N_10 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 NM CK N_36 VPW NCH W=0.15u L=0.06u
MNA1 N_36 M VSS VPW NCH W=0.15u L=0.06u
MPA1 N_10 M VDD VNW PCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.33u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.41u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MN1 N_46 M VSS VPW NCH W=0.51u L=0.06u
MN0 NOUT CK N_46 VPW NCH W=0.51u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.615u L=0.06u
MN0_2 N_44 CK NOUT VPW NCH W=0.51u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.615u L=0.06u
MN1_2 VSS M N_44 VPW NCH W=0.51u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.15u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.435u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.435u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.43u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS PREICGX6BA10TR

****
.SUBCKT PREICGX7P5BA10TR VDD VSS VPW VNW ECK CK E SE
MPA2_2 VDD SE N_17 VNW PCH W=0.405u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.285u L=0.06u
MPA2 VDD SE N_17 VNW PCH W=0.405u L=0.06u
MPA1023 N_17 E NEN VNW PCH W=0.36u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.285u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.285u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.285u L=0.06u
MPOEN07 N_22 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 NM CK N_44 VPW NCH W=0.15u L=0.06u
MNA1 VSS M N_44 VPW NCH W=0.15u L=0.06u
MPA1 N_22 M VDD VNW PCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.39u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.485u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.15u L=0.06u
MN1_2 N_55 M VSS VPW NCH W=0.43u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.2u L=0.06u
MN0_2 NOUT CK N_55 VPW NCH W=0.43u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN0_3 N_57 CK NOUT VPW NCH W=0.43u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MN1_3 VSS M N_57 VPW NCH W=0.43u L=0.06u
MN1 VSS M N_53 VPW NCH W=0.43u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.16u L=0.06u
MN0 N_53 CK NOUT VPW NCH W=0.43u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.52u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.76u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.45u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.69u L=0.06u
.ENDS PREICGX7P5BA10TR

****
.SUBCKT PREICGX9BA10TR VDD VSS VPW VNW ECK CK E SE
MPA2_2 VDD SE N_4 VNW PCH W=0.465u L=0.06u
MNA2 NEN SE VSS VPW NCH W=0.33u L=0.06u
MPA2 VDD SE N_4 VNW PCH W=0.465u L=0.06u
MPA1023 N_4 E NEN VNW PCH W=0.41u L=0.06u
MNA1020 NEN E VSS VPW NCH W=0.33u L=0.06u
MPOEN NM CK NEN VNW PCH W=0.33u L=0.06u
MNOE NM NCLK_ NEN VPW NCH W=0.33u L=0.06u
MPOEN07 N_30 NCLK_ NM VNW PCH W=0.15u L=0.06u
MNOE05 N_75 CK NM VPW NCH W=0.15u L=0.06u
MNA1 N_75 M VSS VPW NCH W=0.15u L=0.06u
MPA1 N_30 M VDD VNW PCH W=0.15u L=0.06u
MNA1016 M NM VSS VPW NCH W=0.45u L=0.06u
MPA1018 M NM VDD VNW PCH W=0.56u L=0.06u
MNA1012 NCLK_ CK VSS VPW NCH W=0.17u L=0.06u
MN1 N_65 M VSS VPW NCH W=0.515u L=0.06u
MPA1014 NCLK_ CK VDD VNW PCH W=0.225u L=0.06u
MN0 NOUT CK N_65 VPW NCH W=0.515u L=0.06u
MP1_3 NOUT CK VDD VNW PCH W=0.62u L=0.06u
MN0_2 N_67 CK NOUT VPW NCH W=0.515u L=0.06u
MP1_2 NOUT CK VDD VNW PCH W=0.62u L=0.06u
MN1_2 VSS M N_67 VPW NCH W=0.515u L=0.06u
MN1_3 VSS M N_63 VPW NCH W=0.515u L=0.06u
MP0 NOUT M VDD VNW PCH W=0.19u L=0.06u
MN0_3 N_63 CK NOUT VPW NCH W=0.515u L=0.06u
MP1 NOUT CK VDD VNW PCH W=0.62u L=0.06u
MNA1026_5 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_2 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_3 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_8 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_6 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026_8 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_5 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026_7 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_4 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026_6 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_3 ECK NOUT VDD VNW PCH W=0.84u L=0.06u
MNA1026_4 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
MNA1026_2 ECK NOUT VSS VPW NCH W=0.405u L=0.06u
MPA1028_7 ECK NOUT VDD VNW PCH W=0.7u L=0.06u
.ENDS PREICGX9BA10TR

****
.SUBCKT TIEHIX1MA10TR VDD VSS VPW VNW Y
MN1 LO HI VSS VPW NCH W=0.15u L=0.06u
MP1 HI LO VDD VNW PCH W=0.15u L=0.06u
MN0 LO LO VSS VPW NCH W=0.15u L=0.06u
MP0 Y LO VDD VNW PCH W=0.7u L=0.06u
.ENDS TIEHIX1MA10TR

****
.SUBCKT TIELOX1MA10TR VDD VSS VPW VNW Y
MN1 LO HI VSS VPW NCH W=0.15u L=0.06u
MP1 HI LO VDD VNW PCH W=0.15u L=0.06u
MN0 Y HI VSS VPW NCH W=0.55u L=0.06u
MP0 HI HI VDD VNW PCH W=0.15u L=0.06u
.ENDS TIELOX1MA10TR
