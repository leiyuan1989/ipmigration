* SPICE INPUT		Tue Jul 31 18:28:43 2018	ad01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d0
.subckt ad01d0 VDD CO S GND CI B A
M1 S N_15 GND GND mn15  l=0.13u w=0.26u m=1
M2 CO N_12 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.27u m=1
M4 N_69 N_6 GND GND mn15  l=0.13u w=0.27u m=1
M5 N_69 N_11 N_5 GND mn15  l=0.13u w=0.27u m=1
M6 N_5 B N_6 GND mn15  l=0.13u w=0.27u m=1
M7 N_11 B GND GND mn15  l=0.13u w=0.27u m=1
M8 GND N_5 N_10 GND mn15  l=0.13u w=0.27u m=1
M9 N_13 N_5 N_12 GND mn15  l=0.13u w=0.27u m=1
M10 N_11 N_10 N_12 GND mn15  l=0.13u w=0.27u m=1
M11 N_10 N_13 N_15 GND mn15  l=0.13u w=0.27u m=1
M12 N_5 CI N_15 GND mn15  l=0.13u w=0.27u m=1
M13 N_13 CI GND GND mn15  l=0.13u w=0.27u m=1
M14 S N_15 VDD VDD mp15  l=0.13u w=0.4u m=1
M15 CO N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_20 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_6 N_11 N_5 VDD mp15  l=0.13u w=0.27u m=1
M19 N_20 B N_5 VDD mp15  l=0.13u w=0.4u m=1
M20 N_11 B VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_10 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 N_11 N_5 N_12 VDD mp15  l=0.13u w=0.27u m=1
M23 N_13 N_10 N_12 VDD mp15  l=0.13u w=0.27u m=1
M24 N_5 N_13 N_15 VDD mp15  l=0.13u w=0.27u m=1
M25 N_10 CI N_15 VDD mp15  l=0.13u w=0.27u m=1
M26 N_13 CI VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ad01d0
* SPICE INPUT		Tue Jul 31 18:28:58 2018	ad01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d1
.subckt ad01d1 GND S CO CI VDD B A
M1 N_2 A GND GND mn15  l=0.13u w=0.38u m=1
M2 N_20 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_20 N_8 N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B N_2 GND mn15  l=0.13u w=0.33u m=1
M5 N_8 B GND GND mn15  l=0.13u w=0.38u m=1
M6 GND N_3 N_6 GND mn15  l=0.13u w=0.38u m=1
M7 N_10 N_3 N_9 GND mn15  l=0.13u w=0.27u m=1
M8 N_8 N_6 N_9 GND mn15  l=0.13u w=0.27u m=1
M9 N_6 N_10 N_12 GND mn15  l=0.13u w=0.27u m=1
M10 N_3 CI N_12 GND mn15  l=0.13u w=0.27u m=1
M11 GND CI N_10 GND mn15  l=0.13u w=0.37u m=1
M12 S N_12 GND GND mn15  l=0.13u w=0.43u m=1
M13 CO N_9 GND GND mn15  l=0.13u w=0.46u m=1
M14 VDD A N_2 VDD mp15  l=0.13u w=0.53u m=1
M15 N_73 N_2 VDD VDD mp15  l=0.13u w=0.66u m=1
M16 N_2 N_8 N_3 VDD mp15  l=0.13u w=0.315u m=1
M17 N_73 B N_3 VDD mp15  l=0.13u w=0.66u m=1
M18 N_8 B VDD VDD mp15  l=0.13u w=0.53u m=1
M19 N_6 N_3 VDD VDD mp15  l=0.13u w=0.53u m=1
M20 N_8 N_3 N_9 VDD mp15  l=0.13u w=0.27u m=1
M21 N_10 N_6 N_9 VDD mp15  l=0.13u w=0.27u m=1
M22 N_3 N_10 N_12 VDD mp15  l=0.13u w=0.27u m=1
M23 N_6 CI N_12 VDD mp15  l=0.13u w=0.27u m=1
M24 N_10 CI VDD VDD mp15  l=0.13u w=0.27u m=1
M25 VDD CI N_10 VDD mp15  l=0.13u w=0.26u m=1
M26 S N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 CO N_9 VDD VDD mp15  l=0.13u w=0.35u m=1
M28 CO N_9 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends ad01d1
* SPICE INPUT		Tue Jul 31 18:29:15 2018	ad01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d2
.subckt ad01d2 VDD S CO GND CI B A
M1 N_3 B N_2 GND mn15  l=0.13u w=0.36u m=1
M2 N_29 N_9 N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.4u m=1
M4 N_29 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_9 N_8 N_19 GND mn15  l=0.13u w=0.36u m=1
M6 N_19 N_3 N_15 GND mn15  l=0.13u w=0.36u m=1
M7 N_8 N_15 N_11 GND mn15  l=0.13u w=0.18u m=1
M8 N_11 N_15 N_8 GND mn15  l=0.13u w=0.18u m=1
M9 N_3 CI N_11 GND mn15  l=0.13u w=0.35u m=1
M10 GND CI N_15 GND mn15  l=0.13u w=0.2u m=1
M11 N_15 CI GND GND mn15  l=0.13u w=0.2u m=1
M12 GND N_11 S GND mn15  l=0.13u w=0.46u m=1
M13 GND N_11 S GND mn15  l=0.13u w=0.46u m=1
M14 GND N_19 CO GND mn15  l=0.13u w=0.46u m=1
M15 CO N_19 GND GND mn15  l=0.13u w=0.46u m=1
M16 N_8 N_3 GND GND mn15  l=0.13u w=0.41u m=1
M17 N_9 B GND GND mn15  l=0.13u w=0.4u m=1
M18 N_23 B N_3 VDD mp15  l=0.13u w=0.66u m=1
M19 N_3 N_9 N_2 VDD mp15  l=0.13u w=0.27u m=1
M20 N_3 N_9 N_2 VDD mp15  l=0.13u w=0.26u m=1
M21 VDD A N_2 VDD mp15  l=0.13u w=0.59u m=1
M22 N_23 N_2 VDD VDD mp15  l=0.13u w=0.66u m=1
M23 N_8 N_3 VDD VDD mp15  l=0.13u w=0.56u m=1
M24 N_9 B VDD VDD mp15  l=0.13u w=0.56u m=1
M25 N_11 CI N_8 VDD mp15  l=0.13u w=0.53u m=1
M26 N_15 CI VDD VDD mp15  l=0.13u w=0.59u m=1
M27 VDD N_11 S VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_11 S VDD mp15  l=0.13u w=0.69u m=1
M29 CO N_19 VDD VDD mp15  l=0.13u w=0.68u m=1
M30 VDD N_19 CO VDD mp15  l=0.13u w=0.69u m=1
M31 N_9 N_3 N_19 VDD mp15  l=0.13u w=0.53u m=1
M32 N_19 N_8 N_15 VDD mp15  l=0.13u w=0.53u m=1
M33 N_3 N_15 N_11 VDD mp15  l=0.13u w=0.49u m=1
.ends ad01d2
* SPICE INPUT		Tue Jul 31 18:29:28 2018	ad01d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d3
.subckt ad01d3 VDD S CO GND CI B A
M1 N_2 A GND GND mn15  l=0.13u w=0.4u m=1
M2 N_92 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_92 N_9 N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B N_2 GND mn15  l=0.13u w=0.36u m=1
M5 N_9 B GND GND mn15  l=0.13u w=0.4u m=1
M6 N_8 N_3 GND GND mn15  l=0.13u w=0.45u m=1
M7 S N_18 GND GND mn15  l=0.13u w=0.46u m=1
M8 S N_18 GND GND mn15  l=0.13u w=0.46u m=1
M9 S N_18 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_14 N_3 N_15 GND mn15  l=0.13u w=0.36u m=1
M11 N_9 N_8 N_14 GND mn15  l=0.13u w=0.36u m=1
M12 N_3 CI N_18 GND mn15  l=0.13u w=0.35u m=1
M13 N_8 N_15 N_18 GND mn15  l=0.13u w=0.19u m=1
M14 N_18 N_15 N_8 GND mn15  l=0.13u w=0.17u m=1
M15 CO N_14 GND GND mn15  l=0.13u w=0.46u m=1
M16 CO N_14 GND GND mn15  l=0.13u w=0.46u m=1
M17 CO N_14 GND GND mn15  l=0.13u w=0.46u m=1
M18 GND CI N_15 GND mn15  l=0.13u w=0.21u m=1
M19 N_15 CI GND GND mn15  l=0.13u w=0.19u m=1
M20 VDD A N_2 VDD mp15  l=0.13u w=0.58u m=1
M21 N_26 N_2 VDD VDD mp15  l=0.13u w=0.66u m=1
M22 N_3 N_9 N_2 VDD mp15  l=0.13u w=0.27u m=1
M23 N_3 N_9 N_2 VDD mp15  l=0.13u w=0.26u m=1
M24 N_26 B N_3 VDD mp15  l=0.13u w=0.66u m=1
M25 N_9 B VDD VDD mp15  l=0.13u w=0.56u m=1
M26 N_8 N_3 VDD VDD mp15  l=0.13u w=0.56u m=1
M27 S N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 S N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 S N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 N_9 N_3 N_14 VDD mp15  l=0.13u w=0.53u m=1
M31 N_15 N_8 N_14 VDD mp15  l=0.13u w=0.53u m=1
M32 N_18 N_15 N_3 VDD mp15  l=0.13u w=0.49u m=1
M33 N_18 CI N_8 VDD mp15  l=0.13u w=0.53u m=1
M34 CO N_14 VDD VDD mp15  l=0.13u w=0.71u m=1
M35 CO N_14 VDD VDD mp15  l=0.13u w=0.71u m=1
M36 CO N_14 VDD VDD mp15  l=0.13u w=0.65u m=1
M37 N_15 CI VDD VDD mp15  l=0.13u w=0.59u m=1
.ends ad01d3
* SPICE INPUT		Tue Jul 31 18:29:41 2018	ad01dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01dm
.subckt ad01dm GND S CO CI VDD B A
M1 S N_17 GND GND mn15  l=0.13u w=0.35u m=1
M2 CO N_14 GND GND mn15  l=0.13u w=0.35u m=1
M3 N_6 CI GND GND mn15  l=0.13u w=0.31u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.31u m=1
M5 N_20 N_7 GND GND mn15  l=0.13u w=0.31u m=1
M6 N_20 N_13 N_8 GND mn15  l=0.13u w=0.31u m=1
M7 N_8 B N_7 GND mn15  l=0.13u w=0.29u m=1
M8 N_13 B GND GND mn15  l=0.13u w=0.31u m=1
M9 GND N_8 N_11 GND mn15  l=0.13u w=0.31u m=1
M10 N_6 N_8 N_14 GND mn15  l=0.13u w=0.29u m=1
M11 N_13 N_11 N_14 GND mn15  l=0.13u w=0.29u m=1
M12 N_11 N_6 N_17 GND mn15  l=0.13u w=0.29u m=1
M13 N_8 CI N_17 GND mn15  l=0.13u w=0.29u m=1
M14 S N_17 VDD VDD mp15  l=0.13u w=0.53u m=1
M15 CO N_14 VDD VDD mp15  l=0.13u w=0.52u m=1
M16 N_6 CI VDD VDD mp15  l=0.13u w=0.48u m=1
M17 N_7 A VDD VDD mp15  l=0.13u w=0.48u m=1
M18 N_27 N_7 VDD VDD mp15  l=0.13u w=0.45u m=1
M19 N_7 N_13 N_8 VDD mp15  l=0.13u w=0.31u m=1
M20 N_27 B N_8 VDD mp15  l=0.13u w=0.45u m=1
M21 N_13 B VDD VDD mp15  l=0.13u w=0.48u m=1
M22 N_11 N_8 VDD VDD mp15  l=0.13u w=0.48u m=1
M23 N_13 N_8 N_14 VDD mp15  l=0.13u w=0.35u m=1
M24 N_6 N_11 N_14 VDD mp15  l=0.13u w=0.35u m=1
M25 N_8 N_6 N_17 VDD mp15  l=0.13u w=0.29u m=1
M26 N_11 CI N_17 VDD mp15  l=0.13u w=0.29u m=1
.ends ad01dm
* SPICE INPUT		Tue Jul 31 18:29:53 2018	adfh01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=adfh01d0
.subckt adfh01d0 GND S CO A B CI VDD
M1 CO N_13 GND GND mn15  l=0.13u w=0.26u m=1
M2 S N_8 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND CI N_5 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M5 N_8 N_14 N_7 GND mn15  l=0.13u w=0.28u m=1
M6 N_13 N_20 N_11 GND mn15  l=0.13u w=0.28u m=1
M7 N_8 N_20 N_5 GND mn15  l=0.13u w=0.28u m=1
M8 N_13 N_14 N_5 GND mn15  l=0.13u w=0.28u m=1
M9 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M10 N_15 N_11 N_14 GND mn15  l=0.13u w=0.3u m=1
M11 N_20 B N_15 GND mn15  l=0.13u w=0.3u m=1
M12 N_14 B N_16 GND mn15  l=0.13u w=0.28u m=1
M13 N_20 N_11 N_16 GND mn15  l=0.13u w=0.28u m=1
M14 N_15 N_21 GND GND mn15  l=0.13u w=0.36u m=1
M15 N_16 A GND GND mn15  l=0.13u w=0.3u m=1
M16 GND A N_21 GND mn15  l=0.13u w=0.18u m=1
M17 CO N_13 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 S N_8 VDD VDD mp15  l=0.13u w=0.4u m=1
M19 VDD CI N_5 VDD mp15  l=0.13u w=0.35u m=1
M20 VDD N_5 N_7 VDD mp15  l=0.13u w=0.35u m=1
M21 N_5 N_14 N_8 VDD mp15  l=0.13u w=0.28u m=1
M22 N_13 N_14 N_11 VDD mp15  l=0.13u w=0.28u m=1
M23 N_7 N_20 N_8 VDD mp15  l=0.13u w=0.28u m=1
M24 N_5 N_20 N_13 VDD mp15  l=0.13u w=0.28u m=1
M25 N_11 B VDD VDD mp15  l=0.13u w=0.35u m=1
M26 VDD B N_11 VDD mp15  l=0.13u w=0.35u m=1
M27 N_16 B N_20 VDD mp15  l=0.13u w=0.4u m=1
M28 N_14 B N_15 VDD mp15  l=0.13u w=0.4u m=1
M29 N_14 N_11 N_16 VDD mp15  l=0.13u w=0.57u m=1
M30 N_20 N_11 N_15 VDD mp15  l=0.13u w=0.56u m=1
M31 N_15 N_21 VDD VDD mp15  l=0.13u w=0.53u m=1
M32 N_21 A VDD VDD mp15  l=0.13u w=0.3u m=1
M33 N_16 A VDD VDD mp15  l=0.13u w=0.46u m=1
.ends adfh01d0
* SPICE INPUT		Tue Jul 31 18:30:06 2018	adfh01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=adfh01d1
.subckt adfh01d1 GND S CO A B CI VDD
M1 N_4 A GND GND mn15  l=0.13u w=0.41u m=1
M2 N_3 A GND GND mn15  l=0.13u w=0.27u m=1
M3 N_8 N_3 GND GND mn15  l=0.13u w=0.41u m=1
M4 N_9 B N_8 GND mn15  l=0.13u w=0.27u m=1
M5 N_6 B N_4 GND mn15  l=0.13u w=0.27u m=1
M6 N_9 N_19 N_4 GND mn15  l=0.13u w=0.27u m=1
M7 CO N_21 GND GND mn15  l=0.13u w=0.46u m=1
M8 S N_16 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND CI N_13 GND mn15  l=0.13u w=0.41u m=1
M10 N_15 N_13 GND GND mn15  l=0.13u w=0.41u m=1
M11 N_16 N_6 N_15 GND mn15  l=0.13u w=0.27u m=1
M12 N_21 N_9 N_19 GND mn15  l=0.13u w=0.27u m=1
M13 N_16 N_9 N_13 GND mn15  l=0.13u w=0.27u m=1
M14 N_21 N_6 N_13 GND mn15  l=0.13u w=0.27u m=1
M15 GND B N_19 GND mn15  l=0.13u w=0.46u m=1
M16 N_8 N_19 N_6 GND mn15  l=0.13u w=0.27u m=1
M17 CO N_21 VDD VDD mp15  l=0.13u w=0.35u m=1
M18 CO N_21 VDD VDD mp15  l=0.13u w=0.35u m=1
M19 S N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_4 A VDD VDD mp15  l=0.13u w=0.59u m=1
M21 N_3 A VDD VDD mp15  l=0.13u w=0.35u m=1
M22 VDD CI N_13 VDD mp15  l=0.13u w=0.59u m=1
M23 VDD N_13 N_15 VDD mp15  l=0.13u w=0.59u m=1
M24 N_13 N_6 N_16 VDD mp15  l=0.13u w=0.4u m=1
M25 N_21 N_6 N_19 VDD mp15  l=0.13u w=0.4u m=1
M26 N_15 N_9 N_16 VDD mp15  l=0.13u w=0.4u m=1
M27 N_13 N_9 N_21 VDD mp15  l=0.13u w=0.4u m=1
M28 N_19 B VDD VDD mp15  l=0.13u w=0.35u m=1
M29 VDD B N_19 VDD mp15  l=0.13u w=0.35u m=1
M30 N_8 N_3 VDD VDD mp15  l=0.13u w=0.59u m=1
M31 N_4 B N_9 VDD mp15  l=0.13u w=0.4u m=1
M32 N_6 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M33 N_6 N_19 N_4 VDD mp15  l=0.13u w=0.4u m=1
M34 N_9 N_19 N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends adfh01d1
* SPICE INPUT		Tue Jul 31 18:30:19 2018	adfh01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=adfh01d2
.subckt adfh01d2 S GND CO VDD CI B A
M1 CO N_26 GND GND mn15  l=0.13u w=0.46u m=1
M2 GND N_26 CO GND mn15  l=0.13u w=0.46u m=1
M3 GND N_10 S GND mn15  l=0.13u w=0.46u m=1
M4 GND N_10 S GND mn15  l=0.13u w=0.46u m=1
M5 GND CI N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_10 N_14 N_9 GND mn15  l=0.13u w=0.41u m=1
M7 N_9 N_7 GND GND mn15  l=0.13u w=0.4u m=1
M8 N_13 A GND GND mn15  l=0.13u w=0.38u m=1
M9 N_12 A GND GND mn15  l=0.13u w=0.27u m=1
M10 N_17 N_12 GND GND mn15  l=0.13u w=0.4u m=1
M11 N_18 B N_17 GND mn15  l=0.13u w=0.41u m=1
M12 N_13 B N_14 GND mn15  l=0.13u w=0.41u m=1
M13 N_18 N_23 N_13 GND mn15  l=0.13u w=0.41u m=1
M14 N_14 N_23 N_17 GND mn15  l=0.13u w=0.41u m=1
M15 GND B N_23 GND mn15  l=0.13u w=0.235u m=1
M16 N_23 B GND GND mn15  l=0.13u w=0.225u m=1
M17 N_26 N_14 N_7 GND mn15  l=0.13u w=0.41u m=1
M18 N_7 N_18 N_10 GND mn15  l=0.13u w=0.41u m=1
M19 N_26 N_18 N_23 GND mn15  l=0.13u w=0.41u m=1
M20 N_13 A VDD VDD mp15  l=0.13u w=0.56u m=1
M21 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M22 VDD N_26 CO VDD mp15  l=0.13u w=0.47u m=1
M23 CO N_26 VDD VDD mp15  l=0.13u w=0.47u m=1
M24 VDD N_26 CO VDD mp15  l=0.13u w=0.46u m=1
M25 VDD N_10 S VDD mp15  l=0.13u w=0.69u m=1
M26 VDD N_10 S VDD mp15  l=0.13u w=0.69u m=1
M27 N_17 N_12 VDD VDD mp15  l=0.13u w=0.59u m=1
M28 N_17 N_23 N_18 VDD mp15  l=0.13u w=0.31u m=1
M29 N_17 N_23 N_18 VDD mp15  l=0.13u w=0.31u m=1
M30 N_18 B N_13 VDD mp15  l=0.13u w=0.62u m=1
M31 N_13 N_23 N_14 VDD mp15  l=0.13u w=0.62u m=1
M32 N_17 B N_14 VDD mp15  l=0.13u w=0.62u m=1
M33 VDD B N_23 VDD mp15  l=0.13u w=0.35u m=1
M34 VDD B N_23 VDD mp15  l=0.13u w=0.35u m=1
M35 N_23 N_14 N_26 VDD mp15  l=0.13u w=0.31u m=1
M36 N_23 N_14 N_26 VDD mp15  l=0.13u w=0.31u m=1
M37 N_7 N_18 N_26 VDD mp15  l=0.13u w=0.62u m=1
M38 N_10 N_18 N_9 VDD mp15  l=0.13u w=0.62u m=1
M39 N_7 N_14 N_10 VDD mp15  l=0.13u w=0.62u m=1
M40 N_7 CI VDD VDD mp15  l=0.13u w=0.59u m=1
M41 N_9 N_7 VDD VDD mp15  l=0.13u w=0.59u m=1
.ends adfh01d2
* SPICE INPUT		Tue Jul 31 18:30:31 2018	ah01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d0
.subckt ah01d0 GND CO S VDD A B
M1 N_12 B GND GND mn15  l=0.13u w=0.26u m=1
M2 CO N_4 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_12 A N_4 GND mn15  l=0.13u w=0.26u m=1
M4 N_11 B N_9 GND mn15  l=0.13u w=0.26u m=1
M5 N_6 B GND GND mn15  l=0.13u w=0.26u m=1
M6 N_9 N_10 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_11 N_6 N_10 GND mn15  l=0.13u w=0.26u m=1
M8 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M9 GND N_11 S GND mn15  l=0.13u w=0.26u m=1
M10 N_4 B VDD VDD mp15  l=0.13u w=0.4u m=1
M11 CO N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_10 B N_11 VDD mp15  l=0.13u w=0.4u m=1
M14 N_6 B VDD VDD mp15  l=0.13u w=0.4u m=1
M15 N_9 N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_9 N_6 N_11 VDD mp15  l=0.13u w=0.4u m=1
M17 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M18 S N_11 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ah01d0
* SPICE INPUT		Tue Jul 31 18:30:44 2018	ah01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d1
.subckt ah01d1 GND S CO A VDD B
M1 S N_8 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_8 B N_6 GND mn15  l=0.13u w=0.28u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.26u m=1
M4 N_6 N_7 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 N_3 N_7 GND mn15  l=0.13u w=0.28u m=1
M6 N_7 A GND GND mn15  l=0.13u w=0.31u m=1
M7 CO N_11 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_12 B GND GND mn15  l=0.13u w=0.28u m=1
M9 N_12 A N_11 GND mn15  l=0.13u w=0.28u m=1
M10 S N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_7 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M12 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_6 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_8 N_3 N_6 VDD mp15  l=0.13u w=0.38u m=1
M15 N_7 A VDD VDD mp15  l=0.13u w=0.46u m=1
M16 CO N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_11 B VDD VDD mp15  l=0.13u w=0.28u m=1
M18 N_11 A VDD VDD mp15  l=0.13u w=0.28u m=1
.ends ah01d1
* SPICE INPUT		Tue Jul 31 18:31:00 2018	ah01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d2
.subckt ah01d2 GND S CO VDD A B
M1 N_3 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_8 B N_7 GND mn15  l=0.13u w=0.31u m=1
M3 S N_8 GND GND mn15  l=0.13u w=0.46u m=1
M4 S N_8 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_9 N_3 N_8 GND mn15  l=0.13u w=0.36u m=1
M6 N_9 A GND GND mn15  l=0.13u w=0.33u m=1
M7 N_7 N_9 GND GND mn15  l=0.13u w=0.31u m=1
M8 N_14 B GND GND mn15  l=0.13u w=0.47u m=1
M9 N_14 A N_12 GND mn15  l=0.13u w=0.47u m=1
M10 GND N_12 CO GND mn15  l=0.13u w=0.46u m=1
M11 GND N_12 CO GND mn15  l=0.13u w=0.46u m=1
M12 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_9 B N_8 VDD mp15  l=0.13u w=0.52u m=1
M14 S N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 S N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_9 A VDD VDD mp15  l=0.13u w=0.51u m=1
M17 N_7 N_9 VDD VDD mp15  l=0.13u w=0.48u m=1
M18 N_8 N_3 N_7 VDD mp15  l=0.13u w=0.48u m=1
M19 VDD B N_12 VDD mp15  l=0.13u w=0.52u m=1
M20 N_12 A VDD VDD mp15  l=0.13u w=0.26u m=1
M21 N_12 A VDD VDD mp15  l=0.13u w=0.26u m=1
M22 VDD N_12 CO VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_12 CO VDD mp15  l=0.13u w=0.69u m=1
.ends ah01d2
* SPICE INPUT		Tue Jul 31 18:31:18 2018	ah01d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d3
.subckt ah01d3 GND CO S VDD A B
M1 GND B N_25 GND mn15  l=0.13u w=0.45u m=1
M2 N_24 B GND GND mn15  l=0.13u w=0.21u m=1
M3 GND B N_4 GND mn15  l=0.13u w=0.28u m=1
M4 N_6 A N_25 GND mn15  l=0.13u w=0.36u m=1
M5 N_6 A N_24 GND mn15  l=0.13u w=0.36u m=1
M6 CO N_6 GND GND mn15  l=0.13u w=0.46u m=1
M7 CO N_6 GND GND mn15  l=0.13u w=0.46u m=1
M8 CO N_6 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_13 S GND mn15  l=0.13u w=0.46u m=1
M10 GND N_13 S GND mn15  l=0.13u w=0.46u m=1
M11 GND N_13 S GND mn15  l=0.13u w=0.46u m=1
M12 N_14 B N_13 GND mn15  l=0.13u w=0.27u m=1
M13 N_13 B N_14 GND mn15  l=0.13u w=0.27u m=1
M14 GND N_20 N_14 GND mn15  l=0.13u w=0.25u m=1
M15 N_14 N_20 GND GND mn15  l=0.13u w=0.24u m=1
M16 N_20 N_4 N_13 GND mn15  l=0.13u w=0.27u m=1
M17 N_13 N_4 N_20 GND mn15  l=0.13u w=0.27u m=1
M18 N_20 A GND GND mn15  l=0.13u w=0.3u m=1
M19 N_20 A GND GND mn15  l=0.13u w=0.3u m=1
M20 VDD N_13 S VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_13 S VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_13 S VDD mp15  l=0.13u w=0.69u m=1
M23 VDD B N_6 VDD mp15  l=0.13u w=0.41u m=1
M24 N_6 B VDD VDD mp15  l=0.13u w=0.41u m=1
M25 VDD B N_4 VDD mp15  l=0.13u w=0.4u m=1
M26 N_6 A VDD VDD mp15  l=0.13u w=0.41u m=1
M27 VDD A N_6 VDD mp15  l=0.13u w=0.39u m=1
M28 CO N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 CO N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 CO N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 N_13 N_4 N_14 VDD mp15  l=0.13u w=0.37u m=1
M32 N_13 N_4 N_14 VDD mp15  l=0.13u w=0.325u m=1
M33 N_14 N_20 VDD VDD mp15  l=0.13u w=0.33u m=1
M34 VDD N_20 N_14 VDD mp15  l=0.13u w=0.33u m=1
M35 N_20 B N_13 VDD mp15  l=0.13u w=0.36u m=1
M36 N_20 B N_13 VDD mp15  l=0.13u w=0.34u m=1
M37 VDD A N_20 VDD mp15  l=0.13u w=0.5u m=1
M38 N_20 A VDD VDD mp15  l=0.13u w=0.5u m=1
.ends ah01d3
* SPICE INPUT		Tue Jul 31 18:31:30 2018	ah01dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01dm
.subckt ah01dm GND S CO A VDD B
M1 S N_8 GND GND mn15  l=0.13u w=0.35u m=1
M2 N_8 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.26u m=1
M4 N_6 N_7 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 N_3 N_7 GND mn15  l=0.13u w=0.26u m=1
M6 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M7 CO N_11 GND GND mn15  l=0.13u w=0.35u m=1
M8 N_12 B GND GND mn15  l=0.13u w=0.26u m=1
M9 N_12 A N_11 GND mn15  l=0.13u w=0.26u m=1
M10 S N_8 VDD VDD mp15  l=0.13u w=0.53u m=1
M11 N_7 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M12 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_6 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_8 N_3 N_6 VDD mp15  l=0.13u w=0.4u m=1
M15 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M16 CO N_11 VDD VDD mp15  l=0.13u w=0.53u m=1
M17 N_11 B VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_11 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ah01dm
* SPICE INPUT		Tue Jul 31 18:31:43 2018	an02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d0
.subckt an02d0 GND Y VDD A B
M1 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 B N_4 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M5 N_4 B VDD VDD mp15  l=0.13u w=0.325u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.325u m=1
.ends an02d0
* SPICE INPUT		Tue Jul 31 18:31:57 2018	an02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d1
.subckt an02d1 GND Y VDD A B
M1 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_5 B N_4 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M5 N_4 B VDD VDD mp15  l=0.13u w=0.325u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.325u m=1
.ends an02d1
* SPICE INPUT		Tue Jul 31 18:32:10 2018	an02d1p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d1p5
.subckt an02d1p5 GND Y VDD A B
M1 N_5 B N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an02d1p5
* SPICE INPUT		Tue Jul 31 18:32:22 2018	an02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d2
.subckt an02d2 Y GND VDD A B
M1 GND A N_6 GND mn15  l=0.13u w=0.46u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 N_6 B N_4 GND mn15  l=0.13u w=0.46u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.57u m=1
M6 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M8 N_4 B VDD VDD mp15  l=0.13u w=0.57u m=1
.ends an02d2
* SPICE INPUT		Tue Jul 31 18:32:34 2018	an02d2p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d2p5
.subckt an02d2p5 Y GND VDD A B
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_8 B N_5 GND mn15  l=0.13u w=0.46u m=1
M6 N_5 B N_7 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an02d2p5
* SPICE INPUT		Tue Jul 31 18:32:46 2018	an02d3p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d3p5
.subckt an02d3p5 Y GND VDD A B
M1 N_10 B N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_12 B N_4 GND mn15  l=0.13u w=0.46u m=1
M5 N_4 B N_11 GND mn15  l=0.13u w=0.46u m=1
M6 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M14 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD B N_4 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an02d3p5
* SPICE INPUT		Tue Jul 31 18:32:58 2018	an02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d4
.subckt an02d4 Y GND VDD A B
M1 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_10 B N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_5 B N_9 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_10 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD B N_5 VDD mp15  l=0.13u w=0.345u m=1
M12 VDD A N_5 VDD mp15  l=0.13u w=0.345u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an02d4
* SPICE INPUT		Tue Jul 31 18:33:10 2018	an02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02dm
.subckt an02dm GND Y VDD A B
M1 N_5 B N_4 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_4 B VDD VDD mp15  l=0.13u w=0.325u m=1
M5 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.325u m=1
.ends an02dm
* SPICE INPUT		Tue Jul 31 18:33:22 2018	an03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d0
.subckt an03d0 GND Y VDD A B C
M1 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_5 C N_4 GND mn15  l=0.13u w=0.26u m=1
M5 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.29u m=1
M7 N_4 B VDD VDD mp15  l=0.13u w=0.29u m=1
M8 N_4 C VDD VDD mp15  l=0.13u w=0.29u m=1
.ends an03d0
* SPICE INPUT		Tue Jul 31 18:33:35 2018	an03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d1
.subckt an03d1 GND Y VDD A B C
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C N_4 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.29u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.29u m=1
M7 N_4 C VDD VDD mp15  l=0.13u w=0.29u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an03d1
* SPICE INPUT		Tue Jul 31 18:33:47 2018	an03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d2
.subckt an03d2 Y GND VDD A B C
M1 N_6 C N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 VDD C N_4 VDD mp15  l=0.13u w=0.51u m=1
M7 N_4 B VDD VDD mp15  l=0.13u w=0.51u m=1
M8 VDD A N_4 VDD mp15  l=0.13u w=0.51u m=1
M9 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends an03d2
* SPICE INPUT		Tue Jul 31 18:34:01 2018	an03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d4
.subckt an03d4 Y GND VDD A B C
M1 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_10 B N_9 GND mn15  l=0.13u w=0.46u m=1
M3 N_11 C N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_5 C N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_12 B N_11 GND mn15  l=0.13u w=0.46u m=1
M6 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_5 A VDD VDD mp15  l=0.13u w=0.505u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.505u m=1
M13 N_5 C VDD VDD mp15  l=0.13u w=0.505u m=1
M14 N_5 C VDD VDD mp15  l=0.13u w=0.505u m=1
M15 N_5 B VDD VDD mp15  l=0.13u w=0.505u m=1
M16 VDD A N_5 VDD mp15  l=0.13u w=0.505u m=1
M17 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an03d4
* SPICE INPUT		Tue Jul 31 18:34:17 2018	an03dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03dm
.subckt an03dm GND Y VDD A B C
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C N_4 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.29u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.29u m=1
M7 N_4 C VDD VDD mp15  l=0.13u w=0.29u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends an03dm
* SPICE INPUT		Tue Jul 31 18:34:33 2018	an04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d0
.subckt an04d0 GND Y D C B A VDD
M1 N_5 D N_4 GND mn15  l=0.13u w=0.26u m=1
M2 N_6 C N_5 GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M5 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M6 N_4 D VDD VDD mp15  l=0.13u w=0.26u m=1
M7 VDD C N_4 VDD mp15  l=0.13u w=0.26u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_4 B VDD VDD mp15  l=0.13u w=0.26u m=1
M10 N_4 A VDD VDD mp15  l=0.13u w=0.26u m=1
.ends an04d0
* SPICE INPUT		Tue Jul 31 18:34:47 2018	an04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d1
.subckt an04d1 GND Y VDD A B C D
M1 N_5 D N_4 GND mn15  l=0.13u w=0.36u m=1
M2 N_6 C N_5 GND mn15  l=0.13u w=0.36u m=1
M3 N_7 B N_6 GND mn15  l=0.13u w=0.36u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.36u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_4 D VDD VDD mp15  l=0.13u w=0.36u m=1
M7 N_4 C VDD VDD mp15  l=0.13u w=0.36u m=1
M8 N_4 B VDD VDD mp15  l=0.13u w=0.36u m=1
M9 N_4 A VDD VDD mp15  l=0.13u w=0.36u m=1
M10 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an04d1
* SPICE INPUT		Tue Jul 31 18:35:00 2018	an04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d2
.subckt an04d2 Y GND VDD A B C D
M1 N_6 D N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 C N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_8 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_4 D VDD VDD mp15  l=0.13u w=0.46u m=1
M8 VDD C N_4 VDD mp15  l=0.13u w=0.46u m=1
M9 N_4 B VDD VDD mp15  l=0.13u w=0.46u m=1
M10 VDD A N_4 VDD mp15  l=0.13u w=0.46u m=1
M11 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends an04d2
* SPICE INPUT		Tue Jul 31 18:35:12 2018	an04d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d4
.subckt an04d4 Y GND VDD D C B A
M1 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_8 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_8 GND mn15  l=0.13u w=0.46u m=1
M7 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M8 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 C N_7 GND mn15  l=0.13u w=0.46u m=1
M10 N_7 C N_12 GND mn15  l=0.13u w=0.46u m=1
M11 N_13 D N_12 GND mn15  l=0.13u w=0.46u m=1
M12 N_12 D N_13 GND mn15  l=0.13u w=0.46u m=1
M13 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_13 A VDD VDD mp15  l=0.13u w=0.46u m=1
M18 N_13 A VDD VDD mp15  l=0.13u w=0.46u m=1
M19 N_13 B VDD VDD mp15  l=0.13u w=0.46u m=1
M20 N_13 B VDD VDD mp15  l=0.13u w=0.46u m=1
M21 N_13 C VDD VDD mp15  l=0.13u w=0.46u m=1
M22 N_13 C VDD VDD mp15  l=0.13u w=0.46u m=1
M23 VDD D N_13 VDD mp15  l=0.13u w=0.46u m=1
M24 VDD D N_13 VDD mp15  l=0.13u w=0.46u m=1
.ends an04d4
* SPICE INPUT		Tue Jul 31 18:35:25 2018	an04dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04dm
.subckt an04dm GND Y VDD A B C D
M1 N_7 B N_6 GND mn15  l=0.13u w=0.3u m=1
M2 N_5 D N_4 GND mn15  l=0.13u w=0.3u m=1
M3 N_6 C N_5 GND mn15  l=0.13u w=0.3u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.3u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.3u m=1
M7 N_4 D VDD VDD mp15  l=0.13u w=0.3u m=1
M8 VDD C N_4 VDD mp15  l=0.13u w=0.3u m=1
M9 N_4 A VDD VDD mp15  l=0.13u w=0.3u m=1
M10 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends an04dm
* SPICE INPUT		Wed Aug  1 08:15:11 2018	antenna
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR


* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d0
.subckt aoi211d0 GND Y VDD D C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y D GND GND mn15  l=0.13u w=0.26u m=1
M4 Y C GND GND mn15  l=0.13u w=0.26u m=1
M5 N_11 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_11 B VDD VDD mp15  l=0.13u w=0.4u m=1
M7 Y D N_14 VDD mp15  l=0.13u w=0.4u m=1
M8 N_11 C N_14 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi211d0
* SPICE INPUT		Tue Jul 31 18:35:58 2018	aoi211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d1
.subckt aoi211d1 Y VDD GND D C B A
M1 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y C GND GND mn15  l=0.13u w=0.26u m=1
M4 Y D GND GND mn15  l=0.13u w=0.26u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_4 C N_6 VDD mp15  l=0.13u w=0.69u m=1
M8 Y D N_6 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi211d1
* SPICE INPUT		Tue Jul 31 18:36:12 2018	aoi211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d2
.subckt aoi211d2 GND Y VDD C D A B
M1 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_8 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND C Y GND mn15  l=0.13u w=0.46u m=1
M6 Y D GND GND mn15  l=0.13u w=0.46u m=1
M7 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_12 B VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_12 B VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_18 C N_12 VDD mp15  l=0.13u w=0.69u m=1
M12 Y D N_17 VDD mp15  l=0.13u w=0.69u m=1
M13 Y D N_18 VDD mp15  l=0.13u w=0.69u m=1
M14 N_12 C N_17 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi211d2
* SPICE INPUT		Tue Jul 31 18:36:31 2018	aoi211d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d4
.subckt aoi211d4 GND Y VDD C D A B
M1 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_11 GND mn15  l=0.13u w=0.46u m=1
M4 GND D Y GND mn15  l=0.13u w=0.46u m=1
M5 Y D GND GND mn15  l=0.13u w=0.46u m=1
M6 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_14 B Y GND mn15  l=0.13u w=0.46u m=1
M9 Y B N_13 GND mn15  l=0.13u w=0.46u m=1
M10 Y C GND GND mn15  l=0.13u w=0.46u m=1
M11 Y C GND GND mn15  l=0.13u w=0.46u m=1
M12 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M13 N_20 C N_70 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD B N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_72 D Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y D N_71 VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M20 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD B N_20 VDD mp15  l=0.13u w=0.69u m=1
M22 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_71 C N_20 VDD mp15  l=0.13u w=0.69u m=1
M24 N_73 C N_20 VDD mp15  l=0.13u w=0.69u m=1
M25 N_20 C N_72 VDD mp15  l=0.13u w=0.69u m=1
M26 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 Y D N_70 VDD mp15  l=0.13u w=0.69u m=1
M28 Y D N_73 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi211d4
* SPICE INPUT		Tue Jul 31 18:36:45 2018	aoi21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d0
.subckt aoi21d0 Y VDD GND C B A
M1 N_19 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_19 B Y GND mn15  l=0.13u w=0.26u m=1
M3 Y C GND GND mn15  l=0.13u w=0.26u m=1
M4 VDD A N_2 VDD mp15  l=0.13u w=0.4u m=1
M5 VDD B N_2 VDD mp15  l=0.13u w=0.4u m=1
M6 Y C N_2 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi21d0
* SPICE INPUT		Tue Jul 31 18:36:57 2018	aoi21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d1
.subckt aoi21d1 Y VDD GND C B A
M1 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_19 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y C GND GND mn15  l=0.13u w=0.26u m=1
M4 VDD A N_2 VDD mp15  l=0.13u w=0.69u m=1
M5 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M6 Y C N_2 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21d1
* SPICE INPUT		Tue Jul 31 18:37:09 2018	aoi21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d2
.subckt aoi21d2 GND Y VDD C A B
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M5 Y C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_12 B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_12 B VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21d2
* SPICE INPUT		Tue Jul 31 18:37:22 2018	aoi21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d4
.subckt aoi21d4 GND Y VDD C A B
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_11 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_13 B Y GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_12 GND mn15  l=0.13u w=0.46u m=1
M8 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M9 Y C GND GND mn15  l=0.13u w=0.31u m=1
M10 Y C GND GND mn15  l=0.13u w=0.31u m=1
M11 Y C GND GND mn15  l=0.13u w=0.31u m=1
M12 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD B N_20 VDD mp15  l=0.13u w=0.69u m=1
M14 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD B N_20 VDD mp15  l=0.13u w=0.69u m=1
M18 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Y C N_20 VDD mp15  l=0.13u w=0.85u m=1
M21 Y C N_20 VDD mp15  l=0.13u w=0.69u m=1
M22 Y C N_20 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21d4
* SPICE INPUT		Tue Jul 31 18:37:34 2018	aoi21dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21dm
.subckt aoi21dm Y VDD GND C B A
M1 N_19 A GND GND mn15  l=0.13u w=0.36u m=1
M2 N_19 B Y GND mn15  l=0.13u w=0.36u m=1
M3 Y C GND GND mn15  l=0.13u w=0.26u m=1
M4 VDD A N_2 VDD mp15  l=0.13u w=0.55u m=1
M5 VDD B N_2 VDD mp15  l=0.13u w=0.55u m=1
M6 Y C N_2 VDD mp15  l=0.13u w=0.55u m=1
.ends aoi21dm
* SPICE INPUT		Tue Jul 31 18:37:46 2018	aoi21md0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21md0
.subckt aoi21md0 GND Y VDD A B CN
M1 GND CN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 GND A N_6 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_3 CN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_10 B VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_10 N_3 Y VDD mp15  l=0.13u w=0.4u m=1
.ends aoi21md0
* SPICE INPUT		Tue Jul 31 18:37:57 2018	aoi21md1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21md1
.subckt aoi21md1 GND Y VDD A B CN
M1 N_3 CN GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_7 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 CN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_11 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M7 N_11 B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21md1
* SPICE INPUT		Tue Jul 31 18:38:09 2018	aoi21md2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21md2
.subckt aoi21md2 GND Y VDD A B CN
M1 N_3 CN GND GND mn15  l=0.13u w=0.3u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M4 Y B N_8 GND mn15  l=0.13u w=0.46u m=1
M5 Y B N_9 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_8 GND mn15  l=0.13u w=0.46u m=1
M7 VDD CN N_3 VDD mp15  l=0.13u w=0.45u m=1
M8 N_13 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M9 Y N_3 N_13 VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_13 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21md2
* SPICE INPUT		Tue Jul 31 18:38:21 2018	aoi21md3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21md3
.subckt aoi21md3 GND Y VDD B A CN
M1 N_3 CN GND GND mn15  l=0.13u w=0.46u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.31u m=1
M3 Y N_3 GND GND mn15  l=0.13u w=0.31u m=1
M4 Y N_3 GND GND mn15  l=0.13u w=0.31u m=1
M5 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_14 B Y GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_13 GND mn15  l=0.13u w=0.46u m=1
M8 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M10 Y B N_12 GND mn15  l=0.13u w=0.46u m=1
M11 Y B N_15 GND mn15  l=0.13u w=0.46u m=1
M12 GND A N_12 GND mn15  l=0.13u w=0.46u m=1
M13 N_3 CN VDD VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_3 N_22 VDD mp15  l=0.13u w=0.85u m=1
M15 N_22 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M16 N_22 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_22 VDD mp15  l=0.13u w=0.69u m=1
M18 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD B N_22 VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_22 VDD mp15  l=0.13u w=0.69u m=1
M21 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21md3
* SPICE INPUT		Tue Jul 31 18:38:33 2018	aoi221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d0
.subckt aoi221d0 GND Y VDD E D C A B
M1 N_6 B Y GND mn15  l=0.13u w=0.26u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_7 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 D Y GND mn15  l=0.13u w=0.26u m=1
M5 Y E GND GND mn15  l=0.13u w=0.26u m=1
M6 N_14 B VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_14 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_12 C N_14 VDD mp15  l=0.13u w=0.4u m=1
M9 N_14 D N_12 VDD mp15  l=0.13u w=0.4u m=1
M10 Y E N_12 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi221d0
* SPICE INPUT		Tue Jul 31 18:38:45 2018	aoi221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d1
.subckt aoi221d1 VDD Y GND E D C A B
M1 N_15 B Y GND mn15  l=0.13u w=0.46u m=1
M2 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_16 D Y GND mn15  l=0.13u w=0.46u m=1
M5 Y E GND GND mn15  l=0.13u w=0.26u m=1
M6 N_3 B VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_3 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_3 C N_5 VDD mp15  l=0.13u w=0.69u m=1
M9 N_3 D N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 Y E N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi221d1
* SPICE INPUT		Tue Jul 31 18:38:57 2018	aoi221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d2
.subckt aoi221d2 GND Y VDD E C D A B
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_9 GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_11 D Y GND mn15  l=0.13u w=0.46u m=1
M6 N_12 C GND GND mn15  l=0.13u w=0.46u m=1
M7 N_11 C GND GND mn15  l=0.13u w=0.46u m=1
M8 N_12 D Y GND mn15  l=0.13u w=0.46u m=1
M9 GND E Y GND mn15  l=0.13u w=0.46u m=1
M10 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD B N_22 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD B N_22 VDD mp15  l=0.13u w=0.69u m=1
M13 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_22 D N_19 VDD mp15  l=0.13u w=0.69u m=1
M15 N_22 C N_19 VDD mp15  l=0.13u w=0.69u m=1
M16 N_19 C N_22 VDD mp15  l=0.13u w=0.69u m=1
M17 N_19 D N_22 VDD mp15  l=0.13u w=0.69u m=1
M18 N_19 E Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_19 E Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi221d2
* SPICE INPUT		Tue Jul 31 18:39:09 2018	aoi221d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d4
.subckt aoi221d4 Y GND VDD E C D A B
M1 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_14 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_13 GND mn15  l=0.13u w=0.46u m=1
M4 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_16 B Y GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_15 GND mn15  l=0.13u w=0.46u m=1
M8 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND E Y GND mn15  l=0.13u w=0.46u m=1
M10 GND E Y GND mn15  l=0.13u w=0.46u m=1
M11 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M12 N_18 D Y GND mn15  l=0.13u w=0.46u m=1
M13 Y D N_17 GND mn15  l=0.13u w=0.46u m=1
M14 N_19 C GND GND mn15  l=0.13u w=0.46u m=1
M15 N_18 C GND GND mn15  l=0.13u w=0.46u m=1
M16 N_20 D Y GND mn15  l=0.13u w=0.46u m=1
M17 Y D N_19 GND mn15  l=0.13u w=0.46u m=1
M18 N_20 C GND GND mn15  l=0.13u w=0.46u m=1
M19 N_33 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_33 B VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD B N_33 VDD mp15  l=0.13u w=0.69u m=1
M22 N_33 A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 VDD A N_33 VDD mp15  l=0.13u w=0.69u m=1
M24 VDD B N_33 VDD mp15  l=0.13u w=0.69u m=1
M25 VDD B N_33 VDD mp15  l=0.13u w=0.69u m=1
M26 VDD A N_33 VDD mp15  l=0.13u w=0.69u m=1
M27 N_30 E Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y E N_30 VDD mp15  l=0.13u w=0.69u m=1
M29 N_30 E Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_30 E Y VDD mp15  l=0.13u w=0.69u m=1
M31 N_33 C N_30 VDD mp15  l=0.13u w=0.69u m=1
M32 N_33 D N_30 VDD mp15  l=0.13u w=0.69u m=1
M33 N_30 D N_33 VDD mp15  l=0.13u w=0.69u m=1
M34 N_33 C N_30 VDD mp15  l=0.13u w=0.69u m=1
M35 N_30 C N_33 VDD mp15  l=0.13u w=0.69u m=1
M36 N_33 D N_30 VDD mp15  l=0.13u w=0.69u m=1
M37 N_30 D N_33 VDD mp15  l=0.13u w=0.69u m=1
M38 N_30 C N_33 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi221d4
* SPICE INPUT		Tue Jul 31 18:39:23 2018	aoi222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi222d0
.subckt aoi222d0 Y GND VDD F E C D B A
M1 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y F N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y B N_7 GND mn15  l=0.13u w=0.26u m=1
M4 N_8 D Y GND mn15  l=0.13u w=0.26u m=1
M5 N_8 C GND GND mn15  l=0.13u w=0.26u m=1
M6 GND E N_6 GND mn15  l=0.13u w=0.26u m=1
M7 VDD A N_17 VDD mp15  l=0.13u w=0.4u m=1
M8 VDD B N_17 VDD mp15  l=0.13u w=0.4u m=1
M9 N_14 F Y VDD mp15  l=0.13u w=0.4u m=1
M10 N_17 D N_14 VDD mp15  l=0.13u w=0.4u m=1
M11 N_14 C N_17 VDD mp15  l=0.13u w=0.4u m=1
M12 N_14 E Y VDD mp15  l=0.13u w=0.4u m=1
.ends aoi222d0
* SPICE INPUT		Tue Jul 31 18:39:38 2018	aoi222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi222d1
.subckt aoi222d1 Y GND VDD F E C D B A
M1 Y F N_6 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 D Y GND mn15  l=0.13u w=0.46u m=1
M5 N_8 C GND GND mn15  l=0.13u w=0.46u m=1
M6 GND E N_6 GND mn15  l=0.13u w=0.46u m=1
M7 VDD A N_17 VDD mp15  l=0.13u w=0.69u m=1
M8 VDD B N_17 VDD mp15  l=0.13u w=0.69u m=1
M9 N_14 F Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_17 D N_14 VDD mp15  l=0.13u w=0.69u m=1
M11 N_14 C N_17 VDD mp15  l=0.13u w=0.69u m=1
M12 N_14 E Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi222d1
* SPICE INPUT		Tue Jul 31 18:39:53 2018	aoi222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi222d2
.subckt aoi222d2 GND Y VDD E F C D A B
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_11 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_12 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_13 D Y GND mn15  l=0.13u w=0.46u m=1
M7 Y D N_12 GND mn15  l=0.13u w=0.46u m=1
M8 N_13 C GND GND mn15  l=0.13u w=0.46u m=1
M9 N_14 E GND GND mn15  l=0.13u w=0.46u m=1
M10 GND E N_9 GND mn15  l=0.13u w=0.46u m=1
M11 Y F N_9 GND mn15  l=0.13u w=0.46u m=1
M12 Y F N_14 GND mn15  l=0.13u w=0.46u m=1
M13 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD B N_26 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD B N_26 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD A N_26 VDD mp15  l=0.13u w=0.69u m=1
M17 N_26 C N_22 VDD mp15  l=0.13u w=0.69u m=1
M18 N_26 D N_22 VDD mp15  l=0.13u w=0.69u m=1
M19 N_22 D N_26 VDD mp15  l=0.13u w=0.69u m=1
M20 N_22 C N_26 VDD mp15  l=0.13u w=0.69u m=1
M21 Y E N_22 VDD mp15  l=0.13u w=0.69u m=1
M22 N_22 E Y VDD mp15  l=0.13u w=0.69u m=1
M23 N_22 F Y VDD mp15  l=0.13u w=0.69u m=1
M24 N_22 F Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi222d2
* SPICE INPUT		Tue Jul 31 18:40:08 2018	aoi222d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi222d4
.subckt aoi222d4 GND Y A D C B VDD F E
M1 GND E N_15 GND mn15  l=0.13u w=0.46u m=1
M2 Y F N_15 GND mn15  l=0.13u w=0.46u m=1
M3 Y F N_26 GND mn15  l=0.13u w=0.46u m=1
M4 N_26 E GND GND mn15  l=0.13u w=0.46u m=1
M5 N_25 E GND GND mn15  l=0.13u w=0.46u m=1
M6 N_25 F Y GND mn15  l=0.13u w=0.46u m=1
M7 Y F N_24 GND mn15  l=0.13u w=0.46u m=1
M8 N_24 E GND GND mn15  l=0.13u w=0.46u m=1
M9 N_23 C GND GND mn15  l=0.13u w=0.46u m=1
M10 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M11 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M12 Y D N_22 GND mn15  l=0.13u w=0.46u m=1
M13 N_22 C GND GND mn15  l=0.13u w=0.46u m=1
M14 N_21 C GND GND mn15  l=0.13u w=0.46u m=1
M15 N_21 D Y GND mn15  l=0.13u w=0.46u m=1
M16 Y D N_20 GND mn15  l=0.13u w=0.46u m=1
M17 N_20 C GND GND mn15  l=0.13u w=0.46u m=1
M18 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M19 N_19 B Y GND mn15  l=0.13u w=0.46u m=1
M20 Y B N_18 GND mn15  l=0.13u w=0.46u m=1
M21 N_18 A GND GND mn15  l=0.13u w=0.46u m=1
M22 N_17 A GND GND mn15  l=0.13u w=0.46u m=1
M23 N_17 B Y GND mn15  l=0.13u w=0.46u m=1
M24 Y B N_16 GND mn15  l=0.13u w=0.46u m=1
M25 N_47 E Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_47 F Y VDD mp15  l=0.13u w=0.69u m=1
M27 N_47 F Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y E N_47 VDD mp15  l=0.13u w=0.69u m=1
M29 N_47 E Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y F N_47 VDD mp15  l=0.13u w=0.69u m=1
M31 N_47 F Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y E N_47 VDD mp15  l=0.13u w=0.69u m=1
M33 N_47 C N_41 VDD mp15  l=0.13u w=0.69u m=1
M34 N_41 D N_47 VDD mp15  l=0.13u w=0.69u m=1
M35 N_47 D N_41 VDD mp15  l=0.13u w=0.69u m=1
M36 N_41 C N_47 VDD mp15  l=0.13u w=0.69u m=1
M37 N_47 C N_41 VDD mp15  l=0.13u w=0.69u m=1
M38 N_41 D N_47 VDD mp15  l=0.13u w=0.69u m=1
M39 N_47 D N_41 VDD mp15  l=0.13u w=0.69u m=1
M40 N_41 C N_47 VDD mp15  l=0.13u w=0.69u m=1
M41 N_41 A VDD VDD mp15  l=0.13u w=0.69u m=1
M42 VDD A N_41 VDD mp15  l=0.13u w=0.69u m=1
M43 VDD B N_41 VDD mp15  l=0.13u w=0.69u m=1
M44 VDD B N_41 VDD mp15  l=0.13u w=0.69u m=1
M45 N_41 A VDD VDD mp15  l=0.13u w=0.69u m=1
M46 VDD A N_41 VDD mp15  l=0.13u w=0.69u m=1
M47 N_41 B VDD VDD mp15  l=0.13u w=0.69u m=1
M48 VDD B N_41 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi222d4
* SPICE INPUT		Tue Jul 31 18:40:20 2018	aoi22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d0
.subckt aoi22d0 GND Y VDD C D B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y D N_5 GND mn15  l=0.13u w=0.26u m=1
M4 GND C N_5 GND mn15  l=0.13u w=0.26u m=1
M5 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_10 B VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_10 D Y VDD mp15  l=0.13u w=0.4u m=1
M8 Y C N_10 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi22d0
* SPICE INPUT		Tue Jul 31 18:40:33 2018	aoi22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d1
.subckt aoi22d1 GND Y VDD C D B A
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 Y D N_5 GND mn15  l=0.13u w=0.46u m=1
M4 GND C N_5 GND mn15  l=0.13u w=0.46u m=1
M5 VDD A N_10 VDD mp15  l=0.13u w=0.69u m=1
M6 N_10 B VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_10 D Y VDD mp15  l=0.13u w=0.69u m=1
M8 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi22d1
* SPICE INPUT		Tue Jul 31 18:40:46 2018	aoi22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d2
.subckt aoi22d2 GND Y VDD D C A B
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_9 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_8 GND mn15  l=0.13u w=0.46u m=1
M4 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_10 C GND GND mn15  l=0.13u w=0.46u m=1
M6 Y D N_7 GND mn15  l=0.13u w=0.46u m=1
M7 Y D N_10 GND mn15  l=0.13u w=0.46u m=1
M8 N_7 C GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M10 VDD B N_16 VDD mp15  l=0.13u w=0.69u m=1
M11 N_16 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y C N_16 VDD mp15  l=0.13u w=0.69u m=1
M14 N_16 D Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_16 D Y VDD mp15  l=0.13u w=0.69u m=1
M16 N_16 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi22d2
* SPICE INPUT		Tue Jul 31 18:40:59 2018	aoi22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d4
.subckt aoi22d4 GND Y VDD D C A B
M1 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_12 GND mn15  l=0.13u w=0.46u m=1
M4 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_15 B Y GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_14 GND mn15  l=0.13u w=0.46u m=1
M8 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M10 N_17 D Y GND mn15  l=0.13u w=0.46u m=1
M11 Y D N_16 GND mn15  l=0.13u w=0.46u m=1
M12 N_18 C GND GND mn15  l=0.13u w=0.46u m=1
M13 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M14 Y D N_11 GND mn15  l=0.13u w=0.46u m=1
M15 Y D N_18 GND mn15  l=0.13u w=0.46u m=1
M16 N_11 C GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD A N_28 VDD mp15  l=0.13u w=0.69u m=1
M18 VDD B N_28 VDD mp15  l=0.13u w=0.69u m=1
M19 N_28 B VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_28 VDD mp15  l=0.13u w=0.69u m=1
M21 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD B N_28 VDD mp15  l=0.13u w=0.69u m=1
M23 N_28 B VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 Y C N_28 VDD mp15  l=0.13u w=0.69u m=1
M26 Y D N_28 VDD mp15  l=0.13u w=0.69u m=1
M27 N_28 D Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y C N_28 VDD mp15  l=0.13u w=0.69u m=1
M29 N_28 C Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_28 D Y VDD mp15  l=0.13u w=0.69u m=1
M31 N_28 D Y VDD mp15  l=0.13u w=0.69u m=1
M32 N_28 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi22d4
* SPICE INPUT		Tue Jul 31 18:41:11 2018	aoi22dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22dm
.subckt aoi22dm GND Y VDD C D B A
M1 N_6 A GND GND mn15  l=0.13u w=0.36u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.36u m=1
M3 Y D N_5 GND mn15  l=0.13u w=0.36u m=1
M4 GND C N_5 GND mn15  l=0.13u w=0.36u m=1
M5 N_10 A VDD VDD mp15  l=0.13u w=0.55u m=1
M6 N_10 B VDD VDD mp15  l=0.13u w=0.55u m=1
M7 N_10 D Y VDD mp15  l=0.13u w=0.55u m=1
M8 N_10 C Y VDD mp15  l=0.13u w=0.55u m=1
.ends aoi22dm
* SPICE INPUT		Tue Jul 31 18:41:24 2018	aoi2m1d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi2m1d0
.subckt aoi2m1d0 Y GND VDD C A BN
M1 N_5 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 N_5 Y GND mn15  l=0.13u w=0.26u m=1
M4 GND C Y GND mn15  l=0.13u w=0.26u m=1
M5 VDD BN N_5 VDD mp15  l=0.13u w=0.4u m=1
M6 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 VDD N_5 N_10 VDD mp15  l=0.13u w=0.4u m=1
M8 Y C N_10 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi2m1d0
* SPICE INPUT		Tue Jul 31 18:41:39 2018	aoi2m1d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi2m1d1
.subckt aoi2m1d1 GND Y VDD C A BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_7 N_3 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND C Y GND mn15  l=0.13u w=0.26u m=1
M5 N_3 BN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 VDD A N_11 VDD mp15  l=0.13u w=0.69u m=1
M7 VDD N_3 N_11 VDD mp15  l=0.13u w=0.69u m=1
M8 Y C N_11 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi2m1d1
* SPICE INPUT		Tue Jul 31 18:41:58 2018	aoi2m1d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi2m1d2
.subckt aoi2m1d2 GND Y VDD C A BN
M1 GND BN N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_8 N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_4 N_7 GND mn15  l=0.13u w=0.46u m=1
M5 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M6 Y C GND GND mn15  l=0.13u w=0.46u m=1
M7 VDD BN N_4 VDD mp15  l=0.13u w=0.69u m=1
M8 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_4 N_13 VDD mp15  l=0.13u w=0.69u m=1
M10 N_13 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
M13 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi2m1d2
* SPICE INPUT		Tue Jul 31 18:42:12 2018	aoi2m1d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi2m1d4
.subckt aoi2m1d4 Y GND VDD C A BN
M1 N_6 BN GND GND mn15  l=0.13u w=0.46u m=1
M2 N_6 BN GND GND mn15  l=0.13u w=0.46u m=1
M3 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_12 N_6 Y GND mn15  l=0.13u w=0.46u m=1
M5 Y N_6 N_11 GND mn15  l=0.13u w=0.46u m=1
M6 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_14 N_6 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_6 N_13 GND mn15  l=0.13u w=0.46u m=1
M10 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M11 GND C Y GND mn15  l=0.13u w=0.46u m=1
M12 GND C Y GND mn15  l=0.13u w=0.46u m=1
M13 VDD BN N_6 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD BN N_6 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_6 N_20 VDD mp15  l=0.13u w=0.69u m=1
M17 N_20 N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M19 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_6 N_20 VDD mp15  l=0.13u w=0.69u m=1
M21 N_20 N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_20 C Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y C N_20 VDD mp15  l=0.13u w=0.69u m=1
M25 N_20 C Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_20 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi2m1d4
* SPICE INPUT		Tue Jul 31 18:42:24 2018	aoi31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d0
.subckt aoi31d0 GND Y VDD D C B A
M1 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y D GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 C Y GND mn15  l=0.13u w=0.26u m=1
M5 N_11 A VDD VDD mp15  l=0.13u w=0.35u m=1
M6 Y D N_11 VDD mp15  l=0.13u w=0.4u m=1
M7 VDD B N_11 VDD mp15  l=0.13u w=0.38u m=1
M8 VDD C N_11 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi31d0
* SPICE INPUT		Tue Jul 31 18:42:36 2018	aoi31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d1
.subckt aoi31d1 GND Y VDD D C B A
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_6 B N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M4 Y D GND GND mn15  l=0.13u w=0.26u m=1
M5 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 VDD B N_11 VDD mp15  l=0.13u w=0.69u m=1
M7 VDD C N_11 VDD mp15  l=0.13u w=0.69u m=1
M8 Y D N_11 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi31d1
* SPICE INPUT		Tue Jul 31 18:42:48 2018	aoi31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d2
.subckt aoi31d2 GND Y C B A D VDD
M1 Y D GND GND mn15  l=0.13u w=0.46u m=1
M2 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_9 B N_8 GND mn15  l=0.13u w=0.46u m=1
M4 Y C N_7 GND mn15  l=0.13u w=0.46u m=1
M5 N_8 C Y GND mn15  l=0.13u w=0.46u m=1
M6 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M7 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_18 D Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_18 D Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_18 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_18 C VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_18 C VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_18 B VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi31d2
* SPICE INPUT		Tue Jul 31 18:43:00 2018	aoi31d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d4
.subckt aoi31d4 GND Y VDD D C B A
M1 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_2 B N_3 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M9 Y C N_3 GND mn15  l=0.13u w=0.46u m=1
M10 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M11 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M12 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M13 Y D GND GND mn15  l=0.13u w=0.46u m=1
M14 Y D GND GND mn15  l=0.13u w=0.46u m=1
M15 N_19 A VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_19 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_19 VDD mp15  l=0.13u w=0.69u m=1
M18 N_19 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_19 B VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_19 B VDD VDD mp15  l=0.13u w=0.61u m=1
M21 N_19 B VDD VDD mp15  l=0.13u w=0.61u m=1
M22 VDD B N_19 VDD mp15  l=0.13u w=0.61u m=1
M23 VDD C N_19 VDD mp15  l=0.13u w=0.575u m=1
M24 VDD C N_19 VDD mp15  l=0.13u w=0.575u m=1
M25 N_19 C VDD VDD mp15  l=0.13u w=0.575u m=1
M26 VDD C N_19 VDD mp15  l=0.13u w=0.575u m=1
M27 N_19 C VDD VDD mp15  l=0.13u w=0.575u m=1
M28 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M29 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M31 Y D N_19 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi31d4
* SPICE INPUT		Tue Jul 31 18:43:11 2018	aoi31dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31dm
.subckt aoi31dm GND Y VDD D C B A
M1 N_5 A GND GND mn15  l=0.13u w=0.36u m=1
M2 N_6 B N_5 GND mn15  l=0.13u w=0.36u m=1
M3 N_6 C Y GND mn15  l=0.13u w=0.36u m=1
M4 Y D GND GND mn15  l=0.13u w=0.26u m=1
M5 N_11 A VDD VDD mp15  l=0.13u w=0.55u m=1
M6 VDD B N_11 VDD mp15  l=0.13u w=0.55u m=1
M7 VDD C N_11 VDD mp15  l=0.13u w=0.55u m=1
M8 Y D N_11 VDD mp15  l=0.13u w=0.55u m=1
.ends aoi31dm
* SPICE INPUT		Tue Jul 31 18:43:23 2018	aoi32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d0
.subckt aoi32d0 GND Y VDD D E C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y C N_7 GND mn15  l=0.13u w=0.26u m=1
M4 Y E N_5 GND mn15  l=0.13u w=0.26u m=1
M5 GND D N_5 GND mn15  l=0.13u w=0.26u m=1
M6 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_13 B VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_13 C VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_13 E Y VDD mp15  l=0.13u w=0.4u m=1
M10 N_13 D Y VDD mp15  l=0.13u w=0.4u m=1
.ends aoi32d0
* SPICE INPUT		Tue Jul 31 18:43:36 2018	aoi32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d1
.subckt aoi32d1 GND Y VDD D E C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_7 C Y GND mn15  l=0.13u w=0.46u m=1
M4 Y E N_5 GND mn15  l=0.13u w=0.36u m=1
M5 GND D N_5 GND mn15  l=0.13u w=0.36u m=1
M6 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 VDD B N_13 VDD mp15  l=0.13u w=0.69u m=1
M8 N_13 C VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_13 E Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_13 D Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi32d1
* SPICE INPUT		Tue Jul 31 18:43:47 2018	aoi32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d2
.subckt aoi32d2 GND Y VDD D E A B C
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_9 B N_8 GND mn15  l=0.13u w=0.46u m=1
M3 GND D N_7 GND mn15  l=0.13u w=0.36u m=1
M4 Y E N_7 GND mn15  l=0.13u w=0.36u m=1
M5 Y E N_12 GND mn15  l=0.13u w=0.36u m=1
M6 N_12 D GND GND mn15  l=0.13u w=0.36u m=1
M7 N_10 C Y GND mn15  l=0.13u w=0.46u m=1
M8 Y C N_9 GND mn15  l=0.13u w=0.46u m=1
M9 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M10 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M11 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_21 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_21 D Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_21 E Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_21 E Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y D N_21 VDD mp15  l=0.13u w=0.69u m=1
M17 N_21 C VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_21 C VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD B N_21 VDD mp15  l=0.13u w=0.69u m=1
M20 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi32d2
* SPICE INPUT		Tue Jul 31 18:43:59 2018	aoi32d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d4
.subckt aoi32d4 GND Y D E C VDD B A
M1 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_2 B N_3 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 D GND GND mn15  l=0.13u w=0.36u m=1
M10 N_12 D GND GND mn15  l=0.13u w=0.36u m=1
M11 N_12 D GND GND mn15  l=0.13u w=0.36u m=1
M12 GND D N_12 GND mn15  l=0.13u w=0.36u m=1
M13 Y C N_3 GND mn15  l=0.13u w=0.46u m=1
M14 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M15 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M16 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M17 N_12 E Y GND mn15  l=0.13u w=0.48u m=1
M18 N_12 E Y GND mn15  l=0.13u w=0.48u m=1
M19 N_12 E Y GND mn15  l=0.13u w=0.48u m=1
M20 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD A N_24 VDD mp15  l=0.13u w=0.69u m=1
M23 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_24 B VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_24 B VDD VDD mp15  l=0.13u w=0.61u m=1
M26 N_24 B VDD VDD mp15  l=0.13u w=0.61u m=1
M27 VDD B N_24 VDD mp15  l=0.13u w=0.61u m=1
M28 N_24 D Y VDD mp15  l=0.13u w=0.69u m=1
M29 N_24 D Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_24 D Y VDD mp15  l=0.13u w=0.69u m=1
M31 Y D N_24 VDD mp15  l=0.13u w=0.69u m=1
M32 N_24 C VDD VDD mp15  l=0.13u w=0.575u m=1
M33 VDD C N_24 VDD mp15  l=0.13u w=0.575u m=1
M34 N_24 C VDD VDD mp15  l=0.13u w=0.575u m=1
M35 VDD C N_24 VDD mp15  l=0.13u w=0.575u m=1
M36 N_24 C VDD VDD mp15  l=0.13u w=0.575u m=1
M37 N_24 E Y VDD mp15  l=0.13u w=0.605u m=1
M38 Y E N_24 VDD mp15  l=0.13u w=0.605u m=1
M39 N_24 E Y VDD mp15  l=0.13u w=0.605u m=1
M40 N_24 E Y VDD mp15  l=0.13u w=0.645u m=1
.ends aoi32d4
* SPICE INPUT		Tue Jul 31 18:44:11 2018	aoi32dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32dm
.subckt aoi32dm GND Y VDD D E C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.36u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.36u m=1
M3 N_7 C Y GND mn15  l=0.13u w=0.36u m=1
M4 Y E N_5 GND mn15  l=0.13u w=0.3u m=1
M5 GND D N_5 GND mn15  l=0.13u w=0.3u m=1
M6 N_13 A VDD VDD mp15  l=0.13u w=0.55u m=1
M7 N_13 B VDD VDD mp15  l=0.13u w=0.55u m=1
M8 N_13 C VDD VDD mp15  l=0.13u w=0.55u m=1
M9 N_13 E Y VDD mp15  l=0.13u w=0.55u m=1
M10 N_13 D Y VDD mp15  l=0.13u w=0.55u m=1
.ends aoi32dm
* SPICE INPUT		Tue Jul 31 18:44:23 2018	aoi33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d0
.subckt aoi33d0 GND Y VDD D E F C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y C N_7 GND mn15  l=0.13u w=0.26u m=1
M4 N_8 F Y GND mn15  l=0.13u w=0.26u m=1
M5 N_8 E N_5 GND mn15  l=0.13u w=0.26u m=1
M6 GND D N_5 GND mn15  l=0.13u w=0.26u m=1
M7 N_15 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_15 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_15 C VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y F N_15 VDD mp15  l=0.13u w=0.4u m=1
M11 Y E N_15 VDD mp15  l=0.13u w=0.4u m=1
M12 Y D N_15 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi33d0
* SPICE INPUT		Tue Jul 31 18:44:36 2018	aoi33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d1
.subckt aoi33d1 GND Y VDD D E F C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 Y C N_7 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 F Y GND mn15  l=0.13u w=0.46u m=1
M5 N_8 E N_5 GND mn15  l=0.13u w=0.46u m=1
M6 GND D N_5 GND mn15  l=0.13u w=0.46u m=1
M7 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_15 B VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_15 C VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y F N_15 VDD mp15  l=0.13u w=0.69u m=1
M11 Y E N_15 VDD mp15  l=0.13u w=0.69u m=1
M12 Y D N_15 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi33d1
* SPICE INPUT		Tue Jul 31 18:44:51 2018	aoi33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d2
.subckt aoi33d2 Y GND A C D E VDD B F
M1 Y F N_10 GND mn15  l=0.13u w=0.46u m=1
M2 N_11 F Y GND mn15  l=0.13u w=0.46u m=1
M3 N_11 E N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 E N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_2 D GND GND mn15  l=0.13u w=0.46u m=1
M7 GND D N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_13 B N_12 GND mn15  l=0.13u w=0.46u m=1
M9 GND A N_15 GND mn15  l=0.13u w=0.46u m=1
M10 N_15 B N_14 GND mn15  l=0.13u w=0.46u m=1
M11 Y C N_13 GND mn15  l=0.13u w=0.46u m=1
M12 N_14 C Y GND mn15  l=0.13u w=0.46u m=1
M13 Y F N_28 VDD mp15  l=0.13u w=0.565u m=1
M14 Y F N_28 VDD mp15  l=0.13u w=0.405u m=1
M15 N_28 F Y VDD mp15  l=0.13u w=0.41u m=1
M16 VDD A N_28 VDD mp15  l=0.13u w=0.69u m=1
M17 N_28 E Y VDD mp15  l=0.13u w=0.69u m=1
M18 N_28 D Y VDD mp15  l=0.13u w=0.69u m=1
M19 Y D N_28 VDD mp15  l=0.13u w=0.69u m=1
M20 N_28 B VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 Y E N_28 VDD mp15  l=0.13u w=0.69u m=1
M23 VDD B N_28 VDD mp15  l=0.13u w=0.69u m=1
M24 N_28 C VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_28 C VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi33d2
* SPICE INPUT		Tue Jul 31 18:45:05 2018	aoi33d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d4
.subckt aoi33d4 GND Y VDD A B C F E D
M1 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 B N_3 GND mn15  l=0.13u w=0.46u m=1
M5 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_12 F Y GND mn15  l=0.13u w=0.46u m=1
M10 Y F N_12 GND mn15  l=0.13u w=0.46u m=1
M11 N_12 F Y GND mn15  l=0.13u w=0.46u m=1
M12 N_12 F Y GND mn15  l=0.13u w=0.46u m=1
M13 Y C N_3 GND mn15  l=0.13u w=0.46u m=1
M14 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M15 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M16 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M17 N_21 D GND GND mn15  l=0.13u w=0.46u m=1
M18 N_21 D GND GND mn15  l=0.13u w=0.46u m=1
M19 N_21 D GND GND mn15  l=0.13u w=0.46u m=1
M20 N_21 D GND GND mn15  l=0.13u w=0.46u m=1
M21 N_21 E N_12 GND mn15  l=0.13u w=0.46u m=1
M22 N_12 E N_21 GND mn15  l=0.13u w=0.46u m=1
M23 N_12 E N_21 GND mn15  l=0.13u w=0.46u m=1
M24 N_12 E N_21 GND mn15  l=0.13u w=0.46u m=1
M25 Y D N_35 VDD mp15  l=0.13u w=0.69u m=1
M26 N_35 D Y VDD mp15  l=0.13u w=0.69u m=1
M27 N_35 D Y VDD mp15  l=0.13u w=0.69u m=1
M28 N_35 D Y VDD mp15  l=0.13u w=0.69u m=1
M29 N_35 E Y VDD mp15  l=0.13u w=0.575u m=1
M30 N_35 E Y VDD mp15  l=0.13u w=0.55u m=1
M31 Y E N_35 VDD mp15  l=0.13u w=0.545u m=1
M32 N_35 E Y VDD mp15  l=0.13u w=0.545u m=1
M33 Y E N_35 VDD mp15  l=0.13u w=0.545u m=1
M34 N_35 F Y VDD mp15  l=0.13u w=0.56u m=1
M35 N_35 F Y VDD mp15  l=0.13u w=0.565u m=1
M36 N_35 F Y VDD mp15  l=0.13u w=0.545u m=1
M37 Y F N_35 VDD mp15  l=0.13u w=0.545u m=1
M38 N_35 F Y VDD mp15  l=0.13u w=0.545u m=1
M39 N_35 C VDD VDD mp15  l=0.13u w=0.545u m=1
M40 N_35 C VDD VDD mp15  l=0.13u w=0.555u m=1
M41 N_35 C VDD VDD mp15  l=0.13u w=0.555u m=1
M42 VDD C N_35 VDD mp15  l=0.13u w=0.555u m=1
M43 N_35 C VDD VDD mp15  l=0.13u w=0.555u m=1
M44 N_35 B VDD VDD mp15  l=0.13u w=0.6u m=1
M45 N_35 B VDD VDD mp15  l=0.13u w=0.6u m=1
M46 VDD B N_35 VDD mp15  l=0.13u w=0.6u m=1
M47 N_35 B VDD VDD mp15  l=0.13u w=0.69u m=1
M48 N_35 B VDD VDD mp15  l=0.13u w=0.265u m=1
M49 N_35 A VDD VDD mp15  l=0.13u w=0.69u m=1
M50 VDD A N_35 VDD mp15  l=0.13u w=0.69u m=1
M51 VDD A N_35 VDD mp15  l=0.13u w=0.69u m=1
M52 N_35 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi33d4
* SPICE INPUT		Tue Jul 31 18:45:20 2018	aoim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d0
.subckt aoim21d0 Y VDD AN C GND BN
M1 GND BN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 GND N_3 Y GND mn15  l=0.13u w=0.26u m=1
M3 GND C Y GND mn15  l=0.13u w=0.26u m=1
M4 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M5 N_8 BN N_3 VDD mp15  l=0.13u w=0.4u m=1
M6 VDD N_3 N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 Y C N_7 VDD mp15  l=0.13u w=0.4u m=1
M8 VDD AN N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends aoim21d0
* SPICE INPUT		Tue Jul 31 18:45:34 2018	aoim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d1
.subckt aoim21d1 Y VDD GND C AN BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_3 Y GND mn15  l=0.13u w=0.35u m=1
M4 GND C Y GND mn15  l=0.13u w=0.35u m=1
M5 N_6 BN N_3 VDD mp15  l=0.13u w=0.52u m=1
M6 VDD AN N_6 VDD mp15  l=0.13u w=0.52u m=1
M7 VDD N_3 N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 Y C N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends aoim21d1
* SPICE INPUT		Tue Jul 31 18:45:47 2018	aoim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d2
.subckt aoim21d2 VDD Y GND C AN BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.36u m=1
M2 GND AN N_3 GND mn15  l=0.13u w=0.36u m=1
M3 Y N_3 GND GND mn15  l=0.13u w=0.36u m=1
M4 GND C Y GND mn15  l=0.13u w=0.36u m=1
M5 GND C Y GND mn15  l=0.13u w=0.36u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.36u m=1
M7 N_7 BN N_3 VDD mp15  l=0.13u w=0.69u m=1
M8 VDD AN N_7 VDD mp15  l=0.13u w=0.69u m=1
M9 N_8 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y C N_6 VDD mp15  l=0.13u w=0.69u m=1
M11 Y C N_8 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_3 N_6 VDD mp15  l=0.13u w=0.69u m=1
.ends aoim21d2
* SPICE INPUT		Tue Jul 31 18:45:59 2018	aoim21d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d3
.subckt aoim21d3 VDD Y GND C AN BN
M1 N_4 AN GND GND mn15  l=0.13u w=0.35u m=1
M2 N_4 BN GND GND mn15  l=0.13u w=0.35u m=1
M3 N_4 BN GND GND mn15  l=0.13u w=0.33u m=1
M4 GND AN N_4 GND mn15  l=0.13u w=0.33u m=1
M5 Y C GND GND mn15  l=0.13u w=0.46u m=1
M6 Y C GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND C Y GND mn15  l=0.13u w=0.46u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M11 N_10 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_11 BN N_4 VDD mp15  l=0.13u w=0.69u m=1
M13 N_4 BN N_10 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD AN N_11 VDD mp15  l=0.13u w=0.69u m=1
M15 N_12 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
M17 N_13 C Y VDD mp15  l=0.13u w=0.62u m=1
M18 N_14 N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
M19 VDD N_4 N_13 VDD mp15  l=0.13u w=0.62u m=1
M20 Y C N_9 VDD mp15  l=0.13u w=0.685u m=1
M21 N_14 C Y VDD mp15  l=0.13u w=0.695u m=1
M22 N_9 N_4 VDD VDD mp15  l=0.13u w=0.685u m=1
.ends aoim21d3
* SPICE INPUT		Tue Jul 31 18:46:11 2018	aoim21dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21dm
.subckt aoim21dm Y VDD GND C AN BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_3 Y GND mn15  l=0.13u w=0.28u m=1
M4 GND C Y GND mn15  l=0.13u w=0.28u m=1
M5 N_8 BN N_3 VDD mp15  l=0.13u w=0.4u m=1
M6 VDD AN N_8 VDD mp15  l=0.13u w=0.4u m=1
M7 VDD N_3 N_7 VDD mp15  l=0.13u w=0.55u m=1
M8 Y C N_7 VDD mp15  l=0.13u w=0.55u m=1
.ends aoim21dm
* SPICE INPUT		Tue Jul 31 18:46:24 2018	aoim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d0
.subckt aoim22d0 GND Y VDD C D BN AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 BN GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M4 Y D N_7 GND mn15  l=0.13u w=0.26u m=1
M5 GND C N_7 GND mn15  l=0.13u w=0.26u m=1
M6 VDD AN N_32 VDD mp15  l=0.13u w=0.4u m=1
M7 N_5 BN N_32 VDD mp15  l=0.13u w=0.4u m=1
M8 N_11 N_5 Y VDD mp15  l=0.13u w=0.4u m=1
M9 N_11 D VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_11 C VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aoim22d0
* SPICE INPUT		Tue Jul 31 18:46:36 2018	aoim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d1
.subckt aoim22d1 GND Y C D VDD BN AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 BN GND GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_7 GND mn15  l=0.13u w=0.46u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M5 Y D N_7 GND mn15  l=0.13u w=0.46u m=1
M6 VDD AN N_32 VDD mp15  l=0.13u w=0.52u m=1
M7 N_32 BN N_5 VDD mp15  l=0.13u w=0.52u m=1
M8 N_11 C VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_11 N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_11 D VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoim22d1
* SPICE INPUT		Tue Jul 31 18:46:50 2018	aoim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d2
.subckt aoim22d2 GND Y VDD C D BN AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.36u m=1
M2 N_5 BN GND GND mn15  l=0.13u w=0.36u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M4 GND C N_9 GND mn15  l=0.13u w=0.47u m=1
M5 N_10 C GND GND mn15  l=0.13u w=0.45u m=1
M6 Y D N_9 GND mn15  l=0.13u w=0.47u m=1
M7 Y D N_10 GND mn15  l=0.13u w=0.45u m=1
M8 VDD AN N_20 VDD mp15  l=0.13u w=0.69u m=1
M9 N_20 BN N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 N_14 C VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_14 N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
M13 N_14 C VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_14 D VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_14 D VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoim22d2
* SPICE INPUT		Tue Jul 31 18:47:10 2018	aoim22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d4
.subckt aoim22d4 GND Y VDD AN BN C D
M1 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M2 N_15 D Y GND mn15  l=0.13u w=0.46u m=1
M3 Y D N_14 GND mn15  l=0.13u w=0.46u m=1
M4 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_15 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_17 D Y GND mn15  l=0.13u w=0.46u m=1
M7 Y D N_16 GND mn15  l=0.13u w=0.46u m=1
M8 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M10 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_3 AN GND GND mn15  l=0.13u w=0.35u m=1
M12 GND AN N_3 GND mn15  l=0.13u w=0.35u m=1
M13 N_3 BN GND GND mn15  l=0.13u w=0.35u m=1
M14 GND BN N_3 GND mn15  l=0.13u w=0.35u m=1
M15 VDD C N_25 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD D N_25 VDD mp15  l=0.13u w=0.69u m=1
M17 N_25 D VDD VDD mp15  l=0.13u w=0.69u m=1
M18 VDD C N_25 VDD mp15  l=0.13u w=0.69u m=1
M19 N_25 C VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD D N_25 VDD mp15  l=0.13u w=0.69u m=1
M21 N_25 D VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_25 C VDD VDD mp15  l=0.13u w=0.69u m=1
M23 Y N_3 N_25 VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_3 N_25 VDD mp15  l=0.13u w=0.69u m=1
M25 N_25 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_25 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M27 N_31 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M28 N_3 BN N_30 VDD mp15  l=0.13u w=0.69u m=1
M29 N_3 BN N_31 VDD mp15  l=0.13u w=0.69u m=1
M30 N_30 AN VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoim22d4
* SPICE INPUT		Tue Jul 31 18:47:24 2018	aoim22dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22dm
.subckt aoim22dm GND Y C D VDD BN AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 BN GND GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_7 GND mn15  l=0.13u w=0.36u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M5 Y D N_7 GND mn15  l=0.13u w=0.36u m=1
M6 VDD AN N_32 VDD mp15  l=0.13u w=0.34u m=1
M7 N_32 BN N_5 VDD mp15  l=0.13u w=0.34u m=1
M8 N_11 C VDD VDD mp15  l=0.13u w=0.55u m=1
M9 N_11 N_5 Y VDD mp15  l=0.13u w=0.55u m=1
M10 N_11 D VDD VDD mp15  l=0.13u w=0.55u m=1
.ends aoim22dm
* SPICE INPUT		Tue Jul 31 18:47:36 2018	aor211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d0
.subckt aor211d0 Y GND VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 C GND GND mn15  l=0.13u w=0.26u m=1
M3 N_7 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.26u m=1
M6 N_16 D N_5 VDD mp15  l=0.13u w=0.38u m=1
M7 N_16 C N_11 VDD mp15  l=0.13u w=0.38u m=1
M8 N_11 B VDD VDD mp15  l=0.13u w=0.38u m=1
M9 N_11 A VDD VDD mp15  l=0.13u w=0.38u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor211d0
* SPICE INPUT		Tue Jul 31 18:47:47 2018	aor211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d1
.subckt aor211d1 GND Y VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 C GND GND mn15  l=0.13u w=0.26u m=1
M3 N_7 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_16 D N_5 VDD mp15  l=0.13u w=0.38u m=1
M7 N_16 C N_11 VDD mp15  l=0.13u w=0.38u m=1
M8 N_11 B VDD VDD mp15  l=0.13u w=0.38u m=1
M9 N_11 A VDD VDD mp15  l=0.13u w=0.38u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor211d1
* SPICE INPUT		Tue Jul 31 18:47:59 2018	aor211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d2
.subckt aor211d2 Y GND A B C D VDD
M1 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_6 D GND GND mn15  l=0.13u w=0.26u m=1
M4 N_6 C GND GND mn15  l=0.13u w=0.26u m=1
M5 N_9 B N_6 GND mn15  l=0.13u w=0.46u m=1
M6 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M7 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_6 D N_37 VDD mp15  l=0.13u w=0.69u m=1
M10 N_13 C N_37 VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
.ends aor211d2
* SPICE INPUT		Tue Jul 31 18:48:13 2018	aor211d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d4
.subckt aor211d4 GND Y VDD C D A B
M1 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 B N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B N_12 GND mn15  l=0.13u w=0.46u m=1
M4 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND C N_3 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 D GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M10 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M11 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_17 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_17 B VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_25 C N_17 VDD mp15  l=0.13u w=0.69u m=1
M16 N_3 D N_24 VDD mp15  l=0.13u w=0.69u m=1
M17 N_3 D N_25 VDD mp15  l=0.13u w=0.69u m=1
M18 N_17 C N_24 VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor211d4
* SPICE INPUT		Tue Jul 31 18:48:25 2018	aor21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d0
.subckt aor21d0 GND Y VDD C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_10 A VDD VDD mp15  l=0.13u w=0.38u m=1
M6 VDD B N_10 VDD mp15  l=0.13u w=0.38u m=1
M7 N_5 C N_10 VDD mp15  l=0.13u w=0.38u m=1
M8 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor21d0
* SPICE INPUT		Tue Jul 31 18:48:36 2018	aor21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d1
.subckt aor21d1 GND Y VDD C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_10 A VDD VDD mp15  l=0.13u w=0.38u m=1
M6 VDD B N_10 VDD mp15  l=0.13u w=0.38u m=1
M7 N_5 C N_10 VDD mp15  l=0.13u w=0.38u m=1
M8 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor21d1
* SPICE INPUT		Tue Jul 31 18:48:48 2018	aor21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d2
.subckt aor21d2 GND Y VDD C B A
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_8 B N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 C GND GND mn15  l=0.13u w=0.26u m=1
M4 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M6 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M7 VDD B N_12 VDD mp15  l=0.13u w=0.69u m=1
M8 N_3 C N_12 VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor21d2
* SPICE INPUT		Tue Jul 31 18:49:02 2018	aor21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d4
.subckt aor21d4 GND Y VDD C A B
M1 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 B N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B N_11 GND mn15  l=0.13u w=0.46u m=1
M4 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M7 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M8 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M10 VDD A N_17 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD B N_17 VDD mp15  l=0.13u w=0.69u m=1
M12 N_17 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_17 C N_3 VDD mp15  l=0.13u w=0.69u m=1
M15 N_17 C N_3 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M19 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor21d4
* SPICE INPUT		Tue Jul 31 18:49:17 2018	aor221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d0
.subckt aor221d0 GND Y VDD E D C A B
M1 N_8 B N_3 GND mn15  l=0.13u w=0.26u m=1
M2 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_9 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_9 D N_3 GND mn15  l=0.13u w=0.26u m=1
M5 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_15 B VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_15 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_15 C N_14 VDD mp15  l=0.13u w=0.4u m=1
M10 N_14 D N_15 VDD mp15  l=0.13u w=0.4u m=1
M11 N_3 E N_14 VDD mp15  l=0.13u w=0.4u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor221d0
* SPICE INPUT		Tue Jul 31 18:49:31 2018	aor221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d1
.subckt aor221d1 GND Y VDD E D C A B
M1 N_8 B N_3 GND mn15  l=0.13u w=0.26u m=1
M2 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_9 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_9 D N_3 GND mn15  l=0.13u w=0.26u m=1
M5 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_15 B VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_15 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_15 C N_14 VDD mp15  l=0.13u w=0.4u m=1
M10 N_14 D N_15 VDD mp15  l=0.13u w=0.4u m=1
M11 N_3 E N_14 VDD mp15  l=0.13u w=0.4u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor221d1
* SPICE INPUT		Tue Jul 31 18:49:44 2018	aor221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d2
.subckt aor221d2 GND Y VDD E C D B A
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 B N_10 GND mn15  l=0.13u w=0.46u m=1
M3 N_4 D N_9 GND mn15  l=0.13u w=0.46u m=1
M4 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_4 E GND GND mn15  l=0.13u w=0.26u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M9 N_16 B VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_16 D N_15 VDD mp15  l=0.13u w=0.69u m=1
M11 N_15 C N_16 VDD mp15  l=0.13u w=0.69u m=1
M12 N_4 E N_15 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor221d2
* SPICE INPUT		Tue Jul 31 18:50:00 2018	aor221d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d4
.subckt aor221d4 Y GND D C B E A VDD
M1 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M2 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M5 N_8 E GND GND mn15  l=0.13u w=0.46u m=1
M6 N_16 D N_8 GND mn15  l=0.13u w=0.46u m=1
M7 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M8 N_15 C GND GND mn15  l=0.13u w=0.46u m=1
M9 N_15 D N_8 GND mn15  l=0.13u w=0.46u m=1
M10 N_8 B N_14 GND mn15  l=0.13u w=0.46u m=1
M11 N_13 B N_8 GND mn15  l=0.13u w=0.46u m=1
M12 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M13 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M14 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M17 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_8 E N_27 VDD mp15  l=0.13u w=0.69u m=1
M19 N_27 E N_8 VDD mp15  l=0.13u w=0.69u m=1
M20 N_27 D N_22 VDD mp15  l=0.13u w=0.69u m=1
M21 N_22 C N_27 VDD mp15  l=0.13u w=0.69u m=1
M22 N_22 C N_27 VDD mp15  l=0.13u w=0.69u m=1
M23 N_27 D N_22 VDD mp15  l=0.13u w=0.69u m=1
M24 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor221d4
* SPICE INPUT		Tue Jul 31 18:50:15 2018	aor222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor222d0
.subckt aor222d0 GND Y A D B VDD C E F
M1 N_9 F N_2 GND mn15  l=0.13u w=0.26u m=1
M2 N_9 E GND GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_8 GND mn15  l=0.13u w=0.26u m=1
M4 N_2 D N_8 GND mn15  l=0.13u w=0.26u m=1
M5 N_10 B N_2 GND mn15  l=0.13u w=0.26u m=1
M6 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_2 F N_19 VDD mp15  l=0.13u w=0.4u m=1
M9 N_19 E N_2 VDD mp15  l=0.13u w=0.4u m=1
M10 N_19 C N_15 VDD mp15  l=0.13u w=0.4u m=1
M11 N_15 D N_19 VDD mp15  l=0.13u w=0.4u m=1
M12 N_15 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_15 A VDD VDD mp15  l=0.13u w=0.4u m=1
M14 Y N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor222d0
* SPICE INPUT		Tue Jul 31 18:50:26 2018	aor222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor222d1
.subckt aor222d1 GND Y VDD B A D C E F
M1 N_9 F N_2 GND mn15  l=0.13u w=0.26u m=1
M2 N_9 E GND GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_8 GND mn15  l=0.13u w=0.26u m=1
M4 N_2 D N_8 GND mn15  l=0.13u w=0.26u m=1
M5 N_10 B N_2 GND mn15  l=0.13u w=0.26u m=1
M6 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_2 F N_19 VDD mp15  l=0.13u w=0.4u m=1
M9 N_19 E N_2 VDD mp15  l=0.13u w=0.4u m=1
M10 N_19 C N_17 VDD mp15  l=0.13u w=0.4u m=1
M11 N_17 D N_19 VDD mp15  l=0.13u w=0.4u m=1
M12 N_17 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_17 A VDD VDD mp15  l=0.13u w=0.4u m=1
M14 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor222d1
* SPICE INPUT		Tue Jul 31 18:50:37 2018	aor222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor222d2
.subckt aor222d2 GND Y VDD A B D C E F
M1 N_10 F N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_10 E GND GND mn15  l=0.13u w=0.46u m=1
M3 GND C N_9 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 D N_9 GND mn15  l=0.13u w=0.46u m=1
M5 N_11 B N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_2 F N_19 VDD mp15  l=0.13u w=0.69u m=1
M10 N_19 E N_2 VDD mp15  l=0.13u w=0.69u m=1
M11 N_19 C N_17 VDD mp15  l=0.13u w=0.69u m=1
M12 N_19 D N_17 VDD mp15  l=0.13u w=0.69u m=1
M13 N_17 B VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_17 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor222d2
* SPICE INPUT		Tue Jul 31 18:50:50 2018	aor222d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor222d4
.subckt aor222d4 Y GND VDD A B D C E F
M1 N_13 E GND GND mn15  l=0.13u w=0.46u m=1
M2 N_14 F N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_5 F N_13 GND mn15  l=0.13u w=0.46u m=1
M4 N_14 E GND GND mn15  l=0.13u w=0.46u m=1
M5 N_15 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_16 D N_5 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 D N_15 GND mn15  l=0.13u w=0.46u m=1
M8 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M9 N_17 A GND GND mn15  l=0.13u w=0.46u m=1
M10 N_18 B N_5 GND mn15  l=0.13u w=0.46u m=1
M11 N_5 B N_17 GND mn15  l=0.13u w=0.46u m=1
M12 N_18 A GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M15 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M16 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M17 N_5 E N_30 VDD mp15  l=0.13u w=0.69u m=1
M18 N_5 F N_30 VDD mp15  l=0.13u w=0.69u m=1
M19 N_30 F N_5 VDD mp15  l=0.13u w=0.69u m=1
M20 N_30 E N_5 VDD mp15  l=0.13u w=0.69u m=1
M21 N_27 C N_30 VDD mp15  l=0.13u w=0.69u m=1
M22 N_30 D N_27 VDD mp15  l=0.13u w=0.69u m=1
M23 N_30 D N_27 VDD mp15  l=0.13u w=0.69u m=1
M24 N_30 C N_27 VDD mp15  l=0.13u w=0.69u m=1
M25 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_27 B VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_27 B VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD A N_27 VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor222d4
* SPICE INPUT		Tue Jul 31 18:51:01 2018	aor22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d0
.subckt aor22d0 GND Y VDD A B D C
M1 GND C N_7 GND mn15  l=0.13u w=0.26u m=1
M2 N_2 D N_7 GND mn15  l=0.13u w=0.26u m=1
M3 N_8 B N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_2 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_13 C N_2 VDD mp15  l=0.13u w=0.4u m=1
M7 N_13 D N_2 VDD mp15  l=0.13u w=0.4u m=1
M8 N_13 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor22d0
* SPICE INPUT		Tue Jul 31 18:51:13 2018	aor22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d1
.subckt aor22d1 GND Y VDD A B D C
M1 GND C N_7 GND mn15  l=0.13u w=0.26u m=1
M2 N_2 D N_7 GND mn15  l=0.13u w=0.26u m=1
M3 N_8 B N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_13 C N_2 VDD mp15  l=0.13u w=0.4u m=1
M7 N_13 D N_2 VDD mp15  l=0.13u w=0.4u m=1
M8 N_13 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor22d1
* SPICE INPUT		Tue Jul 31 18:51:26 2018	aor22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d2
.subckt aor22d2 Y GND VDD A B D C
M1 N_8 B N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND C N_9 GND mn15  l=0.13u w=0.46u m=1
M6 N_4 D N_9 GND mn15  l=0.13u w=0.46u m=1
M7 N_14 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M8 N_4 D N_14 VDD mp15  l=0.13u w=0.69u m=1
M9 N_14 B VDD VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_14 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor22d2
* SPICE INPUT		Tue Jul 31 18:51:37 2018	aor22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d4
.subckt aor22d4 GND Y VDD A B C D
M1 N_13 C GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 D N_12 GND mn15  l=0.13u w=0.46u m=1
M3 N_4 D N_13 GND mn15  l=0.13u w=0.46u m=1
M4 N_12 C GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M10 N_15 B N_4 GND mn15  l=0.13u w=0.46u m=1
M11 N_4 B N_14 GND mn15  l=0.13u w=0.46u m=1
M12 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M13 N_4 C N_22 VDD mp15  l=0.13u w=0.69u m=1
M14 N_22 D N_4 VDD mp15  l=0.13u w=0.69u m=1
M15 N_22 D N_4 VDD mp15  l=0.13u w=0.69u m=1
M16 N_22 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M24 VDD A N_22 VDD mp15  l=0.13u w=0.69u m=1
.ends aor22d4
* SPICE INPUT		Tue Jul 31 18:51:50 2018	aor31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d0
.subckt aor31d0 GND Y VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 C N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_12 D N_5 VDD mp15  l=0.13u w=0.4u m=1
M7 N_12 C VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_12 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor31d0
* SPICE INPUT		Tue Jul 31 18:52:02 2018	aor31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d1
.subckt aor31d1 GND Y VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 C N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_12 D N_5 VDD mp15  l=0.13u w=0.4u m=1
M7 N_12 C VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_12 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor31d1
* SPICE INPUT		Tue Jul 31 18:52:15 2018	aor31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d2
.subckt aor31d2 Y GND VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_7 C N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_13 D N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_13 C VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_13 B VDD VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor31d2
* SPICE INPUT		Tue Jul 31 18:52:29 2018	aor31d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d4
.subckt aor31d4 GND Y VDD D A B C
M1 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 B N_11 GND mn15  l=0.13u w=0.46u m=1
M3 N_13 C N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C N_12 GND mn15  l=0.13u w=0.46u m=1
M5 N_14 B N_13 GND mn15  l=0.13u w=0.46u m=1
M6 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_3 D GND GND mn15  l=0.13u w=0.46u m=1
M8 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M11 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_20 C VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_20 C VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_3 D N_20 VDD mp15  l=0.13u w=0.69u m=1
M19 N_20 D N_3 VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M23 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor31d4
* SPICE INPUT		Tue Jul 31 18:52:45 2018	bh01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=bh01d1
.subckt bh01d1 VDD Y GND
M1 GND Y N_4 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 N_6 GND mn15  l=0.13u w=0.26u m=1
M3 GND N_4 N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_4 Y VDD VDD mp15  l=0.13u w=0.4u m=1
M5 Y N_4 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends bh01d1
* SPICE INPUT		Tue Jul 31 18:52:59 2018	buffd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd0
.subckt buffd0 GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends buffd0
* SPICE INPUT		Tue Jul 31 18:53:12 2018	buffd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd1
.subckt buffd1 GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd1
* SPICE INPUT		Tue Jul 31 18:53:29 2018	buffd12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd12
.subckt buffd12 Y GND VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M16 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M18 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M20 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd12
* SPICE INPUT		Tue Jul 31 18:53:41 2018	buffd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd16
.subckt buffd16 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M6 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M16 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M17 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M18 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M19 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M20 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M21 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M22 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M23 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M24 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M26 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M28 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M33 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M34 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M36 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M37 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M38 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M40 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M42 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M43 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M44 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd16
* SPICE INPUT		Tue Jul 31 18:53:53 2018	buffd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd2
.subckt buffd2 Y GND VDD A
M1 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M6 VDD A N_4 VDD mp15  l=0.13u w=0.55u m=1
.ends buffd2
* SPICE INPUT		Tue Jul 31 18:54:05 2018	buffd20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd20
.subckt buffd20 Y GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M4 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M6 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M11 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M12 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M13 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M14 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M15 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M16 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M17 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M18 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M19 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M20 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M21 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M22 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M23 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M24 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M25 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M26 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M27 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M28 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M29 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M30 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M31 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M32 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M33 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M34 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M36 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M37 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M38 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M40 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M42 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M43 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M44 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M45 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M46 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M47 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M48 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M49 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M50 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M51 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M52 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M53 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M54 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd20
* SPICE INPUT		Tue Jul 31 18:54:17 2018	buffd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd3
.subckt buffd3 GND Y VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd3
* SPICE INPUT		Tue Jul 31 18:54:29 2018	buffd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd4
.subckt buffd4 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.35u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.34u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M7 VDD A N_5 VDD mp15  l=0.13u w=0.54u m=1
M8 N_5 A VDD VDD mp15  l=0.13u w=0.54u m=1
M9 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd4
* SPICE INPUT		Tue Jul 31 18:54:40 2018	buffd5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd5
.subckt buffd5 GND Y VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M8 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M9 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd5
* SPICE INPUT		Tue Jul 31 18:54:52 2018	buffd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd6
.subckt buffd6 Y GND VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd6
* SPICE INPUT		Tue Jul 31 18:55:04 2018	buffd7
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd7
.subckt buffd7 GND Y VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.4u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.39u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.39u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 VDD A N_5 VDD mp15  l=0.13u w=0.6u m=1
M12 N_5 A VDD VDD mp15  l=0.13u w=0.6u m=1
M13 VDD A N_5 VDD mp15  l=0.13u w=0.6u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd7
* SPICE INPUT		Tue Jul 31 18:55:15 2018	buffd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd8
.subckt buffd8 Y GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M11 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M12 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M13 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd8
* SPICE INPUT		Tue Jul 31 18:55:27 2018	buffdm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffdm
.subckt buffdm VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends buffdm
* SPICE INPUT		Tue Jul 31 18:55:40 2018	buftd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd0
.subckt buftd0 GND Y VDD E A
M1 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_6 N_7 GND mn15  l=0.13u w=0.5u m=1
M4 Y E N_7 GND mn15  l=0.13u w=0.5u m=1
M5 VDD A N_6 VDD mp15  l=0.13u w=0.4u m=1
M6 N_14 N_6 VDD VDD mp15  l=0.13u w=0.53u m=1
M7 N_15 N_3 Y VDD mp15  l=0.13u w=0.27u m=1
M8 N_14 N_3 Y VDD mp15  l=0.13u w=0.53u m=1
M9 N_15 N_6 VDD VDD mp15  l=0.13u w=0.27u m=1
M10 N_3 E VDD VDD mp15  l=0.13u w=0.4u m=1
.ends buftd0
* SPICE INPUT		Tue Jul 31 18:55:54 2018	buftd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd1
.subckt buftd1 VDD Y GND E A
M1 N_4 A GND GND mn15  l=0.13u w=0.32u m=1
M2 N_14 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_15 E Y GND mn15  l=0.13u w=0.46u m=1
M4 Y E N_14 GND mn15  l=0.13u w=0.46u m=1
M5 N_15 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 E GND GND mn15  l=0.13u w=0.32u m=1
M7 VDD A N_4 VDD mp15  l=0.13u w=0.48u m=1
M8 N_7 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_8 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y N_3 N_7 VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_3 E VDD VDD mp15  l=0.13u w=0.48u m=1
.ends buftd1
* SPICE INPUT		Tue Jul 31 18:56:09 2018	buftd12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd12
.subckt buftd12 GND Y VDD A E
M1 N_5 E GND GND mn15  l=0.13u w=0.42u m=1
M2 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 A GND GND mn15  l=0.13u w=0.42u m=1
M7 N_2 E N_3 GND mn15  l=0.13u w=0.4u m=1
M8 N_2 E N_3 GND mn15  l=0.13u w=0.4u m=1
M9 N_3 E N_2 GND mn15  l=0.13u w=0.4u m=1
M10 N_3 N_5 GND GND mn15  l=0.13u w=0.38u m=1
M11 N_3 N_5 GND GND mn15  l=0.13u w=0.38u m=1
M12 N_3 N_5 GND GND mn15  l=0.13u w=0.38u m=1
M13 Y N_3 GND GND mn15  l=0.13u w=0.425u m=1
M14 Y N_3 GND GND mn15  l=0.13u w=0.425u m=1
M15 Y N_3 GND GND mn15  l=0.13u w=0.425u m=1
M16 GND N_3 Y GND mn15  l=0.13u w=0.425u m=1
M17 Y N_3 GND GND mn15  l=0.13u w=0.405u m=1
M18 Y N_3 GND GND mn15  l=0.13u w=0.455u m=1
M19 Y N_3 GND GND mn15  l=0.13u w=0.455u m=1
M20 Y N_3 GND GND mn15  l=0.13u w=0.455u m=1
M21 Y N_3 GND GND mn15  l=0.13u w=0.455u m=1
M22 Y N_3 GND GND mn15  l=0.13u w=0.4u m=1
M23 Y N_3 GND GND mn15  l=0.13u w=0.4u m=1
M24 GND N_3 Y GND mn15  l=0.13u w=0.4u m=1
M25 Y N_3 GND GND mn15  l=0.13u w=0.365u m=1
M26 VDD E N_5 VDD mp15  l=0.13u w=0.315u m=1
M27 N_5 E VDD VDD mp15  l=0.13u w=0.315u m=1
M28 N_2 A VDD VDD mp15  l=0.13u w=0.685u m=1
M29 N_2 A VDD VDD mp15  l=0.13u w=0.685u m=1
M30 N_2 A VDD VDD mp15  l=0.13u w=0.685u m=1
M31 N_2 A VDD VDD mp15  l=0.13u w=0.685u m=1
M32 N_2 A VDD VDD mp15  l=0.13u w=0.56u m=1
M33 N_2 E VDD VDD mp15  l=0.13u w=0.605u m=1
M34 N_2 E VDD VDD mp15  l=0.13u w=0.605u m=1
M35 VDD E N_2 VDD mp15  l=0.13u w=0.465u m=1
M36 N_2 N_5 N_3 VDD mp15  l=0.13u w=0.79u m=1
M37 N_3 N_5 N_2 VDD mp15  l=0.13u w=0.8u m=1
M38 N_3 N_5 N_2 VDD mp15  l=0.13u w=0.79u m=1
M39 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M40 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M41 Y N_2 VDD VDD mp15  l=0.13u w=0.71u m=1
M42 Y N_2 VDD VDD mp15  l=0.13u w=0.71u m=1
M43 VDD N_2 Y VDD mp15  l=0.13u w=0.71u m=1
M44 Y N_2 VDD VDD mp15  l=0.13u w=0.71u m=1
M45 VDD N_2 Y VDD mp15  l=0.13u w=0.71u m=1
M46 Y N_2 VDD VDD mp15  l=0.13u w=0.71u m=1
M47 VDD N_2 Y VDD mp15  l=0.13u w=0.71u m=1
M48 Y N_2 VDD VDD mp15  l=0.13u w=0.68u m=1
M49 VDD N_2 Y VDD mp15  l=0.13u w=0.67u m=1
M50 Y N_2 VDD VDD mp15  l=0.13u w=0.58u m=1
.ends buftd12
* SPICE INPUT		Tue Jul 31 18:56:22 2018	buftd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd16
.subckt buftd16 GND Y VDD E A
M1 GND A N_2 GND mn15  l=0.13u w=0.43u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M3 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M4 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M5 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M6 N_2 A GND GND mn15  l=0.13u w=0.4u m=1
M7 N_2 A GND GND mn15  l=0.13u w=0.37u m=1
M8 N_2 N_14 GND GND mn15  l=0.13u w=0.37u m=1
M9 N_2 N_14 GND GND mn15  l=0.13u w=0.37u m=1
M10 GND N_14 N_2 GND mn15  l=0.13u w=0.37u m=1
M11 GND N_14 N_2 GND mn15  l=0.13u w=0.35u m=1
M12 GND E N_14 GND mn15  l=0.13u w=0.44u m=1
M13 N_17 E N_2 GND mn15  l=0.13u w=0.55u m=1
M14 N_2 E N_17 GND mn15  l=0.13u w=0.55u m=1
M15 N_2 E N_17 GND mn15  l=0.13u w=0.48u m=1
M16 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M17 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M18 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M19 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M20 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M21 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M22 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M23 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M24 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M25 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M26 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M27 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M28 Y N_2 GND GND mn15  l=0.13u w=0.4u m=1
M29 Y N_2 GND GND mn15  l=0.13u w=0.4u m=1
M30 GND N_2 Y GND mn15  l=0.13u w=0.4u m=1
M31 Y N_2 GND GND mn15  l=0.13u w=0.4u m=1
M32 Y N_2 GND GND mn15  l=0.13u w=0.36u m=1
M33 N_17 A VDD VDD mp15  l=0.13u w=0.65u m=1
M34 VDD A N_17 VDD mp15  l=0.13u w=0.65u m=1
M35 N_17 A VDD VDD mp15  l=0.13u w=0.65u m=1
M36 VDD A N_17 VDD mp15  l=0.13u w=0.65u m=1
M37 N_17 A VDD VDD mp15  l=0.13u w=0.65u m=1
M38 VDD A N_17 VDD mp15  l=0.13u w=0.65u m=1
M39 N_17 A VDD VDD mp15  l=0.13u w=0.64u m=1
M40 N_17 E VDD VDD mp15  l=0.13u w=0.76u m=1
M41 N_17 E VDD VDD mp15  l=0.13u w=0.76u m=1
M42 VDD E N_17 VDD mp15  l=0.13u w=0.73u m=1
M43 N_14 E VDD VDD mp15  l=0.13u w=0.67u m=1
M44 N_2 N_14 N_17 VDD mp15  l=0.13u w=0.56u m=1
M45 N_17 N_14 N_2 VDD mp15  l=0.13u w=0.56u m=1
M46 N_17 N_14 N_2 VDD mp15  l=0.13u w=0.56u m=1
M47 N_2 N_14 N_17 VDD mp15  l=0.13u w=0.56u m=1
M48 N_17 N_14 N_2 VDD mp15  l=0.13u w=0.56u m=1
M49 N_2 N_14 N_17 VDD mp15  l=0.13u w=0.28u m=1
M50 Y N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M51 Y N_17 VDD VDD mp15  l=0.13u w=0.67u m=1
M52 Y N_17 VDD VDD mp15  l=0.13u w=0.67u m=1
M53 VDD N_17 Y VDD mp15  l=0.13u w=0.67u m=1
M54 Y N_17 VDD VDD mp15  l=0.13u w=0.67u m=1
M55 VDD N_17 Y VDD mp15  l=0.13u w=0.69u m=1
M56 VDD N_17 Y VDD mp15  l=0.13u w=0.69u m=1
M57 Y N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M58 VDD N_17 Y VDD mp15  l=0.13u w=0.69u m=1
M59 Y N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M60 VDD N_17 Y VDD mp15  l=0.13u w=0.69u m=1
M61 Y N_17 VDD VDD mp15  l=0.13u w=0.65u m=1
M62 Y N_17 VDD VDD mp15  l=0.13u w=0.62u m=1
M63 VDD N_17 Y VDD mp15  l=0.13u w=0.57u m=1
M64 Y N_17 VDD VDD mp15  l=0.13u w=0.57u m=1
M65 VDD N_17 Y VDD mp15  l=0.13u w=0.57u m=1
M66 Y N_17 VDD VDD mp15  l=0.13u w=0.57u m=1
.ends buftd16
* SPICE INPUT		Tue Jul 31 18:56:36 2018	buftd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd2
.subckt buftd2 GND Y VDD E A
M1 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 E GND GND mn15  l=0.13u w=0.46u m=1
M3 N_6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_6 E Y GND mn15  l=0.13u w=0.565u m=1
M8 N_6 E Y GND mn15  l=0.13u w=0.565u m=1
M9 N_6 E Y GND mn15  l=0.13u w=0.43u m=1
M10 Y E N_6 GND mn15  l=0.13u w=0.29u m=1
M11 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD E N_3 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_4 N_15 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_4 N_15 VDD mp15  l=0.13u w=0.69u m=1
M15 N_15 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_4 N_15 VDD mp15  l=0.13u w=0.69u m=1
M17 Y N_3 N_15 VDD mp15  l=0.13u w=0.595u m=1
M18 Y N_3 N_15 VDD mp15  l=0.13u w=0.595u m=1
M19 Y N_3 N_15 VDD mp15  l=0.13u w=0.595u m=1
M20 N_15 N_3 Y VDD mp15  l=0.13u w=0.595u m=1
M21 Y N_3 N_15 VDD mp15  l=0.13u w=0.46u m=1
.ends buftd2
* SPICE INPUT		Tue Jul 31 18:56:52 2018	buftd20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd20
.subckt buftd20 GND Y VDD E A
M1 N_5 N_2 GND GND mn15  l=0.13u w=0.47u m=1
M2 N_5 N_2 GND GND mn15  l=0.13u w=0.47u m=1
M3 GND N_2 N_5 GND mn15  l=0.13u w=0.47u m=1
M4 N_5 N_2 GND GND mn15  l=0.13u w=0.47u m=1
M5 GND E N_2 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M8 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M9 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M10 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M11 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M12 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M13 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M14 N_5 E N_16 GND mn15  l=0.13u w=0.56u m=1
M15 N_5 E N_16 GND mn15  l=0.13u w=0.56u m=1
M16 N_5 E N_16 GND mn15  l=0.13u w=0.56u m=1
M17 N_16 E N_5 GND mn15  l=0.13u w=0.32u m=1
M18 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M19 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M20 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M21 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M22 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M23 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M24 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M25 Y N_5 GND GND mn15  l=0.13u w=0.39u m=1
M26 Y N_5 GND GND mn15  l=0.13u w=0.39u m=1
M27 Y N_5 GND GND mn15  l=0.13u w=0.27u m=1
M28 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M29 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M30 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M31 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M32 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M33 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M34 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M35 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M36 Y N_5 GND GND mn15  l=0.13u w=0.39u m=1
M37 Y N_5 GND GND mn15  l=0.13u w=0.39u m=1
M38 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M39 N_2 E VDD VDD mp15  l=0.13u w=0.69u m=1
M40 N_16 E VDD VDD mp15  l=0.13u w=0.69u m=1
M41 N_16 E VDD VDD mp15  l=0.13u w=0.69u m=1
M42 VDD E N_16 VDD mp15  l=0.13u w=0.69u m=1
M43 N_16 E VDD VDD mp15  l=0.13u w=0.69u m=1
M44 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M45 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M46 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M47 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M48 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M49 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M50 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M51 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M52 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.575u m=1
M53 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.575u m=1
M54 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.575u m=1
M55 N_16 N_2 N_5 VDD mp15  l=0.13u w=0.575u m=1
M56 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.57u m=1
M57 N_16 N_2 N_5 VDD mp15  l=0.13u w=0.57u m=1
M58 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.42u m=1
M59 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M60 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M61 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M62 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M63 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M64 Y N_16 VDD VDD mp15  l=0.13u w=0.64u m=1
M65 Y N_16 VDD VDD mp15  l=0.13u w=0.64u m=1
M66 VDD N_16 Y VDD mp15  l=0.13u w=0.64u m=1
M67 Y N_16 VDD VDD mp15  l=0.13u w=0.64u m=1
M68 VDD N_16 Y VDD mp15  l=0.13u w=0.62u m=1
M69 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M70 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M71 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M72 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M73 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M74 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M75 Y N_16 VDD VDD mp15  l=0.13u w=0.6u m=1
M76 VDD N_16 Y VDD mp15  l=0.13u w=0.57u m=1
M77 Y N_16 VDD VDD mp15  l=0.13u w=0.57u m=1
M78 VDD N_16 Y VDD mp15  l=0.13u w=0.57u m=1
M79 Y N_16 VDD VDD mp15  l=0.13u w=0.57u m=1
.ends buftd20
* SPICE INPUT		Tue Jul 31 18:57:04 2018	buftd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd3
.subckt buftd3 GND Y VDD E A
M1 N_5 E GND GND mn15  l=0.13u w=0.3u m=1
M2 N_2 A GND GND mn15  l=0.13u w=0.28u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.27u m=1
M4 GND N_5 N_2 GND mn15  l=0.13u w=0.28u m=1
M5 N_3 E N_2 GND mn15  l=0.13u w=0.3u m=1
M6 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M8 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M9 N_5 E VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_3 A VDD VDD mp15  l=0.13u w=0.83u m=1
M11 N_3 N_5 N_2 VDD mp15  l=0.13u w=0.6u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD E N_3 VDD mp15  l=0.13u w=0.41u m=1
.ends buftd3
* SPICE INPUT		Tue Jul 31 18:57:15 2018	buftd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd4
.subckt buftd4 GND Y VDD E A
M1 N_4 E GND GND mn15  l=0.13u w=0.3u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.37u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.37u m=1
M4 N_6 N_4 GND GND mn15  l=0.13u w=0.37u m=1
M5 N_6 E N_2 GND mn15  l=0.13u w=0.39u m=1
M6 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_4 E VDD VDD mp15  l=0.13u w=0.4u m=1
M11 VDD A N_2 VDD mp15  l=0.13u w=0.55u m=1
M12 N_2 A VDD VDD mp15  l=0.13u w=0.55u m=1
M13 VDD E N_2 VDD mp15  l=0.13u w=0.55u m=1
M14 N_6 N_4 N_2 VDD mp15  l=0.13u w=0.64u m=1
M15 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buftd4
* SPICE INPUT		Tue Jul 31 18:57:27 2018	buftd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd6
.subckt buftd6 GND Y VDD A E
M1 GND E N_4 GND mn15  l=0.13u w=0.3u m=1
M2 GND A N_3 GND mn15  l=0.13u w=0.37u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.37u m=1
M4 N_3 A GND GND mn15  l=0.13u w=0.37u m=1
M5 N_3 E N_2 GND mn15  l=0.13u w=0.59u m=1
M6 N_3 N_4 GND GND mn15  l=0.13u w=0.55u m=1
M7 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M13 VDD E N_4 VDD mp15  l=0.13u w=0.42u m=1
M14 N_2 A VDD VDD mp15  l=0.13u w=0.66u m=1
M15 N_2 A VDD VDD mp15  l=0.13u w=0.57u m=1
M16 N_2 A VDD VDD mp15  l=0.13u w=0.45u m=1
M17 N_2 E VDD VDD mp15  l=0.13u w=0.41u m=1
M18 VDD E N_2 VDD mp15  l=0.13u w=0.41u m=1
M19 N_2 N_4 N_3 VDD mp15  l=0.13u w=0.59u m=1
M20 N_3 N_4 N_2 VDD mp15  l=0.13u w=0.57u m=1
M21 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buftd6
* SPICE INPUT		Tue Jul 31 18:57:39 2018	buftd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd8
.subckt buftd8 GND Y VDD E A
M1 N_4 E GND GND mn15  l=0.13u w=0.4u m=1
M2 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_8 E N_2 GND mn15  l=0.13u w=0.42u m=1
M6 N_2 E N_8 GND mn15  l=0.13u w=0.38u m=1
M7 GND N_4 N_2 GND mn15  l=0.13u w=0.35u m=1
M8 GND N_4 N_2 GND mn15  l=0.13u w=0.35u m=1
M9 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M10 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M16 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD E N_4 VDD mp15  l=0.13u w=0.3u m=1
M18 N_4 E VDD VDD mp15  l=0.13u w=0.3u m=1
M19 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_8 E VDD VDD mp15  l=0.13u w=0.595u m=1
M23 VDD E N_8 VDD mp15  l=0.13u w=0.445u m=1
M24 N_2 N_4 N_8 VDD mp15  l=0.13u w=0.81u m=1
M25 N_2 N_4 N_8 VDD mp15  l=0.13u w=0.75u m=1
M26 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M27 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M29 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M31 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M33 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buftd8
* SPICE INPUT		Tue Jul 31 18:57:51 2018	buftdm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftdm
.subckt buftdm VDD Y GND E A
M1 GND A N_5 GND mn15  l=0.13u w=0.26u m=1
M2 N_31 N_5 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_32 N_5 GND GND mn15  l=0.13u w=0.24u m=1
M4 N_31 E Y GND mn15  l=0.13u w=0.46u m=1
M5 N_32 E Y GND mn15  l=0.13u w=0.24u m=1
M6 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M7 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_7 N_5 VDD VDD mp15  l=0.13u w=0.53u m=1
M9 N_8 N_3 Y VDD mp15  l=0.13u w=0.53u m=1
M10 Y N_3 N_7 VDD mp15  l=0.13u w=0.53u m=1
M11 N_8 N_5 VDD VDD mp15  l=0.13u w=0.53u m=1
M12 N_3 E VDD VDD mp15  l=0.13u w=0.4u m=1
.ends buftdm
* SPICE INPUT		Tue Jul 31 18:58:03 2018	ckandd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckandd0
.subckt ckandd0 Y GND VDD A B
M1 GND N_4 Y GND mn15  l=0.13u w=0.2u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.2u m=1
M3 N_5 B N_4 GND mn15  l=0.13u w=0.2u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.5u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.5u m=1
.ends ckandd0
* SPICE INPUT		Tue Jul 31 18:58:15 2018	ckandd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckandd1
.subckt ckandd1 GND Y VDD A B
M1 Y N_4 GND GND mn15  l=0.13u w=0.39u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_5 B N_4 GND mn15  l=0.13u w=0.26u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.59u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.59u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.6u m=1
M7 N_4 B VDD VDD mp15  l=0.13u w=0.6u m=1
.ends ckandd1
* SPICE INPUT		Tue Jul 31 18:58:27 2018	ckandd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckandd2
.subckt ckandd2 GND Y VDD A B
M1 N_5 A GND GND mn15  l=0.13u w=0.3u m=1
M2 N_5 B N_4 GND mn15  l=0.13u w=0.3u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M5 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M6 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckandd2
* SPICE INPUT		Tue Jul 31 18:58:39 2018	ckandd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckandd4
.subckt ckandd4 Y GND VDD A B
M1 GND A N_9 GND mn15  l=0.13u w=0.33u m=1
M2 Y N_5 GND GND mn15  l=0.13u w=0.265u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.265u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.265u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.265u m=1
M6 GND A N_10 GND mn15  l=0.13u w=0.27u m=1
M7 N_5 B N_10 GND mn15  l=0.13u w=0.3u m=1
M8 N_5 B N_9 GND mn15  l=0.13u w=0.3u m=1
M9 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.865u m=1
M11 Y N_5 VDD VDD mp15  l=0.13u w=0.865u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.79u m=1
M13 Y N_5 VDD VDD mp15  l=0.13u w=0.24u m=1
M14 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M15 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M16 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends ckandd4
* SPICE INPUT		Tue Jul 31 18:58:51 2018	ckbufd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd0
.subckt ckbufd0 VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.2u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd0
* SPICE INPUT		Tue Jul 31 18:59:05 2018	ckbufd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd1
.subckt ckbufd1 GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.4u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
.ends ckbufd1
* SPICE INPUT		Tue Jul 31 18:59:19 2018	ckbufd10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd10
.subckt ckbufd10 GND Y VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M2 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.35u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_4 A VDD VDD mp15  l=0.13u w=0.735u m=1
M11 VDD A N_4 VDD mp15  l=0.13u w=0.72u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.72u m=1
M13 N_4 A VDD VDD mp15  l=0.13u w=0.705u m=1
M14 Y N_4 VDD VDD mp15  l=0.13u w=1.38u m=1
M15 Y N_4 VDD VDD mp15  l=0.13u w=0.795u m=1
M16 VDD N_4 Y VDD mp15  l=0.13u w=0.72u m=1
M17 Y N_4 VDD VDD mp15  l=0.13u w=0.72u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.72u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.72u m=1
M20 VDD N_4 Y VDD mp15  l=0.13u w=0.72u m=1
M21 Y N_4 VDD VDD mp15  l=0.13u w=0.72u m=1
M22 Y N_4 VDD VDD mp15  l=0.13u w=0.71u m=1
.ends ckbufd10
* SPICE INPUT		Tue Jul 31 18:59:34 2018	ckbufd12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd12
.subckt ckbufd12 Y GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M2 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.35u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M6 Y N_4 GND GND mn15  l=0.13u w=0.41u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.41u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M11 Y N_4 GND GND mn15  l=0.13u w=0.41u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.73u m=1
M13 N_4 A VDD VDD mp15  l=0.13u w=0.72u m=1
M14 N_4 A VDD VDD mp15  l=0.13u w=0.72u m=1
M15 N_4 A VDD VDD mp15  l=0.13u w=0.67u m=1
M16 Y N_4 VDD VDD mp15  l=0.13u w=1.23u m=1
M17 Y N_4 VDD VDD mp15  l=0.13u w=0.91u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.71u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
M21 VDD N_4 Y VDD mp15  l=0.13u w=0.695u m=1
M22 Y N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
M23 VDD N_4 Y VDD mp15  l=0.13u w=0.695u m=1
M24 Y N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
M25 VDD N_4 Y VDD mp15  l=0.13u w=0.695u m=1
M26 Y N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
.ends ckbufd12
* SPICE INPUT		Tue Jul 31 18:59:47 2018	ckbufd14
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd14
.subckt ckbufd14 GND Y VDD A
M1 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.44u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.44u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.43u m=1
M8 Y N_4 GND GND mn15  l=0.13u w=0.43u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.43u m=1
M10 GND A N_4 GND mn15  l=0.13u w=0.44u m=1
M11 N_4 A GND GND mn15  l=0.13u w=0.435u m=1
M12 GND A N_4 GND mn15  l=0.13u w=0.435u m=1
M13 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M14 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M15 Y N_4 VDD VDD mp15  l=0.13u w=0.8u m=1
M16 VDD N_4 Y VDD mp15  l=0.13u w=0.735u m=1
M17 Y N_4 VDD VDD mp15  l=0.13u w=0.735u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.735u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.725u m=1
M20 VDD N_4 Y VDD mp15  l=0.13u w=0.725u m=1
M21 Y N_4 VDD VDD mp15  l=0.13u w=0.725u m=1
M22 VDD N_4 Y VDD mp15  l=0.13u w=0.725u m=1
M23 Y N_4 VDD VDD mp15  l=0.13u w=0.725u m=1
M24 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M25 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M26 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M27 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M28 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M29 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd14
* SPICE INPUT		Tue Jul 31 19:00:03 2018	ckbufd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd16
.subckt ckbufd16 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.405u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.405u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.405u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.405u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 VDD A N_5 VDD mp15  l=0.13u w=0.72u m=1
M15 VDD A N_5 VDD mp15  l=0.13u w=0.72u m=1
M16 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M18 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M21 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M22 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M23 Y N_5 VDD VDD mp15  l=0.13u w=0.785u m=1
M24 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M25 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M26 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M27 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M28 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M29 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M30 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M31 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M32 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
.ends ckbufd16
* SPICE INPUT		Tue Jul 31 19:00:16 2018	ckbufd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd2
.subckt ckbufd2 GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd2
* SPICE INPUT		Tue Jul 31 19:00:27 2018	ckbufd20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd20
.subckt ckbufd20 GND Y VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M10 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M16 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M18 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M21 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M23 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M25 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M26 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M27 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M28 Y N_5 VDD VDD mp15  l=0.13u w=0.83u m=1
M29 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M30 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M31 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
M32 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M33 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
M34 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M35 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
M36 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M37 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
M38 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M39 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
.ends ckbufd20
* SPICE INPUT		Tue Jul 31 19:00:39 2018	ckbufd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd3
.subckt ckbufd3 GND Y VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.2u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M5 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd3
* SPICE INPUT		Tue Jul 31 19:00:51 2018	ckbufd30
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd30
.subckt ckbufd30 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.41u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.41u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.41u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.41u m=1
M5 GND A N_5 GND mn15  l=0.13u w=0.41u m=1
M6 N_5 A GND GND mn15  l=0.13u w=0.41u m=1
M7 GND A N_5 GND mn15  l=0.13u w=0.41u m=1
M8 N_5 A GND GND mn15  l=0.13u w=0.41u m=1
M9 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M10 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M11 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M12 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M13 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M14 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M15 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M16 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M17 Y N_5 GND GND mn15  l=0.13u w=0.44u m=1
M18 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M19 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M20 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M21 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M22 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M23 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M24 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M25 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M26 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M27 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M28 N_5 A VDD VDD mp15  l=0.13u w=0.71u m=1
M29 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M30 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M31 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M32 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M33 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M34 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M35 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M36 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M37 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M38 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M39 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M40 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M41 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M42 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M43 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M44 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M45 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M46 Y N_5 VDD VDD mp15  l=0.13u w=0.875u m=1
M47 VDD N_5 Y VDD mp15  l=0.13u w=0.725u m=1
M48 Y N_5 VDD VDD mp15  l=0.13u w=0.725u m=1
M49 VDD N_5 Y VDD mp15  l=0.13u w=0.725u m=1
M50 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M51 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M52 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M53 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M54 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M55 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M56 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M57 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M58 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M59 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M60 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M61 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M62 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M63 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
.ends ckbufd30
* SPICE INPUT		Tue Jul 31 19:01:03 2018	ckbufd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd4
.subckt ckbufd4 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.26u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.23u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.27u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.27u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.27u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_5 A VDD VDD mp15  l=0.13u w=0.71u m=1
M8 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_5 Y VDD mp15  l=0.13u w=0.7u m=1
M10 VDD N_5 Y VDD mp15  l=0.13u w=0.7u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.7u m=1
M12 Y N_5 VDD VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd4
* SPICE INPUT		Tue Jul 31 19:01:15 2018	ckbufd40
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd40
.subckt ckbufd40 GND Y VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M2 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M3 N_4 A GND GND mn15  l=0.13u w=0.43u m=1
M4 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M5 N_4 A GND GND mn15  l=0.13u w=0.43u m=1
M6 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M7 N_4 A GND GND mn15  l=0.13u w=0.43u m=1
M8 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M9 GND A N_4 GND mn15  l=0.13u w=0.4u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M11 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M12 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M13 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M14 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M15 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M16 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M17 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M18 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M19 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M20 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M21 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M22 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M23 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M24 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M25 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M26 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M27 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M28 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M29 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M30 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M31 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M32 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M33 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M34 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M35 N_4 A VDD VDD mp15  l=0.13u w=0.71u m=1
M36 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M37 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M38 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M39 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M40 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M41 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M42 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M43 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M44 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M45 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M46 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M47 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M48 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M49 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M50 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M51 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M52 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M53 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M54 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M55 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M56 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M57 VDD N_4 Y VDD mp15  l=0.13u w=1.28u m=1
M58 VDD N_4 Y VDD mp15  l=0.13u w=0.705u m=1
M59 Y N_4 VDD VDD mp15  l=0.13u w=0.705u m=1
M60 VDD N_4 Y VDD mp15  l=0.13u w=0.705u m=1
M61 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M62 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M63 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M64 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M65 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M66 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M67 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M68 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M69 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M70 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M71 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M72 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M73 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M74 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M75 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M76 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M77 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M78 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M79 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M80 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd40
* SPICE INPUT		Tue Jul 31 19:01:27 2018	ckbufd5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd5
.subckt ckbufd5 GND Y VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.26u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.27u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.27u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.27u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.27u m=1
M7 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M8 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M9 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd5
* SPICE INPUT		Tue Jul 31 19:01:39 2018	ckbufd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd6
.subckt ckbufd6 Y GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.44u m=1
M2 GND A N_4 GND mn15  l=0.13u w=0.32u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.27u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.27u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.27u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.27u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.27u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.27u m=1
M9 VDD A N_4 VDD mp15  l=0.13u w=0.72u m=1
M10 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_4 VDD VDD mp15  l=0.13u w=0.88u m=1
M13 Y N_4 VDD VDD mp15  l=0.13u w=0.88u m=1
M14 VDD N_4 Y VDD mp15  l=0.13u w=0.88u m=1
M15 Y N_4 VDD VDD mp15  l=0.13u w=0.88u m=1
M16 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd6
* SPICE INPUT		Tue Jul 31 19:01:51 2018	ckbufd7
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd7
.subckt ckbufd7 GND Y VDD A
M1 N_6 A GND GND mn15  l=0.13u w=0.39u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.39u m=1
M3 Y N_6 GND GND mn15  l=0.13u w=0.27u m=1
M4 GND N_6 Y GND mn15  l=0.13u w=0.26u m=1
M5 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M6 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M7 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M8 GND N_6 Y GND mn15  l=0.13u w=0.26u m=1
M9 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M10 VDD A N_6 VDD mp15  l=0.13u w=0.705u m=1
M11 N_6 A VDD VDD mp15  l=0.13u w=0.705u m=1
M12 VDD A N_6 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.89u m=1
M14 VDD N_6 Y VDD mp15  l=0.13u w=0.89u m=1
M15 Y N_6 VDD VDD mp15  l=0.13u w=0.89u m=1
M16 VDD N_6 Y VDD mp15  l=0.13u w=0.775u m=1
M17 Y N_6 VDD VDD mp15  l=0.13u w=0.775u m=1
M18 VDD N_6 Y VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd7
* SPICE INPUT		Tue Jul 31 19:02:03 2018	ckbufd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd8
.subckt ckbufd8 Y GND VDD A
M1 N_6 A GND GND mn15  l=0.13u w=0.39u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.39u m=1
M3 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M4 Y N_6 GND GND mn15  l=0.13u w=0.27u m=1
M5 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M6 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M7 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M8 Y N_6 GND GND mn15  l=0.13u w=0.27u m=1
M9 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M10 Y N_6 GND GND mn15  l=0.13u w=0.27u m=1
M11 VDD A N_6 VDD mp15  l=0.13u w=0.755u m=1
M12 N_6 A VDD VDD mp15  l=0.13u w=0.7u m=1
M13 VDD A N_6 VDD mp15  l=0.13u w=0.7u m=1
M14 Y N_6 VDD VDD mp15  l=0.13u w=0.825u m=1
M15 VDD N_6 Y VDD mp15  l=0.13u w=0.895u m=1
M16 VDD N_6 Y VDD mp15  l=0.13u w=0.895u m=1
M17 Y N_6 VDD VDD mp15  l=0.13u w=0.895u m=1
M18 VDD N_6 Y VDD mp15  l=0.13u w=0.775u m=1
M19 Y N_6 VDD VDD mp15  l=0.13u w=0.775u m=1
M20 Y N_6 VDD VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd8
* SPICE INPUT		Tue Jul 31 19:02:16 2018	ckbufd80
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd80
.subckt ckbufd80 GND Y VDD A
M1 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M2 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M3 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M4 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M5 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M6 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M7 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M8 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M9 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M10 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M12 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M13 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M14 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M15 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M16 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M17 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M18 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M19 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M20 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M21 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M22 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M23 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M24 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M25 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M26 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M27 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M28 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M29 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M30 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M31 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M32 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M33 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M34 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M35 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M36 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M37 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M38 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M39 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M40 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M41 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M42 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M43 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M44 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M45 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M46 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M47 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M48 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M49 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M50 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M51 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M52 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M53 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M54 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M55 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M56 Y N_2 GND GND mn15  l=0.13u w=0.44u m=1
M57 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M58 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M59 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M60 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M61 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M62 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M63 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M64 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M65 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M66 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M67 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M68 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M69 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M70 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M71 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M72 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M73 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M74 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M75 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M76 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M77 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M78 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M79 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M80 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M81 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M82 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M83 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M84 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M85 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M86 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M87 VDD N_2 Y VDD mp15  l=0.13u w=1.28u m=1
M88 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M89 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M90 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M91 Y N_2 VDD VDD mp15  l=0.13u w=0.715u m=1
M92 VDD N_2 Y VDD mp15  l=0.13u w=0.715u m=1
M93 VDD N_2 Y VDD mp15  l=0.13u w=0.715u m=1
M94 VDD N_2 Y VDD mp15  l=0.13u w=0.71u m=1
M95 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M96 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M97 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M98 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M99 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M100 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M101 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M102 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M103 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M104 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M105 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M106 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M107 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M108 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M109 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M110 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M111 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M112 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M113 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M114 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M115 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M116 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M117 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M118 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M119 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M120 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M121 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M122 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M123 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M124 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M125 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M126 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M127 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M128 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M129 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M130 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M131 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M132 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M133 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M134 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M135 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M136 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M137 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M138 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M139 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M140 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M141 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M142 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M143 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M144 VDD A N_2 VDD mp15  l=0.13u w=0.71u m=1
M145 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M146 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M147 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M148 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M149 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M150 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M151 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M152 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M153 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M154 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M155 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M156 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M157 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M158 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M159 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M160 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M161 N_2 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd80
* SPICE INPUT		Tue Jul 31 19:02:31 2018	ckbufdm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufdm
.subckt ckbufdm GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.3u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.37u m=1
.ends ckbufdm
* SPICE INPUT		Tue Jul 31 19:02:46 2018	ckinvd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd0
.subckt ckinvd0 GND VDD Y A
M1 GND A Y GND mn15  l=0.13u w=0.2u m=1
M2 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd0
* SPICE INPUT		Tue Jul 31 19:03:00 2018	ckinvd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd1
.subckt ckinvd1 Y VDD GND A
M1 Y A GND GND mn15  l=0.13u w=0.4u m=1
M2 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
.ends ckinvd1
* SPICE INPUT		Tue Jul 31 19:03:15 2018	ckinvd10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd10
.subckt ckinvd10 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.3u m=1
M2 Y A GND GND mn15  l=0.13u w=0.3u m=1
M3 Y A GND GND mn15  l=0.13u w=0.3u m=1
M4 Y A GND GND mn15  l=0.13u w=0.295u m=1
M5 Y A GND GND mn15  l=0.13u w=0.295u m=1
M6 Y A GND GND mn15  l=0.13u w=0.295u m=1
M7 Y A GND GND mn15  l=0.13u w=0.295u m=1
M8 Y A GND GND mn15  l=0.13u w=0.295u m=1
M9 GND A Y GND mn15  l=0.13u w=0.295u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.805u m=1
M11 Y A VDD VDD mp15  l=0.13u w=0.805u m=1
M12 VDD A Y VDD mp15  l=0.13u w=0.805u m=1
M13 Y A VDD VDD mp15  l=0.13u w=0.805u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.805u m=1
M15 Y A VDD VDD mp15  l=0.13u w=0.805u m=1
M16 VDD A Y VDD mp15  l=0.13u w=0.805u m=1
M17 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 Y A VDD VDD mp15  l=0.13u w=0.685u m=1
.ends ckinvd10
* SPICE INPUT		Tue Jul 31 19:03:31 2018	ckinvd12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd12
.subckt ckinvd12 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.3u m=1
M2 Y A GND GND mn15  l=0.13u w=0.295u m=1
M3 Y A GND GND mn15  l=0.13u w=0.295u m=1
M4 Y A GND GND mn15  l=0.13u w=0.295u m=1
M5 GND A Y GND mn15  l=0.13u w=0.295u m=1
M6 Y A GND GND mn15  l=0.13u w=0.295u m=1
M7 GND A Y GND mn15  l=0.13u w=0.295u m=1
M8 Y A GND GND mn15  l=0.13u w=0.295u m=1
M9 GND A Y GND mn15  l=0.13u w=0.295u m=1
M10 Y A GND GND mn15  l=0.13u w=0.295u m=1
M11 GND A Y GND mn15  l=0.13u w=0.295u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.79u m=1
M13 Y A VDD VDD mp15  l=0.13u w=0.79u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M15 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M16 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M17 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M18 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M19 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M20 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M21 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd12
* SPICE INPUT		Tue Jul 31 19:03:43 2018	ckinvd14
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd14
.subckt ckinvd14 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.345u m=1
M2 GND A Y GND mn15  l=0.13u w=0.315u m=1
M3 Y A GND GND mn15  l=0.13u w=0.315u m=1
M4 Y A GND GND mn15  l=0.13u w=0.315u m=1
M5 Y A GND GND mn15  l=0.13u w=0.315u m=1
M6 Y A GND GND mn15  l=0.13u w=0.315u m=1
M7 Y A GND GND mn15  l=0.13u w=0.315u m=1
M8 Y A GND GND mn15  l=0.13u w=0.315u m=1
M9 Y A GND GND mn15  l=0.13u w=0.315u m=1
M10 Y A GND GND mn15  l=0.13u w=0.315u m=1
M11 Y A GND GND mn15  l=0.13u w=0.315u m=1
M12 Y A GND GND mn15  l=0.13u w=0.315u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M15 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M16 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M17 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M18 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M19 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M20 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M21 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M22 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M23 Y A VDD VDD mp15  l=0.13u w=0.782u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd14
* SPICE INPUT		Tue Jul 31 19:03:55 2018	ckinvd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd16
.subckt ckinvd16 Y GND VDD A
M1 Y A GND GND mn15  l=0.13u w=0.315u m=1
M2 Y A GND GND mn15  l=0.13u w=0.315u m=1
M3 Y A GND GND mn15  l=0.13u w=0.315u m=1
M4 Y A GND GND mn15  l=0.13u w=0.315u m=1
M5 GND A Y GND mn15  l=0.13u w=0.31u m=1
M6 GND A Y GND mn15  l=0.13u w=0.31u m=1
M7 GND A Y GND mn15  l=0.13u w=0.31u m=1
M8 Y A GND GND mn15  l=0.13u w=0.31u m=1
M9 GND A Y GND mn15  l=0.13u w=0.31u m=1
M10 Y A GND GND mn15  l=0.13u w=0.31u m=1
M11 GND A Y GND mn15  l=0.13u w=0.31u m=1
M12 Y A GND GND mn15  l=0.13u w=0.31u m=1
M13 GND A Y GND mn15  l=0.13u w=0.31u m=1
M14 Y A GND GND mn15  l=0.13u w=0.31u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M16 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M17 Y A VDD VDD mp15  l=0.13u w=0.825u m=1
M18 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M19 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M20 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M21 Y A VDD VDD mp15  l=0.13u w=0.82u m=1
M22 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M23 Y A VDD VDD mp15  l=0.13u w=0.82u m=1
M24 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M25 Y A VDD VDD mp15  l=0.13u w=0.82u m=1
M26 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M27 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd16
* SPICE INPUT		Tue Jul 31 19:04:07 2018	ckinvd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd2
.subckt ckinvd2 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.26u m=1
M2 Y A GND GND mn15  l=0.13u w=0.23u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M4 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd2
* SPICE INPUT		Tue Jul 31 19:04:18 2018	ckinvd20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd20
.subckt ckinvd20 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.31u m=1
M2 GND A Y GND mn15  l=0.13u w=0.31u m=1
M3 GND A Y GND mn15  l=0.13u w=0.31u m=1
M4 Y A GND GND mn15  l=0.13u w=0.31u m=1
M5 GND A Y GND mn15  l=0.13u w=0.31u m=1
M6 Y A GND GND mn15  l=0.13u w=0.31u m=1
M7 GND A Y GND mn15  l=0.13u w=0.31u m=1
M8 Y A GND GND mn15  l=0.13u w=0.31u m=1
M9 GND A Y GND mn15  l=0.13u w=0.31u m=1
M10 Y A GND GND mn15  l=0.13u w=0.31u m=1
M11 GND A Y GND mn15  l=0.13u w=0.31u m=1
M12 Y A GND GND mn15  l=0.13u w=0.31u m=1
M13 GND A Y GND mn15  l=0.13u w=0.31u m=1
M14 Y A GND GND mn15  l=0.13u w=0.31u m=1
M15 GND A Y GND mn15  l=0.13u w=0.31u m=1
M16 Y A GND GND mn15  l=0.13u w=0.31u m=1
M17 GND A Y GND mn15  l=0.13u w=0.31u m=1
M18 Y A GND GND mn15  l=0.13u w=0.31u m=1
M19 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M20 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M21 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M23 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M25 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M26 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M27 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M29 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M30 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M31 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M32 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M33 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M34 Y A VDD VDD mp15  l=0.13u w=0.7u m=1
M35 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M36 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M37 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd20
* SPICE INPUT		Tue Jul 31 19:04:30 2018	ckinvd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd3
.subckt ckinvd3 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M5 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd3
* SPICE INPUT		Tue Jul 31 19:04:42 2018	ckinvd30
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd30
.subckt ckinvd30 Y GND VDD A
M1 Y A GND GND mn15  l=0.13u w=0.325u m=1
M2 Y A GND GND mn15  l=0.13u w=0.325u m=1
M3 GND A Y GND mn15  l=0.13u w=0.325u m=1
M4 Y A GND GND mn15  l=0.13u w=0.325u m=1
M5 GND A Y GND mn15  l=0.13u w=0.325u m=1
M6 Y A GND GND mn15  l=0.13u w=0.325u m=1
M7 GND A Y GND mn15  l=0.13u w=0.325u m=1
M8 Y A GND GND mn15  l=0.13u w=0.325u m=1
M9 GND A Y GND mn15  l=0.13u w=0.325u m=1
M10 Y A GND GND mn15  l=0.13u w=0.325u m=1
M11 GND A Y GND mn15  l=0.13u w=0.325u m=1
M12 Y A GND GND mn15  l=0.13u w=0.325u m=1
M13 GND A Y GND mn15  l=0.13u w=0.32u m=1
M14 Y A GND GND mn15  l=0.13u w=0.32u m=1
M15 GND A Y GND mn15  l=0.13u w=0.32u m=1
M16 GND A Y GND mn15  l=0.13u w=0.32u m=1
M17 GND A Y GND mn15  l=0.13u w=0.32u m=1
M18 Y A GND GND mn15  l=0.13u w=0.32u m=1
M19 GND A Y GND mn15  l=0.13u w=0.32u m=1
M20 Y A GND GND mn15  l=0.13u w=0.32u m=1
M21 GND A Y GND mn15  l=0.13u w=0.32u m=1
M22 Y A GND GND mn15  l=0.13u w=0.32u m=1
M23 GND A Y GND mn15  l=0.13u w=0.32u m=1
M24 Y A GND GND mn15  l=0.13u w=0.32u m=1
M25 GND A Y GND mn15  l=0.13u w=0.32u m=1
M26 Y A GND GND mn15  l=0.13u w=0.32u m=1
M27 Y A VDD VDD mp15  l=0.13u w=0.83u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.83u m=1
M29 VDD A Y VDD mp15  l=0.13u w=0.83u m=1
M30 Y A VDD VDD mp15  l=0.13u w=0.83u m=1
M31 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M32 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M33 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M34 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M35 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M36 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M37 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M38 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M39 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M40 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M41 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M42 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M43 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M44 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M45 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M46 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M47 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M48 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M49 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M50 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M51 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M52 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M53 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd30
* SPICE INPUT		Tue Jul 31 19:04:55 2018	ckinvd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd4
.subckt ckinvd4 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.29u m=1
M2 GND A Y GND mn15  l=0.13u w=0.26u m=1
M3 GND A Y GND mn15  l=0.13u w=0.26u m=1
M4 GND A Y GND mn15  l=0.13u w=0.26u m=1
M5 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M6 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd4
* SPICE INPUT		Tue Jul 31 19:05:07 2018	ckinvd40
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd40
.subckt ckinvd40 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.32u m=1
M2 GND A Y GND mn15  l=0.13u w=0.32u m=1
M3 Y A GND GND mn15  l=0.13u w=0.32u m=1
M4 GND A Y GND mn15  l=0.13u w=0.32u m=1
M5 Y A GND GND mn15  l=0.13u w=0.32u m=1
M6 GND A Y GND mn15  l=0.13u w=0.32u m=1
M7 Y A GND GND mn15  l=0.13u w=0.32u m=1
M8 GND A Y GND mn15  l=0.13u w=0.32u m=1
M9 Y A GND GND mn15  l=0.13u w=0.32u m=1
M10 Y A GND GND mn15  l=0.13u w=0.32u m=1
M11 GND A Y GND mn15  l=0.13u w=0.32u m=1
M12 Y A GND GND mn15  l=0.13u w=0.32u m=1
M13 GND A Y GND mn15  l=0.13u w=0.32u m=1
M14 Y A GND GND mn15  l=0.13u w=0.32u m=1
M15 GND A Y GND mn15  l=0.13u w=0.32u m=1
M16 Y A GND GND mn15  l=0.13u w=0.32u m=1
M17 GND A Y GND mn15  l=0.13u w=0.32u m=1
M18 GND A Y GND mn15  l=0.13u w=0.32u m=1
M19 Y A GND GND mn15  l=0.13u w=0.32u m=1
M20 GND A Y GND mn15  l=0.13u w=0.32u m=1
M21 Y A GND GND mn15  l=0.13u w=0.32u m=1
M22 GND A Y GND mn15  l=0.13u w=0.32u m=1
M23 Y A GND GND mn15  l=0.13u w=0.32u m=1
M24 GND A Y GND mn15  l=0.13u w=0.32u m=1
M25 Y A GND GND mn15  l=0.13u w=0.32u m=1
M26 Y A GND GND mn15  l=0.13u w=0.315u m=1
M27 Y A GND GND mn15  l=0.13u w=0.315u m=1
M28 Y A GND GND mn15  l=0.13u w=0.315u m=1
M29 GND A Y GND mn15  l=0.13u w=0.315u m=1
M30 Y A GND GND mn15  l=0.13u w=0.315u m=1
M31 GND A Y GND mn15  l=0.13u w=0.315u m=1
M32 GND A Y GND mn15  l=0.13u w=0.32u m=1
M33 GND A Y GND mn15  l=0.13u w=0.32u m=1
M34 Y A GND GND mn15  l=0.13u w=0.32u m=1
M35 GND A Y GND mn15  l=0.13u w=0.32u m=1
M36 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M37 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M38 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M39 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M40 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M41 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M42 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M43 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M44 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M45 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M46 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M47 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M48 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M49 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M50 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M51 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M52 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M53 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M54 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M55 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M56 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M57 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M58 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M59 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M60 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M61 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M62 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M63 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M64 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M65 Y A VDD VDD mp15  l=0.13u w=0.825u m=1
M66 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M67 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M68 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M69 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M70 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M71 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd40
* SPICE INPUT		Tue Jul 31 19:05:20 2018	ckinvd5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd5
.subckt ckinvd5 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.3u m=1
M2 Y A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y A GND GND mn15  l=0.13u w=0.26u m=1
M5 GND A Y GND mn15  l=0.13u w=0.26u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd5
* SPICE INPUT		Tue Jul 31 19:05:35 2018	ckinvd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd6
.subckt ckinvd6 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.27u m=1
M2 GND A Y GND mn15  l=0.13u w=0.27u m=1
M3 GND A Y GND mn15  l=0.13u w=0.27u m=1
M4 Y A GND GND mn15  l=0.13u w=0.27u m=1
M5 GND A Y GND mn15  l=0.13u w=0.27u m=1
M6 Y A GND GND mn15  l=0.13u w=0.27u m=1
M7 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd6
* SPICE INPUT		Tue Jul 31 19:05:49 2018	ckinvd7
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd7
.subckt ckinvd7 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.28u m=1
M2 Y A GND GND mn15  l=0.13u w=0.27u m=1
M3 Y A GND GND mn15  l=0.13u w=0.27u m=1
M4 Y A GND GND mn15  l=0.13u w=0.27u m=1
M5 GND A Y GND mn15  l=0.13u w=0.27u m=1
M6 Y A GND GND mn15  l=0.13u w=0.27u m=1
M7 GND A Y GND mn15  l=0.13u w=0.27u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd7
* SPICE INPUT		Tue Jul 31 19:06:02 2018	ckinvd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd8
.subckt ckinvd8 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.3u m=1
M2 GND A Y GND mn15  l=0.13u w=0.3u m=1
M3 Y A GND GND mn15  l=0.13u w=0.3u m=1
M4 GND A Y GND mn15  l=0.13u w=0.3u m=1
M5 Y A GND GND mn15  l=0.13u w=0.3u m=1
M6 Y A GND GND mn15  l=0.13u w=0.295u m=1
M7 Y A GND GND mn15  l=0.13u w=0.295u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.85u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.85u m=1
M10 VDD A Y VDD mp15  l=0.13u w=0.85u m=1
M11 Y A VDD VDD mp15  l=0.13u w=0.845u m=1
M12 VDD A Y VDD mp15  l=0.13u w=0.845u m=1
M13 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd8
* SPICE INPUT		Tue Jul 31 19:06:17 2018	ckinvd80
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd80
.subckt ckinvd80 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.315u m=1
M2 Y A GND GND mn15  l=0.13u w=0.315u m=1
M3 GND A Y GND mn15  l=0.13u w=0.315u m=1
M4 Y A GND GND mn15  l=0.13u w=0.315u m=1
M5 GND A Y GND mn15  l=0.13u w=0.315u m=1
M6 Y A GND GND mn15  l=0.13u w=0.315u m=1
M7 GND A Y GND mn15  l=0.13u w=0.315u m=1
M8 Y A GND GND mn15  l=0.13u w=0.315u m=1
M9 GND A Y GND mn15  l=0.13u w=0.315u m=1
M10 GND A Y GND mn15  l=0.13u w=0.315u m=1
M11 GND A Y GND mn15  l=0.13u w=0.27u m=1
M12 Y A GND GND mn15  l=0.13u w=0.27u m=1
M13 GND A Y GND mn15  l=0.13u w=0.27u m=1
M14 Y A GND GND mn15  l=0.13u w=0.27u m=1
M15 GND A Y GND mn15  l=0.13u w=0.275u m=1
M16 Y A GND GND mn15  l=0.13u w=0.315u m=1
M17 GND A Y GND mn15  l=0.13u w=0.315u m=1
M18 Y A GND GND mn15  l=0.13u w=0.315u m=1
M19 Y A GND GND mn15  l=0.13u w=0.315u m=1
M20 GND A Y GND mn15  l=0.13u w=0.325u m=1
M21 GND A Y GND mn15  l=0.13u w=0.325u m=1
M22 Y A GND GND mn15  l=0.13u w=0.325u m=1
M23 Y A GND GND mn15  l=0.13u w=0.325u m=1
M24 GND A Y GND mn15  l=0.13u w=0.325u m=1
M25 Y A GND GND mn15  l=0.13u w=0.325u m=1
M26 GND A Y GND mn15  l=0.13u w=0.325u m=1
M27 Y A GND GND mn15  l=0.13u w=0.325u m=1
M28 GND A Y GND mn15  l=0.13u w=0.325u m=1
M29 Y A GND GND mn15  l=0.13u w=0.325u m=1
M30 GND A Y GND mn15  l=0.13u w=0.325u m=1
M31 GND A Y GND mn15  l=0.13u w=0.325u m=1
M32 GND A Y GND mn15  l=0.13u w=0.325u m=1
M33 Y A GND GND mn15  l=0.13u w=0.325u m=1
M34 GND A Y GND mn15  l=0.13u w=0.325u m=1
M35 Y A GND GND mn15  l=0.13u w=0.325u m=1
M36 GND A Y GND mn15  l=0.13u w=0.325u m=1
M37 Y A GND GND mn15  l=0.13u w=0.325u m=1
M38 Y A GND GND mn15  l=0.13u w=0.325u m=1
M39 Y A GND GND mn15  l=0.13u w=0.325u m=1
M40 GND A Y GND mn15  l=0.13u w=0.325u m=1
M41 Y A GND GND mn15  l=0.13u w=0.325u m=1
M42 Y A GND GND mn15  l=0.13u w=0.325u m=1
M43 Y A GND GND mn15  l=0.13u w=0.325u m=1
M44 GND A Y GND mn15  l=0.13u w=0.325u m=1
M45 Y A GND GND mn15  l=0.13u w=0.325u m=1
M46 GND A Y GND mn15  l=0.13u w=0.325u m=1
M47 Y A GND GND mn15  l=0.13u w=0.325u m=1
M48 GND A Y GND mn15  l=0.13u w=0.325u m=1
M49 Y A GND GND mn15  l=0.13u w=0.325u m=1
M50 Y A GND GND mn15  l=0.13u w=0.325u m=1
M51 GND A Y GND mn15  l=0.13u w=0.325u m=1
M52 Y A GND GND mn15  l=0.13u w=0.325u m=1
M53 GND A Y GND mn15  l=0.13u w=0.325u m=1
M54 Y A GND GND mn15  l=0.13u w=0.325u m=1
M55 GND A Y GND mn15  l=0.13u w=0.325u m=1
M56 Y A GND GND mn15  l=0.13u w=0.325u m=1
M57 Y A GND GND mn15  l=0.13u w=0.325u m=1
M58 GND A Y GND mn15  l=0.13u w=0.325u m=1
M59 Y A GND GND mn15  l=0.13u w=0.325u m=1
M60 GND A Y GND mn15  l=0.13u w=0.325u m=1
M61 Y A GND GND mn15  l=0.13u w=0.325u m=1
M62 GND A Y GND mn15  l=0.13u w=0.325u m=1
M63 Y A GND GND mn15  l=0.13u w=0.325u m=1
M64 GND A Y GND mn15  l=0.13u w=0.325u m=1
M65 Y A GND GND mn15  l=0.13u w=0.325u m=1
M66 GND A Y GND mn15  l=0.13u w=0.325u m=1
M67 Y A GND GND mn15  l=0.13u w=0.325u m=1
M68 GND A Y GND mn15  l=0.13u w=0.325u m=1
M69 Y A GND GND mn15  l=0.13u w=0.325u m=1
M70 GND A Y GND mn15  l=0.13u w=0.325u m=1
M71 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M72 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M73 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M74 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M75 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M76 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M77 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M78 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M79 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M80 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M81 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M82 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M83 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M84 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M85 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M86 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M87 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M88 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M89 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M90 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M91 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M92 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M93 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M94 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M95 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M96 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M97 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M98 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M99 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M100 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M101 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M102 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M103 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M104 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M105 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M106 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M107 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M108 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M109 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M110 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M111 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M112 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M113 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M114 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M115 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M116 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M117 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M118 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M119 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M120 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M121 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M122 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M123 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M124 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M125 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M126 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M127 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M128 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M129 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M130 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M131 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M132 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M133 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M134 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M135 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M136 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M137 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M138 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M139 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M140 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M141 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
.ends ckinvd80
* SPICE INPUT		Tue Jul 31 19:06:32 2018	ckinvdm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvdm
.subckt ckinvdm Y VDD GND A
M1 Y A GND GND mn15  l=0.13u w=0.3u m=1
M2 VDD A Y VDD mp15  l=0.13u w=0.49u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.49u m=1
.ends ckinvdm
* SPICE INPUT		Tue Jul 31 19:06:44 2018	ckmx02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckmx02d0
.subckt ckmx02d0 VDD Y GND S0 B A
M1 N_16 B GND GND mn15  l=0.13u w=0.19u m=1
M2 GND S0 N_3 GND mn15  l=0.13u w=0.18u m=1
M3 N_15 N_3 N_6 GND mn15  l=0.13u w=0.19u m=1
M4 N_15 A GND GND mn15  l=0.13u w=0.19u m=1
M5 GND N_6 Y GND mn15  l=0.13u w=0.19u m=1
M6 N_16 S0 N_6 GND mn15  l=0.13u w=0.19u m=1
M7 N_8 B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_8 N_3 N_6 VDD mp15  l=0.13u w=0.69u m=1
M9 N_3 S0 VDD VDD mp15  l=0.13u w=0.26u m=1
M10 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M12 N_6 S0 N_7 VDD mp15  l=0.13u w=0.69u m=1
.ends ckmx02d0
* SPICE INPUT		Tue Jul 31 19:06:55 2018	ckmx02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckmx02d1
.subckt ckmx02d1 VDD Y GND S0 B A
M1 N_16 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_7 GND GND mn15  l=0.13u w=0.39u m=1
M3 GND S0 N_2 GND mn15  l=0.13u w=0.18u m=1
M4 N_17 B GND GND mn15  l=0.13u w=0.2u m=1
M5 N_7 N_2 N_16 GND mn15  l=0.13u w=0.2u m=1
M6 N_17 S0 N_7 GND mn15  l=0.13u w=0.2u m=1
M7 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_7 Y VDD mp15  l=0.13u w=0.59u m=1
M9 Y N_7 VDD VDD mp15  l=0.13u w=0.59u m=1
M10 VDD S0 N_2 VDD mp15  l=0.13u w=0.24u m=1
M11 N_9 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_9 N_2 N_7 VDD mp15  l=0.13u w=0.69u m=1
M13 N_7 S0 N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends ckmx02d1
* SPICE INPUT		Tue Jul 31 19:07:07 2018	ckmx02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckmx02d2
.subckt ckmx02d2 GND Y VDD S0 B A
M1 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.19u m=1
M3 N_3 S0 GND GND mn15  l=0.13u w=0.32u m=1
M4 N_8 S0 N_6 GND mn15  l=0.13u w=0.32u m=1
M5 N_8 B GND GND mn15  l=0.13u w=0.18u m=1
M6 N_7 N_3 N_6 GND mn15  l=0.13u w=0.32u m=1
M7 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_3 S0 VDD VDD mp15  l=0.13u w=0.46u m=1
M11 N_6 S0 N_7 VDD mp15  l=0.13u w=0.5u m=1
M12 N_8 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_8 N_3 N_6 VDD mp15  l=0.13u w=0.5u m=1
.ends ckmx02d2
* SPICE INPUT		Tue Jul 31 19:07:19 2018	ckmx02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckmx02d4
.subckt ckmx02d4 GND Y A B S0 VDD
M1 N_5 S0 N_4 GND mn15  l=0.13u w=0.45u m=1
M2 N_3 S0 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_5 B GND GND mn15  l=0.13u w=0.155u m=1
M4 GND B N_5 GND mn15  l=0.13u w=0.155u m=1
M5 N_5 B GND GND mn15  l=0.13u w=0.15u m=1
M6 N_9 N_3 N_4 GND mn15  l=0.13u w=0.45u m=1
M7 GND A N_9 GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.3u m=1
M10 Y N_4 GND GND mn15  l=0.13u w=0.29u m=1
M11 VDD S0 N_3 VDD mp15  l=0.13u w=0.42u m=1
M12 N_9 S0 N_4 VDD mp15  l=0.13u w=0.67u m=1
M13 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_5 N_3 N_4 VDD mp15  l=0.13u w=0.64u m=1
M16 N_9 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_9 VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckmx02d4
* SPICE INPUT		Tue Jul 31 19:07:31 2018	cknd02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknd02d0
.subckt cknd02d0 Y VDD A GND B
M1 GND A N_14 GND mn15  l=0.13u w=0.27u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.27u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.6u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.6u m=1
.ends cknd02d0
* SPICE INPUT		Tue Jul 31 19:07:43 2018	cknd02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknd02d1
.subckt cknd02d1 Y VDD A B GND
M1 GND A N_9 GND mn15  l=0.13u w=0.36u m=1
M2 Y B N_9 GND mn15  l=0.13u w=0.36u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
.ends cknd02d1
* SPICE INPUT		Tue Jul 31 19:07:56 2018	cknd02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknd02d2
.subckt cknd02d2 GND Y VDD A B
M1 N_6 A GND GND mn15  l=0.13u w=0.43u m=1
M2 N_6 B Y GND mn15  l=0.13u w=0.43u m=1
M3 Y B N_5 GND mn15  l=0.13u w=0.42u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.42u m=1
M5 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends cknd02d2
* SPICE INPUT		Tue Jul 31 19:08:08 2018	cknd02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknd02d4
.subckt cknd02d4 Y GND A B VDD
M1 Y B N_7 GND mn15  l=0.13u w=0.4u m=1
M2 GND A N_7 GND mn15  l=0.13u w=0.4u m=1
M3 N_10 A GND GND mn15  l=0.13u w=0.4u m=1
M4 N_10 B Y GND mn15  l=0.13u w=0.4u m=1
M5 Y B N_9 GND mn15  l=0.13u w=0.4u m=1
M6 N_8 A GND GND mn15  l=0.13u w=0.4u m=1
M7 N_9 A GND GND mn15  l=0.13u w=0.4u m=1
M8 N_8 B Y GND mn15  l=0.13u w=0.4u m=1
M9 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
.ends cknd02d4
* SPICE INPUT		Tue Jul 31 19:08:21 2018	cknr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknr02d0
.subckt cknr02d0 GND Y VDD B A
M1 GND A Y GND mn15  l=0.13u w=0.18u m=1
M2 Y B GND GND mn15  l=0.13u w=0.18u m=1
M3 N_10 A VDD VDD mp15  l=0.13u w=0.6u m=1
M4 N_11 A VDD VDD mp15  l=0.13u w=0.6u m=1
M5 Y B N_10 VDD mp15  l=0.13u w=0.6u m=1
M6 Y B N_11 VDD mp15  l=0.13u w=0.6u m=1
.ends cknr02d0
* SPICE INPUT		Tue Jul 31 19:08:36 2018	cknr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknr02d1
.subckt cknr02d1 GND Y VDD B A
M1 Y B GND GND mn15  l=0.13u w=0.23u m=1
M2 GND A Y GND mn15  l=0.13u w=0.23u m=1
M3 N_10 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 Y B N_10 VDD mp15  l=0.13u w=0.69u m=1
M5 Y B N_11 VDD mp15  l=0.13u w=0.69u m=1
M6 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends cknr02d1
* SPICE INPUT		Tue Jul 31 19:08:51 2018	cknr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknr02d2
.subckt cknr02d2 Y GND VDD B A
M1 GND B Y GND mn15  l=0.13u w=0.4u m=1
M2 GND A Y GND mn15  l=0.13u w=0.4u m=1
M3 N_9 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 N_10 B Y VDD mp15  l=0.13u w=0.69u m=1
M5 Y B N_9 VDD mp15  l=0.13u w=0.69u m=1
M6 VDD A N_8 VDD mp15  l=0.13u w=0.69u m=1
M7 N_10 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y B N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends cknr02d2
* SPICE INPUT		Tue Jul 31 19:09:04 2018	cknr02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknr02d4
.subckt cknr02d4 Y GND VDD A B
M1 GND A Y GND mn15  l=0.13u w=0.3u m=1
M2 GND A Y GND mn15  l=0.13u w=0.3u m=1
M3 GND B Y GND mn15  l=0.13u w=0.3u m=1
M4 GND B Y GND mn15  l=0.13u w=0.3u m=1
M5 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 N_17 B Y VDD mp15  l=0.13u w=0.69u m=1
M7 Y B N_16 VDD mp15  l=0.13u w=0.69u m=1
M8 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y B N_15 VDD mp15  l=0.13u w=0.69u m=1
M11 Y B N_18 VDD mp15  l=0.13u w=0.69u m=1
M12 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends cknr02d4
* SPICE INPUT		Tue Jul 31 19:09:21 2018	ckor02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckor02d0
.subckt ckor02d0 GND Y B VDD A
M1 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.26u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M5 N_19 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M6 N_19 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckor02d0
* SPICE INPUT		Tue Jul 31 19:09:34 2018	ckor02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckor02d1
.subckt ckor02d1 GND Y VDD A B
M1 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M3 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_13 A VDD VDD mp15  l=0.13u w=0.68u m=1
M5 N_13 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M6 N_3 B N_12 VDD mp15  l=0.13u w=0.68u m=1
M7 N_12 A VDD VDD mp15  l=0.13u w=0.68u m=1
M8 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckor02d1
* SPICE INPUT		Tue Jul 31 19:09:45 2018	ckor02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckor02d2
.subckt ckor02d2 GND Y VDD A B
M1 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M7 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_43 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M10 N_3 B N_42 VDD mp15  l=0.13u w=0.68u m=1
M11 N_43 A VDD VDD mp15  l=0.13u w=0.68u m=1
M12 N_40 A VDD VDD mp15  l=0.13u w=0.68u m=1
M13 N_41 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M14 N_3 B N_40 VDD mp15  l=0.13u w=0.68u m=1
M15 N_42 A VDD VDD mp15  l=0.13u w=0.68u m=1
M16 VDD A N_41 VDD mp15  l=0.13u w=0.68u m=1
.ends ckor02d2
* SPICE INPUT		Tue Jul 31 19:09:57 2018	ckor02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckor02d4
.subckt ckor02d4 GND Y A B VDD
M1 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND B N_3 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_60 A VDD VDD mp15  l=0.13u w=0.68u m=1
M12 N_61 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M13 N_3 B N_60 VDD mp15  l=0.13u w=0.68u m=1
M14 N_62 A VDD VDD mp15  l=0.13u w=0.68u m=1
M15 VDD A N_61 VDD mp15  l=0.13u w=0.68u m=1
M16 N_63 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M17 N_3 B N_62 VDD mp15  l=0.13u w=0.68u m=1
M18 N_64 A VDD VDD mp15  l=0.13u w=0.68u m=1
M19 VDD A N_63 VDD mp15  l=0.13u w=0.68u m=1
M20 N_65 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M21 N_3 B N_64 VDD mp15  l=0.13u w=0.68u m=1
M22 N_65 A VDD VDD mp15  l=0.13u w=0.68u m=1
M23 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckor02d4
* SPICE INPUT		Tue Jul 31 19:10:09 2018	ckxn02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxn02d0
.subckt ckxn02d0 GND Y VDD A B
M1 GND B N_2 GND mn15  l=0.13u w=0.2u m=1
M2 N_9 N_2 GND GND mn15  l=0.13u w=0.2u m=1
M3 N_9 N_8 N_3 GND mn15  l=0.13u w=0.2u m=1
M4 N_3 A N_2 GND mn15  l=0.13u w=0.2u m=1
M5 GND N_3 Y GND mn15  l=0.13u w=0.2u m=1
M6 N_8 A GND GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M8 N_16 N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_16 A N_3 VDD mp15  l=0.13u w=0.69u m=1
M10 N_2 N_8 N_3 VDD mp15  l=0.13u w=0.345u m=1
M11 N_2 N_8 N_3 VDD mp15  l=0.13u w=0.345u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckxn02d0
* SPICE INPUT		Tue Jul 31 19:10:20 2018	ckxn02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxn02d1
.subckt ckxn02d1 GND Y VDD A B
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_6 GND GND mn15  l=0.13u w=0.4u m=1
M3 N_6 A N_5 GND mn15  l=0.13u w=0.2u m=1
M4 GND B N_5 GND mn15  l=0.13u w=0.2u m=1
M5 N_9 N_5 GND GND mn15  l=0.13u w=0.2u m=1
M6 N_9 N_4 N_6 GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_38 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_38 A N_6 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.35u m=1
M11 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.34u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.59u m=1
M14 VDD N_6 Y VDD mp15  l=0.13u w=0.59u m=1
.ends ckxn02d1
* SPICE INPUT		Tue Jul 31 19:10:32 2018	ckxn02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxn02d2
.subckt ckxn02d2 GND Y VDD A B
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_6 A N_5 GND mn15  l=0.13u w=0.2u m=1
M4 GND B N_5 GND mn15  l=0.13u w=0.2u m=1
M5 N_9 N_5 GND GND mn15  l=0.13u w=0.2u m=1
M6 N_9 N_4 N_6 GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_38 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_38 A N_6 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.35u m=1
M11 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.34u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckxn02d2
* SPICE INPUT		Tue Jul 31 19:10:44 2018	ckxn02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxn02d4
.subckt ckxn02d4 GND Y VDD B A
M1 N_3 N_6 N_2 GND mn15  l=0.13u w=0.39u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.18u m=1
M3 N_2 N_8 GND GND mn15  l=0.13u w=0.39u m=1
M4 N_8 A N_3 GND mn15  l=0.13u w=0.39u m=1
M5 N_8 B GND GND mn15  l=0.13u w=0.39u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.355u m=1
M7 Y N_3 GND GND mn15  l=0.13u w=0.355u m=1
M8 Y N_3 GND GND mn15  l=0.13u w=0.35u m=1
M9 N_8 N_6 N_3 VDD mp15  l=0.13u w=0.59u m=1
M10 N_3 N_6 N_8 VDD mp15  l=0.13u w=0.59u m=1
M11 N_20 A N_3 VDD mp15  l=0.13u w=0.59u m=1
M12 N_3 A N_19 VDD mp15  l=0.13u w=0.59u m=1
M13 N_6 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_8 B VDD VDD mp15  l=0.13u w=0.59u m=1
M15 N_8 B VDD VDD mp15  l=0.13u w=0.59u m=1
M16 N_19 N_8 VDD VDD mp15  l=0.13u w=0.59u m=1
M17 N_20 N_8 VDD VDD mp15  l=0.13u w=0.59u m=1
M18 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M21 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckxn02d4
* SPICE INPUT		Tue Jul 31 19:10:57 2018	ckxr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxr02d0
.subckt ckxr02d0 GND Y A VDD B
M1 GND B N_2 GND mn15  l=0.13u w=0.2u m=1
M2 N_9 N_2 GND GND mn15  l=0.13u w=0.2u m=1
M3 N_3 N_8 N_2 GND mn15  l=0.13u w=0.2u m=1
M4 N_9 A N_3 GND mn15  l=0.13u w=0.2u m=1
M5 N_8 A GND GND mn15  l=0.13u w=0.2u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M8 N_37 N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_37 N_8 N_3 VDD mp15  l=0.13u w=0.69u m=1
M10 N_2 A N_3 VDD mp15  l=0.13u w=0.345u m=1
M11 N_3 A N_2 VDD mp15  l=0.13u w=0.345u m=1
M12 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckxr02d0
* SPICE INPUT		Tue Jul 31 19:11:08 2018	ckxr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxr02d1
.subckt ckxr02d1 GND Y A VDD B
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_8 GND GND mn15  l=0.13u w=0.4u m=1
M3 GND B N_5 GND mn15  l=0.13u w=0.2u m=1
M4 N_9 N_5 GND GND mn15  l=0.13u w=0.2u m=1
M5 N_8 N_4 N_5 GND mn15  l=0.13u w=0.2u m=1
M6 N_8 A N_9 GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_16 N_4 N_8 VDD mp15  l=0.13u w=0.69u m=1
M9 N_16 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_8 A N_5 VDD mp15  l=0.13u w=0.345u m=1
M11 N_5 A N_8 VDD mp15  l=0.13u w=0.345u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_8 Y VDD mp15  l=0.13u w=0.61u m=1
M14 VDD N_8 Y VDD mp15  l=0.13u w=0.61u m=1
.ends ckxr02d1
* SPICE INPUT		Tue Jul 31 19:11:22 2018	ckxr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxr02d2
.subckt ckxr02d2 GND Y A VDD B
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_5 GND mn15  l=0.13u w=0.2u m=1
M4 N_9 N_5 GND GND mn15  l=0.13u w=0.2u m=1
M5 N_8 N_4 N_5 GND mn15  l=0.13u w=0.2u m=1
M6 N_8 A N_9 GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_16 N_4 N_8 VDD mp15  l=0.13u w=0.69u m=1
M9 N_16 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_8 A N_5 VDD mp15  l=0.13u w=0.345u m=1
M11 N_5 A N_8 VDD mp15  l=0.13u w=0.345u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckxr02d2
* SPICE INPUT		Tue Jul 31 19:11:37 2018	ckxr02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxr02d4
.subckt ckxr02d4 GND Y VDD A B
M1 N_3 B GND GND mn15  l=0.13u w=0.39u m=1
M2 N_11 N_3 GND GND mn15  l=0.13u w=0.39u m=1
M3 N_11 A N_2 GND mn15  l=0.13u w=0.39u m=1
M4 N_3 N_8 N_2 GND mn15  l=0.13u w=0.39u m=1
M5 GND A N_8 GND mn15  l=0.13u w=0.19u m=1
M6 Y N_2 GND GND mn15  l=0.13u w=0.355u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.355u m=1
M8 Y N_2 GND GND mn15  l=0.13u w=0.35u m=1
M9 VDD B N_3 VDD mp15  l=0.13u w=0.59u m=1
M10 N_3 B VDD VDD mp15  l=0.13u w=0.59u m=1
M11 N_16 N_3 VDD VDD mp15  l=0.13u w=0.59u m=1
M12 VDD N_3 N_16 VDD mp15  l=0.13u w=0.59u m=1
M13 N_16 N_8 N_2 VDD mp15  l=0.13u w=0.59u m=1
M14 N_16 N_8 N_2 VDD mp15  l=0.13u w=0.59u m=1
M15 N_2 A N_3 VDD mp15  l=0.13u w=1.18u m=1
M16 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckxr02d4

* SPICE INPUT		Tue Jul 31 19:23:44 2018	dl01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d1
.subckt dl01d1 VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.14u m=1
M2 GND N_4 N_3 GND mn15  l=0.13u w=0.14u m=1
M3 N_7 N_3 GND GND mn15  l=0.13u w=0.14u m=1
M4 GND N_7 Y GND mn15  l=0.13u w=0.2u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.49u m=1
M6 N_3 N_4 VDD VDD mp15  l=0.13u w=0.49u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.13u w=0.49u m=1
M8 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends dl01d1
* SPICE INPUT		Tue Jul 31 19:23:56 2018	dl01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d2
.subckt dl01d2 Y VDD GND A
M1 N_8 A GND GND mn15  l=0.13u w=0.14u m=1
M2 GND N_8 N_7 GND mn15  l=0.13u w=0.14u m=1
M3 GND N_7 N_4 GND mn15  l=0.13u w=0.14u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.24u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.24u m=1
M6 VDD N_7 N_4 VDD mp15  l=0.13u w=0.49u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_8 A VDD VDD mp15  l=0.13u w=0.49u m=1
M10 N_7 N_8 VDD VDD mp15  l=0.13u w=0.49u m=1
.ends dl01d2
* SPICE INPUT		Tue Jul 31 19:24:09 2018	dl01dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01dm
.subckt dl01dm VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.14u m=1
M2 GND N_4 N_3 GND mn15  l=0.13u w=0.14u m=1
M3 N_7 N_3 GND GND mn15  l=0.13u w=0.14u m=1
M4 GND N_7 Y GND mn15  l=0.13u w=0.18u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.49u m=1
M6 N_3 N_4 VDD VDD mp15  l=0.13u w=0.49u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.13u w=0.49u m=1
M8 Y N_7 VDD VDD mp15  l=0.13u w=0.63u m=1
.ends dl01dm
* SPICE INPUT		Tue Jul 31 19:24:22 2018	dl02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d1
.subckt dl02d1 VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.14u m=1
M2 GND N_4 N_3 GND mn15  l=0.26u w=0.14u m=1
M3 N_7 N_3 GND GND mn15  l=0.26u w=0.14u m=1
M4 GND N_7 Y GND mn15  l=0.13u w=0.2u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.49u m=1
M6 N_3 N_4 VDD VDD mp15  l=0.26u w=0.49u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.26u w=0.49u m=1
M8 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends dl02d1
* SPICE INPUT		Tue Jul 31 19:24:35 2018	dl02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d2
.subckt dl02d2 VDD Y GND A
M1 GND N_3 N_7 GND mn15  l=0.26u w=0.14u m=1
M2 GND N_7 Y GND mn15  l=0.13u w=0.34u m=1
M3 GND N_7 Y GND mn15  l=0.13u w=0.14u m=1
M4 N_4 A GND GND mn15  l=0.13u w=0.14u m=1
M5 GND N_4 N_3 GND mn15  l=0.26u w=0.14u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.49u m=1
M7 N_3 N_4 VDD VDD mp15  l=0.26u w=0.49u m=1
M8 VDD N_3 N_7 VDD mp15  l=0.26u w=0.49u m=1
M9 VDD N_7 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_7 Y VDD mp15  l=0.13u w=0.69u m=1
.ends dl02d2
* SPICE INPUT		Tue Jul 31 19:24:48 2018	dmnrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dmnrq0
.subckt dmnrq0 GND Q VDD CK D1 S0 D0
M1 GND S0 N_4 GND mn15  l=0.13u w=0.18u m=1
M2 N_18 D0 GND GND mn15  l=0.13u w=0.18u m=1
M3 N_18 N_4 N_6 GND mn15  l=0.13u w=0.18u m=1
M4 N_19 S0 N_6 GND mn15  l=0.13u w=0.18u m=1
M5 N_19 D1 GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.17u m=1
M7 N_20 N_12 N_9 GND mn15  l=0.13u w=0.17u m=1
M8 N_20 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M9 GND N_9 N_7 GND mn15  l=0.13u w=0.18u m=1
M10 N_6 N_2 N_9 GND mn15  l=0.13u w=0.28u m=1
M11 GND N_2 N_12 GND mn15  l=0.13u w=0.17u m=1
M12 N_22 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M13 N_22 N_12 N_14 GND mn15  l=0.13u w=0.17u m=1
M14 N_14 N_2 N_21 GND mn15  l=0.13u w=0.17u m=1
M15 N_21 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M16 Q N_14 GND GND mn15  l=0.13u w=0.26u m=1
M17 N_17 N_14 GND GND mn15  l=0.13u w=0.18u m=1
M18 N_4 S0 VDD VDD mp15  l=0.13u w=0.26u m=1
M19 N_39 D0 VDD VDD mp15  l=0.13u w=0.28u m=1
M20 N_39 S0 N_6 VDD mp15  l=0.13u w=0.28u m=1
M21 N_40 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M22 N_40 D1 VDD VDD mp15  l=0.13u w=0.28u m=1
M23 N_2 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M24 N_6 N_12 N_9 VDD mp15  l=0.13u w=0.42u m=1
M25 N_41 N_7 VDD VDD mp15  l=0.13u w=0.17u m=1
M26 VDD N_9 N_7 VDD mp15  l=0.13u w=0.26u m=1
M27 N_41 N_2 N_9 VDD mp15  l=0.13u w=0.17u m=1
M28 N_12 N_2 VDD VDD mp15  l=0.13u w=0.42u m=1
M29 N_43 N_7 VDD VDD mp15  l=0.13u w=0.27u m=1
M30 N_14 N_12 N_42 VDD mp15  l=0.13u w=0.17u m=1
M31 N_14 N_2 N_43 VDD mp15  l=0.13u w=0.27u m=1
M32 N_42 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M33 VDD N_14 Q VDD mp15  l=0.13u w=0.4u m=1
M34 N_17 N_14 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends dmnrq0
* SPICE INPUT		Tue Jul 31 19:25:01 2018	dmnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dmnrq1
.subckt dmnrq1 GND Q VDD CK D1 S0 D0
M1 N_5 N_6 N_18 GND mn15  l=0.13u w=0.17u m=1
M2 N_19 N_3 N_5 GND mn15  l=0.13u w=0.36u m=1
M3 GND N_6 N_3 GND mn15  l=0.13u w=0.2u m=1
M4 N_18 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_19 N_15 GND GND mn15  l=0.13u w=0.36u m=1
M6 GND S0 N_8 GND mn15  l=0.13u w=0.17u m=1
M7 N_20 D0 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_20 N_8 N_10 GND mn15  l=0.13u w=0.28u m=1
M9 N_21 S0 N_10 GND mn15  l=0.13u w=0.28u m=1
M10 N_21 D1 GND GND mn15  l=0.13u w=0.28u m=1
M11 GND CK N_6 GND mn15  l=0.13u w=0.2u m=1
M12 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_13 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M14 N_10 N_6 N_16 GND mn15  l=0.13u w=0.28u m=1
M15 N_15 N_16 GND GND mn15  l=0.13u w=0.28u m=1
M16 N_22 N_3 N_16 GND mn15  l=0.13u w=0.17u m=1
M17 N_22 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M18 VDD S0 N_8 VDD mp15  l=0.13u w=0.24u m=1
M19 N_39 D0 VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_10 S0 N_39 VDD mp15  l=0.13u w=0.42u m=1
M21 N_40 N_8 N_10 VDD mp15  l=0.13u w=0.42u m=1
M22 N_40 D1 VDD VDD mp15  l=0.13u w=0.42u m=1
M23 N_6 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M24 N_41 N_6 N_16 VDD mp15  l=0.13u w=0.17u m=1
M25 VDD N_16 N_15 VDD mp15  l=0.13u w=0.42u m=1
M26 N_10 N_3 N_16 VDD mp15  l=0.13u w=0.42u m=1
M27 N_41 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 N_43 N_6 N_5 VDD mp15  l=0.13u w=0.52u m=1
M29 N_5 N_3 N_42 VDD mp15  l=0.13u w=0.17u m=1
M30 N_3 N_6 VDD VDD mp15  l=0.13u w=0.51u m=1
M31 N_42 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_43 N_15 VDD VDD mp15  l=0.13u w=0.52u m=1
M33 VDD N_5 Q VDD mp15  l=0.13u w=0.69u m=1
M34 N_13 N_5 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends dmnrq1
* SPICE INPUT		Tue Jul 31 19:25:14 2018	dmnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dmnrq2
.subckt dmnrq2 GND Q VDD CK D1 S0 D0
M1 GND S0 N_4 GND mn15  l=0.13u w=0.24u m=1
M2 N_19 D0 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_6 N_4 N_19 GND mn15  l=0.13u w=0.28u m=1
M4 N_20 S0 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_20 D1 GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 CK GND GND mn15  l=0.13u w=0.28u m=1
M7 N_21 N_18 GND GND mn15  l=0.13u w=0.41u m=1
M8 N_21 N_13 N_10 GND mn15  l=0.13u w=0.41u m=1
M9 N_22 N_3 N_10 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_8 N_22 GND mn15  l=0.13u w=0.17u m=1
M11 Q N_10 GND GND mn15  l=0.13u w=0.46u m=1
M12 Q N_10 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_8 N_10 GND GND mn15  l=0.13u w=0.37u m=1
M14 N_23 N_13 N_16 GND mn15  l=0.13u w=0.17u m=1
M15 N_16 N_3 N_6 GND mn15  l=0.13u w=0.41u m=1
M16 GND N_18 N_23 GND mn15  l=0.13u w=0.17u m=1
M17 N_18 N_16 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_18 N_16 GND GND mn15  l=0.13u w=0.15u m=1
M19 GND N_3 N_13 GND mn15  l=0.13u w=0.23u m=1
M20 VDD S0 N_4 VDD mp15  l=0.13u w=0.37u m=1
M21 N_41 D0 VDD VDD mp15  l=0.13u w=0.42u m=1
M22 N_6 S0 N_41 VDD mp15  l=0.13u w=0.42u m=1
M23 N_42 N_4 N_6 VDD mp15  l=0.13u w=0.42u m=1
M24 N_42 D1 VDD VDD mp15  l=0.13u w=0.42u m=1
M25 N_3 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M26 N_16 N_13 N_6 VDD mp15  l=0.13u w=0.63u m=1
M27 N_43 N_3 N_16 VDD mp15  l=0.13u w=0.17u m=1
M28 N_43 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 VDD N_16 N_18 VDD mp15  l=0.13u w=0.63u m=1
M30 VDD N_3 N_13 VDD mp15  l=0.13u w=0.57u m=1
M31 N_44 N_18 VDD VDD mp15  l=0.13u w=0.62u m=1
M32 N_44 N_3 N_10 VDD mp15  l=0.13u w=0.62u m=1
M33 N_45 N_13 N_10 VDD mp15  l=0.13u w=0.17u m=1
M34 VDD N_8 N_45 VDD mp15  l=0.13u w=0.17u m=1
M35 N_8 N_10 VDD VDD mp15  l=0.13u w=0.55u m=1
M36 Q N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M37 Q N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends dmnrq2
* SPICE INPUT		Tue Jul 31 19:26:49 2018	fillercap16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap16
.subckt fillercap16 GND VDD
M1 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M2 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M3 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M4 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
.ends fillercap16
* SPICE INPUT		Tue Jul 31 19:27:11 2018	fillercap3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap3
.subckt fillercap3 VDD GND
M1 VDD GND VDD VDD mp15  l=0.33u w=0.69u m=1
.ends fillercap3
* SPICE INPUT		Tue Jul 31 19:27:24 2018	fillercap32
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap32
.subckt fillercap32 GND VDD
M1 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M2 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M3 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M4 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M5 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M6 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M7 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M8 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M9 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M10 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
.ends fillercap32
* SPICE INPUT		Tue Jul 31 19:27:37 2018	fillercap4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap4
.subckt fillercap4 VDD GND
M1 VDD GND VDD VDD mp15  l=0.67u w=0.69u m=1
.ends fillercap4
* SPICE INPUT		Tue Jul 31 19:27:50 2018	fillercap6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap6
.subckt fillercap6 VDD GND
M1 VDD GND VDD VDD mp15  l=0.33u w=1.22u m=1
.ends fillercap6
* SPICE INPUT		Tue Jul 31 19:28:03 2018	fillercap64
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap64
.subckt fillercap64 GND VDD
M1 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M2 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M3 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M4 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M5 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M6 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M7 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M8 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M9 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M10 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M11 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M12 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M13 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M14 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M15 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M16 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M17 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M18 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M19 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M20 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M21 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M22 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
.ends fillercap64
* SPICE INPUT		Tue Jul 31 19:28:16 2018	fillercap8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap8
.subckt fillercap8 VDD GND
M1 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
.ends fillercap8
* SPICE INPUT		Tue Jul 31 19:28:38 2018	inv0d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d0
.subckt inv0d0 GND VDD Y A
M1 Y A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends inv0d0
* SPICE INPUT		Tue Jul 31 19:28:51 2018	inv0d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d1
.subckt inv0d1 GND VDD Y A
M1 Y A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d1
* SPICE INPUT		Tue Jul 31 19:29:04 2018	inv0d12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d12
.subckt inv0d12 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A Y GND mn15  l=0.13u w=0.46u m=1
M8 Y A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND A Y GND mn15  l=0.13u w=0.46u m=1
M10 Y A GND GND mn15  l=0.13u w=0.46u m=1
M11 GND A Y GND mn15  l=0.13u w=0.46u m=1
M12 Y A GND GND mn15  l=0.13u w=0.46u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d12
* SPICE INPUT		Tue Jul 31 19:29:17 2018	inv0d16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d16
.subckt inv0d16 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A Y GND mn15  l=0.13u w=0.46u m=1
M8 Y A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND A Y GND mn15  l=0.13u w=0.46u m=1
M10 Y A GND GND mn15  l=0.13u w=0.46u m=1
M11 GND A Y GND mn15  l=0.13u w=0.46u m=1
M12 Y A GND GND mn15  l=0.13u w=0.46u m=1
M13 GND A Y GND mn15  l=0.13u w=0.46u m=1
M14 Y A GND GND mn15  l=0.13u w=0.46u m=1
M15 GND A Y GND mn15  l=0.13u w=0.46u m=1
M16 Y A GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M31 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d16
* SPICE INPUT		Tue Jul 31 19:29:30 2018	inv0d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d2
.subckt inv0d2 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M4 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d2
* SPICE INPUT		Tue Jul 31 19:29:42 2018	inv0d20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d20
.subckt inv0d20 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A Y GND mn15  l=0.13u w=0.46u m=1
M8 Y A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND A Y GND mn15  l=0.13u w=0.46u m=1
M10 Y A GND GND mn15  l=0.13u w=0.46u m=1
M11 GND A Y GND mn15  l=0.13u w=0.46u m=1
M12 Y A GND GND mn15  l=0.13u w=0.46u m=1
M13 GND A Y GND mn15  l=0.13u w=0.46u m=1
M14 Y A GND GND mn15  l=0.13u w=0.46u m=1
M15 GND A Y GND mn15  l=0.13u w=0.46u m=1
M16 Y A GND GND mn15  l=0.13u w=0.46u m=1
M17 GND A Y GND mn15  l=0.13u w=0.46u m=1
M18 Y A GND GND mn15  l=0.13u w=0.46u m=1
M19 GND A Y GND mn15  l=0.13u w=0.46u m=1
M20 Y A GND GND mn15  l=0.13u w=0.46u m=1
M21 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M31 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M33 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M34 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M35 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M36 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M37 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M38 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M39 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M40 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d20
* SPICE INPUT		Tue Jul 31 19:29:55 2018	inv0d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d3
.subckt inv0d3 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y A GND GND mn15  l=0.13u w=0.46u m=1
M4 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M5 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d3
* SPICE INPUT		Tue Jul 31 19:30:08 2018	inv0d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d4
.subckt inv0d4 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M6 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d4
* SPICE INPUT		Tue Jul 31 19:30:21 2018	inv0d5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d5
.subckt inv0d5 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A Y GND mn15  l=0.13u w=0.46u m=1
M5 Y A GND GND mn15  l=0.13u w=0.46u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d5
* SPICE INPUT		Tue Jul 31 19:30:34 2018	inv0d6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d6
.subckt inv0d6 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d6
* SPICE INPUT		Tue Jul 31 19:30:47 2018	inv0d7
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d7
.subckt inv0d7 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A Y GND mn15  l=0.13u w=0.46u m=1
M5 Y A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A Y GND mn15  l=0.13u w=0.46u m=1
M7 Y A GND GND mn15  l=0.13u w=0.46u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d7
* SPICE INPUT		Tue Jul 31 19:31:00 2018	inv0d8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d8
.subckt inv0d8 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A Y GND mn15  l=0.13u w=0.46u m=1
M8 Y A GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d8
* SPICE INPUT		Tue Jul 31 19:31:13 2018	inv0dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0dm
.subckt inv0dm GND VDD Y A
M1 Y A GND GND mn15  l=0.13u w=0.36u m=1
M2 Y A VDD VDD mp15  l=0.13u w=0.55u m=1
.ends inv0dm
* SPICE INPUT		Tue Jul 31 19:31:26 2018	inv0dp
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0dp
.subckt inv0dp Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.355u m=1
M2 GND A Y GND mn15  l=0.13u w=0.355u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
M4 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
.ends inv0dp
* SPICE INPUT		Tue Jul 31 19:31:40 2018	invod8d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invod8d1
.subckt invod8d1 GND Y0 Y6 Y5 Y2 Y1 Y7 Y4 Y3 VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y0 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 Y5 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 Y1 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y2 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y7 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M8 Y4 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y3 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M10 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
.ends invod8d1
* SPICE INPUT		Tue Jul 31 19:31:52 2018	invtld0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld0
.subckt invtld0 GND Y VDD A E
M1 GND E N_3 GND mn15  l=0.13u w=0.26u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y E N_6 GND mn15  l=0.13u w=0.26u m=1
M4 Y E N_7 GND mn15  l=0.13u w=0.26u m=1
M5 GND A N_6 GND mn15  l=0.13u w=0.26u m=1
M6 VDD E N_3 VDD mp15  l=0.13u w=0.4u m=1
M7 N_14 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 Y N_3 N_13 VDD mp15  l=0.13u w=0.4u m=1
M9 Y N_3 N_14 VDD mp15  l=0.13u w=0.4u m=1
M10 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends invtld0
* SPICE INPUT		Tue Jul 31 19:32:06 2018	invtld1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld1
.subckt invtld1 Y VDD GND A E
M1 GND E N_3 GND mn15  l=0.13u w=0.31u m=1
M2 GND A N_13 GND mn15  l=0.13u w=0.46u m=1
M3 Y E N_15 GND mn15  l=0.13u w=0.46u m=1
M4 Y E N_13 GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_15 GND mn15  l=0.13u w=0.46u m=1
M6 VDD E N_3 VDD mp15  l=0.13u w=0.46u m=1
M7 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_7 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M9 Y N_3 N_8 VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends invtld1
* SPICE INPUT		Tue Jul 31 19:32:19 2018	invtld12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld12
.subckt invtld12 GND Y VDD E A
M1 GND E N_2 GND mn15  l=0.13u w=0.42u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.31u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.31u m=1
M4 N_7 N_5 GND GND mn15  l=0.13u w=0.455u m=1
M5 N_7 N_5 GND GND mn15  l=0.13u w=0.45u m=1
M6 N_7 N_5 GND GND mn15  l=0.13u w=0.45u m=1
M7 N_7 N_5 GND GND mn15  l=0.13u w=0.45u m=1
M8 N_7 N_5 GND GND mn15  l=0.13u w=0.415u m=1
M9 N_6 E N_7 GND mn15  l=0.13u w=0.4u m=1
M10 N_6 E N_7 GND mn15  l=0.13u w=0.405u m=1
M11 N_7 E N_6 GND mn15  l=0.13u w=0.395u m=1
M12 GND N_2 N_7 GND mn15  l=0.13u w=0.37u m=1
M13 N_7 N_2 GND GND mn15  l=0.13u w=0.37u m=1
M14 N_7 N_2 GND GND mn15  l=0.13u w=0.37u m=1
M15 Y N_7 GND GND mn15  l=0.13u w=0.43u m=1
M16 GND N_7 Y GND mn15  l=0.13u w=0.4u m=1
M17 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M18 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M19 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M20 GND N_7 Y GND mn15  l=0.13u w=0.42u m=1
M21 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M22 GND N_7 Y GND mn15  l=0.13u w=0.42u m=1
M23 Y N_7 GND GND mn15  l=0.13u w=0.4u m=1
M24 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M25 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M26 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M27 Y N_7 GND GND mn15  l=0.13u w=0.37u m=1
M28 N_2 E VDD VDD mp15  l=0.13u w=0.63u m=1
M29 N_5 A VDD VDD mp15  l=0.13u w=0.47u m=1
M30 N_5 A VDD VDD mp15  l=0.13u w=0.47u m=1
M31 VDD N_6 Y VDD mp15  l=0.13u w=0.72u m=1
M32 VDD N_6 Y VDD mp15  l=0.13u w=0.72u m=1
M33 Y N_6 VDD VDD mp15  l=0.13u w=0.72u m=1
M34 VDD N_6 Y VDD mp15  l=0.13u w=0.72u m=1
M35 Y N_6 VDD VDD mp15  l=0.13u w=0.72u m=1
M36 VDD N_6 Y VDD mp15  l=0.13u w=0.71u m=1
M37 VDD N_6 Y VDD mp15  l=0.13u w=0.71u m=1
M38 Y N_6 VDD VDD mp15  l=0.13u w=0.71u m=1
M39 VDD N_6 Y VDD mp15  l=0.13u w=0.68u m=1
M40 VDD N_6 Y VDD mp15  l=0.13u w=0.64u m=1
M41 VDD N_6 Y VDD mp15  l=0.13u w=0.64u m=1
M42 VDD N_6 Y VDD mp15  l=0.13u w=0.59u m=1
M43 N_6 N_5 VDD VDD mp15  l=0.13u w=0.54u m=1
M44 N_6 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M45 N_6 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M46 N_6 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M47 N_6 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M48 N_6 E VDD VDD mp15  l=0.13u w=0.57u m=1
M49 N_6 E VDD VDD mp15  l=0.13u w=0.57u m=1
M50 VDD E N_6 VDD mp15  l=0.13u w=0.48u m=1
M51 N_7 N_2 N_6 VDD mp15  l=0.13u w=0.76u m=1
M52 N_6 N_2 N_7 VDD mp15  l=0.13u w=0.78u m=1
M53 N_7 N_2 N_6 VDD mp15  l=0.13u w=0.78u m=1
.ends invtld12
* SPICE INPUT		Tue Jul 31 19:32:33 2018	invtld16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld16
.subckt invtld16 GND Y A VDD E
M1 N_3 N_16 GND GND mn15  l=0.13u w=0.37u m=1
M2 N_3 N_16 GND GND mn15  l=0.13u w=0.37u m=1
M3 GND N_16 N_3 GND mn15  l=0.13u w=0.37u m=1
M4 N_3 N_16 GND GND mn15  l=0.13u w=0.35u m=1
M5 GND N_5 N_3 GND mn15  l=0.13u w=0.41u m=1
M6 GND N_5 N_3 GND mn15  l=0.13u w=0.44u m=1
M7 GND N_5 N_3 GND mn15  l=0.13u w=0.44u m=1
M8 N_3 N_5 GND GND mn15  l=0.13u w=0.44u m=1
M9 GND N_5 N_3 GND mn15  l=0.13u w=0.44u m=1
M10 N_3 N_5 GND GND mn15  l=0.13u w=0.39u m=1
M11 N_3 N_5 GND GND mn15  l=0.13u w=0.37u m=1
M12 GND A N_5 GND mn15  l=0.13u w=0.39u m=1
M13 N_5 A GND GND mn15  l=0.13u w=0.39u m=1
M14 GND E N_16 GND mn15  l=0.13u w=0.44u m=1
M15 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M16 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M17 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M18 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M19 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M20 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M21 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M22 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M23 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M24 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M25 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M26 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M27 Y N_3 GND GND mn15  l=0.13u w=0.39u m=1
M28 GND N_3 Y GND mn15  l=0.13u w=0.39u m=1
M29 Y N_3 GND GND mn15  l=0.13u w=0.39u m=1
M30 Y N_3 GND GND mn15  l=0.13u w=0.39u m=1
M31 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M32 N_37 E N_3 GND mn15  l=0.13u w=0.55u m=1
M33 N_3 E N_37 GND mn15  l=0.13u w=0.55u m=1
M34 N_3 E N_37 GND mn15  l=0.13u w=0.46u m=1
M35 N_37 E VDD VDD mp15  l=0.13u w=0.76u m=1
M36 N_37 E VDD VDD mp15  l=0.13u w=0.76u m=1
M37 VDD E N_37 VDD mp15  l=0.13u w=0.67u m=1
M38 N_16 E VDD VDD mp15  l=0.13u w=0.67u m=1
M39 N_37 N_5 VDD VDD mp15  l=0.13u w=0.63u m=1
M40 VDD N_5 N_37 VDD mp15  l=0.13u w=0.63u m=1
M41 N_37 N_5 VDD VDD mp15  l=0.13u w=0.63u m=1
M42 VDD N_5 N_37 VDD mp15  l=0.13u w=0.63u m=1
M43 N_37 N_5 VDD VDD mp15  l=0.13u w=0.63u m=1
M44 VDD N_5 N_37 VDD mp15  l=0.13u w=0.63u m=1
M45 N_37 N_5 VDD VDD mp15  l=0.13u w=0.62u m=1
M46 VDD A N_5 VDD mp15  l=0.13u w=0.59u m=1
M47 N_5 A VDD VDD mp15  l=0.13u w=0.59u m=1
M48 N_3 N_16 N_37 VDD mp15  l=0.13u w=0.54u m=1
M49 N_37 N_16 N_3 VDD mp15  l=0.13u w=0.54u m=1
M50 N_37 N_16 N_3 VDD mp15  l=0.13u w=0.54u m=1
M51 N_3 N_16 N_37 VDD mp15  l=0.13u w=0.54u m=1
M52 N_37 N_16 N_3 VDD mp15  l=0.13u w=0.54u m=1
M53 N_37 N_16 N_3 VDD mp15  l=0.13u w=0.4u m=1
M54 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M55 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M56 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M57 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M58 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M59 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M60 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M61 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M62 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M63 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M64 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M65 Y N_37 VDD VDD mp15  l=0.13u w=0.64u m=1
M66 Y N_37 VDD VDD mp15  l=0.13u w=0.61u m=1
M67 VDD N_37 Y VDD mp15  l=0.13u w=0.55u m=1
M68 Y N_37 VDD VDD mp15  l=0.13u w=0.55u m=1
M69 VDD N_37 Y VDD mp15  l=0.13u w=0.55u m=1
M70 Y N_37 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends invtld16
* SPICE INPUT		Tue Jul 31 19:32:46 2018	invtld2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld2
.subckt invtld2 GND Y VDD E A
M1 N_3 E GND GND mn15  l=0.13u w=0.46u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_5 E Y GND mn15  l=0.13u w=0.42u m=1
M7 N_5 E Y GND mn15  l=0.13u w=0.57u m=1
M8 N_5 E Y GND mn15  l=0.13u w=0.57u m=1
M9 Y E N_5 GND mn15  l=0.13u w=0.29u m=1
M10 VDD E N_3 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A N_14 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_14 VDD mp15  l=0.13u w=0.69u m=1
M13 N_14 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_14 VDD mp15  l=0.13u w=0.69u m=1
M15 Y N_3 N_14 VDD mp15  l=0.13u w=0.57u m=1
M16 Y N_3 N_14 VDD mp15  l=0.13u w=0.57u m=1
M17 Y N_3 N_14 VDD mp15  l=0.13u w=0.57u m=1
M18 N_14 N_3 Y VDD mp15  l=0.13u w=0.57u m=1
M19 Y N_3 N_14 VDD mp15  l=0.13u w=0.46u m=1
.ends invtld2
* SPICE INPUT		Tue Jul 31 19:33:00 2018	invtld20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld20
.subckt invtld20 GND Y VDD E A
M1 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M2 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_25 GND GND mn15  l=0.13u w=0.4u m=1
M4 Y N_25 GND GND mn15  l=0.13u w=0.4u m=1
M5 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M8 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_25 GND GND mn15  l=0.13u w=0.385u m=1
M10 Y N_25 GND GND mn15  l=0.13u w=0.315u m=1
M11 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M12 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M13 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M14 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M15 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M16 Y N_25 GND GND mn15  l=0.13u w=0.4u m=1
M17 Y N_25 GND GND mn15  l=0.13u w=0.4u m=1
M18 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M19 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M20 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M21 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M22 N_25 E N_24 GND mn15  l=0.13u w=0.56u m=1
M23 N_25 E N_24 GND mn15  l=0.13u w=0.56u m=1
M24 N_25 E N_24 GND mn15  l=0.13u w=0.56u m=1
M25 N_24 E N_25 GND mn15  l=0.13u w=0.27u m=1
M26 GND A N_32 GND mn15  l=0.13u w=0.46u m=1
M27 N_32 A GND GND mn15  l=0.13u w=0.46u m=1
M28 GND N_32 N_25 GND mn15  l=0.13u w=0.46u m=1
M29 N_25 N_32 GND GND mn15  l=0.13u w=0.46u m=1
M30 GND N_32 N_25 GND mn15  l=0.13u w=0.46u m=1
M31 N_25 N_32 GND GND mn15  l=0.13u w=0.46u m=1
M32 GND N_32 N_25 GND mn15  l=0.13u w=0.46u m=1
M33 N_25 N_32 GND GND mn15  l=0.13u w=0.46u m=1
M34 GND N_32 N_25 GND mn15  l=0.13u w=0.46u m=1
M35 N_25 N_32 GND GND mn15  l=0.13u w=0.46u m=1
M36 GND E N_29 GND mn15  l=0.13u w=0.46u m=1
M37 N_25 N_29 GND GND mn15  l=0.13u w=0.46u m=1
M38 N_25 N_29 GND GND mn15  l=0.13u w=0.46u m=1
M39 GND N_29 N_25 GND mn15  l=0.13u w=0.46u m=1
M40 N_25 N_29 GND GND mn15  l=0.13u w=0.46u m=1
M41 VDD A N_32 VDD mp15  l=0.13u w=0.69u m=1
M42 N_32 A VDD VDD mp15  l=0.13u w=0.69u m=1
M43 VDD N_32 N_24 VDD mp15  l=0.13u w=0.69u m=1
M44 N_24 N_32 VDD VDD mp15  l=0.13u w=0.69u m=1
M45 VDD N_32 N_24 VDD mp15  l=0.13u w=0.69u m=1
M46 N_24 N_32 VDD VDD mp15  l=0.13u w=0.69u m=1
M47 VDD N_32 N_24 VDD mp15  l=0.13u w=0.69u m=1
M48 N_24 N_32 VDD VDD mp15  l=0.13u w=0.69u m=1
M49 VDD N_32 N_24 VDD mp15  l=0.13u w=0.69u m=1
M50 N_24 N_32 VDD VDD mp15  l=0.13u w=0.69u m=1
M51 N_29 E VDD VDD mp15  l=0.13u w=0.69u m=1
M52 N_24 E VDD VDD mp15  l=0.13u w=0.69u m=1
M53 N_24 E VDD VDD mp15  l=0.13u w=0.69u m=1
M54 VDD E N_24 VDD mp15  l=0.13u w=0.69u m=1
M55 N_24 E VDD VDD mp15  l=0.13u w=0.69u m=1
M56 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.58u m=1
M57 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.58u m=1
M58 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.58u m=1
M59 N_24 N_29 N_25 VDD mp15  l=0.13u w=0.58u m=1
M60 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.58u m=1
M61 N_24 N_29 N_25 VDD mp15  l=0.13u w=0.58u m=1
M62 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.4u m=1
M63 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M64 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M65 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M66 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M67 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M68 Y N_24 VDD VDD mp15  l=0.13u w=0.665u m=1
M69 Y N_24 VDD VDD mp15  l=0.13u w=0.665u m=1
M70 VDD N_24 Y VDD mp15  l=0.13u w=0.665u m=1
M71 Y N_24 VDD VDD mp15  l=0.13u w=0.665u m=1
M72 VDD N_24 Y VDD mp15  l=0.13u w=0.65u m=1
M73 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M74 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M75 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M76 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M77 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M78 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M79 Y N_24 VDD VDD mp15  l=0.13u w=0.61u m=1
M80 VDD N_24 Y VDD mp15  l=0.13u w=0.57u m=1
M81 Y N_24 VDD VDD mp15  l=0.13u w=0.57u m=1
M82 VDD N_24 Y VDD mp15  l=0.13u w=0.57u m=1
M83 Y N_24 VDD VDD mp15  l=0.13u w=0.57u m=1
.ends invtld20
* SPICE INPUT		Tue Jul 31 19:33:13 2018	invtld3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld3
.subckt invtld3 GND Y VDD E A
M1 N_4 A GND GND mn15  l=0.13u w=0.3u m=1
M2 N_3 N_4 GND GND mn15  l=0.13u w=0.56u m=1
M3 GND N_5 N_3 GND mn15  l=0.13u w=0.28u m=1
M4 GND E N_5 GND mn15  l=0.13u w=0.3u m=1
M5 N_7 E N_3 GND mn15  l=0.13u w=0.3u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M8 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A N_4 VDD mp15  l=0.13u w=0.42u m=1
M10 VDD N_4 N_7 VDD mp15  l=0.13u w=0.42u m=1
M11 VDD N_4 N_7 VDD mp15  l=0.13u w=0.41u m=1
M12 N_3 N_5 N_7 VDD mp15  l=0.13u w=0.58u m=1
M13 VDD E N_7 VDD mp15  l=0.13u w=0.41u m=1
M14 VDD E N_5 VDD mp15  l=0.13u w=0.42u m=1
M15 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends invtld3
* SPICE INPUT		Tue Jul 31 19:33:26 2018	invtld4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld4
.subckt invtld4 Y GND E A VDD
M1 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_8 E GND GND mn15  l=0.13u w=0.3u m=1
M6 N_9 A GND GND mn15  l=0.13u w=0.34u m=1
M7 N_13 N_9 GND GND mn15  l=0.13u w=0.37u m=1
M8 N_13 N_9 GND GND mn15  l=0.13u w=0.37u m=1
M9 N_13 N_8 GND GND mn15  l=0.13u w=0.37u m=1
M10 N_13 E N_10 GND mn15  l=0.13u w=0.39u m=1
M11 N_8 E VDD VDD mp15  l=0.13u w=0.4u m=1
M12 N_9 A VDD VDD mp15  l=0.13u w=0.48u m=1
M13 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_9 N_10 VDD mp15  l=0.13u w=0.55u m=1
M18 N_10 N_9 VDD VDD mp15  l=0.13u w=0.55u m=1
M19 VDD E N_10 VDD mp15  l=0.13u w=0.55u m=1
M20 N_13 N_8 N_10 VDD mp15  l=0.13u w=0.64u m=1
.ends invtld4
* SPICE INPUT		Tue Jul 31 19:33:40 2018	invtld6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld6
.subckt invtld6 GND Y VDD E A
M1 N_4 A GND GND mn15  l=0.13u w=0.39u m=1
M2 N_3 E GND GND mn15  l=0.13u w=0.3u m=1
M3 GND N_4 N_5 GND mn15  l=0.13u w=0.37u m=1
M4 N_5 N_4 GND GND mn15  l=0.13u w=0.37u m=1
M5 N_5 N_4 GND GND mn15  l=0.13u w=0.37u m=1
M6 N_6 E N_5 GND mn15  l=0.13u w=0.59u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_5 N_3 GND GND mn15  l=0.13u w=0.55u m=1
M14 N_4 A VDD VDD mp15  l=0.13u w=0.58u m=1
M15 N_3 E VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_6 N_4 VDD VDD mp15  l=0.13u w=0.57u m=1
M17 N_6 N_4 VDD VDD mp15  l=0.13u w=0.64u m=1
M18 N_6 N_4 VDD VDD mp15  l=0.13u w=0.45u m=1
M19 N_6 E VDD VDD mp15  l=0.13u w=0.41u m=1
M20 VDD E N_6 VDD mp15  l=0.13u w=0.41u m=1
M21 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.595u m=1
M22 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.565u m=1
M23 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends invtld6
* SPICE INPUT		Tue Jul 31 19:33:52 2018	invtld8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld8
.subckt invtld8 GND Y VDD E A
M1 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 E GND GND mn15  l=0.13u w=0.39u m=1
M3 N_5 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_5 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_10 E N_5 GND mn15  l=0.13u w=0.41u m=1
M7 N_5 E N_10 GND mn15  l=0.13u w=0.38u m=1
M8 GND N_3 N_5 GND mn15  l=0.13u w=0.345u m=1
M9 GND N_3 N_5 GND mn15  l=0.13u w=0.345u m=1
M10 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M13 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M14 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M15 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M16 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M17 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M18 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD E N_3 VDD mp15  l=0.13u w=0.58u m=1
M20 N_10 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_10 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_10 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_10 E VDD VDD mp15  l=0.13u w=0.605u m=1
M24 VDD E N_10 VDD mp15  l=0.13u w=0.415u m=1
M25 N_5 N_3 N_10 VDD mp15  l=0.13u w=0.77u m=1
M26 N_5 N_3 N_10 VDD mp15  l=0.13u w=0.77u m=1
M27 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M33 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M34 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends invtld8
* SPICE INPUT		Tue Jul 31 19:34:05 2018	invtldm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtldm
.subckt invtldm VDD Y A E GND
M1 Y E N_13 GND mn15  l=0.13u w=0.47u m=1
M2 N_14 E Y GND mn15  l=0.13u w=0.24u m=1
M3 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M4 N_14 A GND GND mn15  l=0.13u w=0.24u m=1
M5 GND A N_13 GND mn15  l=0.13u w=0.47u m=1
M6 N_3 E VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_7 A VDD VDD mp15  l=0.13u w=0.55u m=1
M8 N_7 N_3 Y VDD mp15  l=0.13u w=0.55u m=1
M9 Y N_3 N_6 VDD mp15  l=0.13u w=0.55u m=1
M10 N_6 A VDD VDD mp15  l=0.13u w=0.55u m=1
.ends invtldm

* SPICE INPUT		Tue Jul 31 19:41:16 2018	mi02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d0
.subckt mi02d0 GND Y S0 VDD B A
M1 GND B N_2 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y S0 N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M5 GND S0 N_4 GND mn15  l=0.13u w=0.26u m=1
M6 VDD B N_2 VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 N_2 VDD mp15  l=0.13u w=0.4u m=1
M8 Y S0 N_6 VDD mp15  l=0.13u w=0.4u m=1
M9 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_4 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mi02d0
* SPICE INPUT		Tue Jul 31 19:41:29 2018	mi02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d1
.subckt mi02d1 GND Y S0 A B VDD
M1 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M2 Y S0 N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M4 Y N_4 N_6 GND mn15  l=0.13u w=0.46u m=1
M5 GND S0 N_4 GND mn15  l=0.13u w=0.28u m=1
M6 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M7 Y S0 N_6 VDD mp15  l=0.13u w=0.59u m=1
M8 N_6 A VDD VDD mp15  l=0.13u w=0.59u m=1
M9 Y N_4 N_2 VDD mp15  l=0.13u w=0.69u m=1
M10 N_4 S0 VDD VDD mp15  l=0.13u w=0.39u m=1
.ends mi02d1
* SPICE INPUT		Tue Jul 31 19:41:43 2018	mi02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d2
.subckt mi02d2 GND Y S0 B A VDD
M1 GND S0 N_4 GND mn15  l=0.13u w=0.37u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_7 N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_7 N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y S0 N_2 GND mn15  l=0.13u w=0.46u m=1
M9 N_2 S0 Y GND mn15  l=0.13u w=0.46u m=1
M10 N_4 S0 VDD VDD mp15  l=0.13u w=0.55u m=1
M11 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M13 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_7 S0 Y VDD mp15  l=0.13u w=0.595u m=1
M16 N_7 S0 Y VDD mp15  l=0.13u w=0.595u m=1
M17 N_2 N_4 Y VDD mp15  l=0.13u w=0.565u m=1
M18 N_2 N_4 Y VDD mp15  l=0.13u w=0.565u m=1
.ends mi02d2
* SPICE INPUT		Tue Jul 31 19:41:56 2018	mi02d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d3
.subckt mi02d3 Y GND S0 A B VDD
M1 N_3 S0 Y GND mn15  l=0.13u w=0.46u m=1
M2 N_3 S0 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_3 S0 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_14 N_6 GND mn15  l=0.13u w=0.46u m=1
M5 N_6 N_14 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_6 N_14 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M10 GND S0 N_14 GND mn15  l=0.13u w=0.45u m=1
M11 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M12 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M13 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M14 N_14 S0 VDD VDD mp15  l=0.13u w=0.67u m=1
M15 N_3 B VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_3 B VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_3 B VDD VDD mp15  l=0.13u w=0.69u m=1
M18 Y S0 N_6 VDD mp15  l=0.13u w=0.59u m=1
M19 Y S0 N_6 VDD mp15  l=0.13u w=0.57u m=1
M20 N_6 S0 Y VDD mp15  l=0.13u w=0.57u m=1
M21 Y N_14 N_3 VDD mp15  l=0.13u w=0.61u m=1
M22 N_3 N_14 Y VDD mp15  l=0.13u w=0.575u m=1
M23 N_3 N_14 Y VDD mp15  l=0.13u w=0.575u m=1
M24 N_6 A VDD VDD mp15  l=0.13u w=0.65u m=1
M25 VDD A N_6 VDD mp15  l=0.13u w=0.65u m=1
M26 VDD A N_6 VDD mp15  l=0.13u w=0.66u m=1
.ends mi02d3
* SPICE INPUT		Tue Jul 31 19:42:10 2018	mi02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02dm
.subckt mi02dm GND Y VDD B A S0
M1 GND S0 N_4 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.36u m=1
M3 Y S0 N_2 GND mn15  l=0.13u w=0.36u m=1
M4 Y N_4 N_6 GND mn15  l=0.13u w=0.36u m=1
M5 N_6 A GND GND mn15  l=0.13u w=0.36u m=1
M6 N_4 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M7 VDD B N_2 VDD mp15  l=0.13u w=0.55u m=1
M8 Y N_4 N_2 VDD mp15  l=0.13u w=0.55u m=1
M9 Y S0 N_6 VDD mp15  l=0.13u w=0.55u m=1
M10 N_6 A VDD VDD mp15  l=0.13u w=0.55u m=1
.ends mi02dm
* SPICE INPUT		Tue Jul 31 19:42:23 2018	mx02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d0
.subckt mx02d0 VDD Y B A GND S0
M1 N_16 B GND GND mn15  l=0.13u w=0.18u m=1
M2 N_15 A GND GND mn15  l=0.13u w=0.18u m=1
M3 N_15 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M4 N_16 S0 N_6 GND mn15  l=0.13u w=0.18u m=1
M5 GND S0 N_5 GND mn15  l=0.13u w=0.18u m=1
M6 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_10 B VDD VDD mp15  l=0.13u w=0.26u m=1
M8 N_9 A VDD VDD mp15  l=0.13u w=0.26u m=1
M9 N_10 N_5 N_6 VDD mp15  l=0.13u w=0.26u m=1
M10 N_5 S0 VDD VDD mp15  l=0.13u w=0.26u m=1
M11 N_6 S0 N_9 VDD mp15  l=0.13u w=0.26u m=1
M12 Y N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mx02d0
* SPICE INPUT		Tue Jul 31 19:42:36 2018	mx02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d1
.subckt mx02d1 VDD Y GND B A S0
M1 GND S0 N_4 GND mn15  l=0.13u w=0.18u m=1
M2 N_16 S0 N_6 GND mn15  l=0.13u w=0.22u m=1
M3 N_15 A GND GND mn15  l=0.13u w=0.22u m=1
M4 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_16 B GND GND mn15  l=0.13u w=0.22u m=1
M6 N_15 N_4 N_6 GND mn15  l=0.13u w=0.22u m=1
M7 N_6 S0 N_7 VDD mp15  l=0.13u w=0.37u m=1
M8 VDD S0 N_4 VDD mp15  l=0.13u w=0.24u m=1
M9 N_7 A VDD VDD mp15  l=0.13u w=0.37u m=1
M10 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 B VDD VDD mp15  l=0.13u w=0.37u m=1
M12 N_8 N_4 N_6 VDD mp15  l=0.13u w=0.37u m=1
.ends mx02d1
* SPICE INPUT		Tue Jul 31 19:42:49 2018	mx02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d2
.subckt mx02d2 Y GND VDD B A S0
M1 N_8 N_4 N_6 GND mn15  l=0.13u w=0.32u m=1
M2 GND B N_7 GND mn15  l=0.13u w=0.3u m=1
M3 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M5 N_6 A GND GND mn15  l=0.13u w=0.3u m=1
M6 GND S0 N_4 GND mn15  l=0.13u w=0.32u m=1
M7 N_8 S0 N_7 GND mn15  l=0.13u w=0.32u m=1
M8 N_8 N_4 N_7 VDD mp15  l=0.13u w=0.5u m=1
M9 VDD B N_7 VDD mp15  l=0.13u w=0.48u m=1
M10 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M12 N_6 A VDD VDD mp15  l=0.13u w=0.48u m=1
M13 N_4 S0 VDD VDD mp15  l=0.13u w=0.46u m=1
M14 N_8 S0 N_6 VDD mp15  l=0.13u w=0.5u m=1
.ends mx02d2
* SPICE INPUT		Tue Jul 31 19:43:02 2018	mx02d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d3
.subckt mx02d3 VDD Y GND B A S0
M1 N_16 S0 GND GND mn15  l=0.13u w=0.27u m=1
M2 N_12 A GND GND mn15  l=0.13u w=0.23u m=1
M3 GND A N_12 GND mn15  l=0.13u w=0.22u m=1
M4 N_6 S0 N_9 GND mn15  l=0.13u w=0.23u m=1
M5 N_6 S0 N_9 GND mn15  l=0.13u w=0.22u m=1
M6 N_9 N_16 N_12 GND mn15  l=0.13u w=0.23u m=1
M7 N_12 N_16 N_9 GND mn15  l=0.13u w=0.22u m=1
M8 Y N_9 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_9 GND GND mn15  l=0.13u w=0.46u m=1
M10 Y N_9 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND B N_6 GND mn15  l=0.13u w=0.23u m=1
M12 N_6 B GND GND mn15  l=0.13u w=0.22u m=1
M13 Y N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 Y N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_6 B VDD VDD mp15  l=0.13u w=0.335u m=1
M17 N_6 B VDD VDD mp15  l=0.13u w=0.335u m=1
M18 N_12 S0 N_9 VDD mp15  l=0.13u w=0.335u m=1
M19 N_12 S0 N_9 VDD mp15  l=0.13u w=0.335u m=1
M20 N_9 N_16 N_6 VDD mp15  l=0.13u w=0.32u m=1
M21 N_9 N_16 N_6 VDD mp15  l=0.13u w=0.32u m=1
M22 N_16 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M23 N_12 A VDD VDD mp15  l=0.13u w=0.32u m=1
M24 VDD A N_12 VDD mp15  l=0.13u w=0.32u m=1
.ends mx02d3
* SPICE INPUT		Tue Jul 31 19:43:14 2018	mx02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02dm
.subckt mx02dm GND Y VDD B A S0
M1 N_7 A GND GND mn15  l=0.13u w=0.27u m=1
M2 Y N_6 GND GND mn15  l=0.13u w=0.36u m=1
M3 N_8 B GND GND mn15  l=0.13u w=0.27u m=1
M4 N_6 N_5 N_7 GND mn15  l=0.13u w=0.27u m=1
M5 N_8 S0 N_6 GND mn15  l=0.13u w=0.27u m=1
M6 N_5 S0 GND GND mn15  l=0.13u w=0.27u m=1
M7 N_15 A VDD VDD mp15  l=0.13u w=0.41u m=1
M8 Y N_6 VDD VDD mp15  l=0.13u w=0.55u m=1
M9 N_16 B VDD VDD mp15  l=0.13u w=0.41u m=1
M10 N_5 S0 VDD VDD mp15  l=0.13u w=0.41u m=1
M11 N_6 S0 N_15 VDD mp15  l=0.13u w=0.41u m=1
M12 N_16 N_5 N_6 VDD mp15  l=0.13u w=0.41u m=1
.ends mx02dm
* SPICE INPUT		Tue Jul 31 19:43:27 2018	mx03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx03d0
.subckt mx03d0 VDD Y C S1 A GND B S0
M1 N_6 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_8 S0 N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 S0 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_8 N_5 N_7 GND mn15  l=0.13u w=0.26u m=1
M5 GND S1 N_3 GND mn15  l=0.13u w=0.26u m=1
M6 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M7 Y N_12 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_12 N_3 N_8 GND mn15  l=0.13u w=0.26u m=1
M9 N_12 S1 N_13 GND mn15  l=0.13u w=0.26u m=1
M10 N_13 C GND GND mn15  l=0.13u w=0.26u m=1
M11 N_6 B VDD VDD mp15  l=0.13u w=0.4u m=1
M12 N_8 N_5 N_6 VDD mp15  l=0.13u w=0.26u m=1
M13 N_5 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_8 S0 N_7 VDD mp15  l=0.13u w=0.26u m=1
M15 N_3 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M17 Y N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_13 N_3 N_12 VDD mp15  l=0.13u w=0.26u m=1
M19 N_12 S1 N_8 VDD mp15  l=0.13u w=0.26u m=1
M20 N_13 C VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mx03d0
* SPICE INPUT		Tue Jul 31 19:43:41 2018	mx03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx03d1
.subckt mx03d1 VDD Y GND C S1 A B S0
M1 N_12 N_3 N_7 GND mn15  l=0.13u w=0.28u m=1
M2 N_12 S1 N_13 GND mn15  l=0.13u w=0.28u m=1
M3 N_13 C GND GND mn15  l=0.13u w=0.28u m=1
M4 Y N_12 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 B GND GND mn15  l=0.13u w=0.33u m=1
M6 N_5 S0 GND GND mn15  l=0.13u w=0.28u m=1
M7 N_7 S0 N_6 GND mn15  l=0.13u w=0.28u m=1
M8 N_8 N_5 N_7 GND mn15  l=0.13u w=0.28u m=1
M9 N_8 A GND GND mn15  l=0.13u w=0.33u m=1
M10 GND S1 N_3 GND mn15  l=0.13u w=0.28u m=1
M11 N_6 B VDD VDD mp15  l=0.13u w=0.5u m=1
M12 N_7 N_5 N_6 VDD mp15  l=0.13u w=0.28u m=1
M13 N_8 S0 N_7 VDD mp15  l=0.13u w=0.28u m=1
M14 N_5 S0 VDD VDD mp15  l=0.13u w=0.39u m=1
M15 N_8 A VDD VDD mp15  l=0.13u w=0.5u m=1
M16 N_3 S1 VDD VDD mp15  l=0.13u w=0.39u m=1
M17 N_13 N_3 N_12 VDD mp15  l=0.13u w=0.28u m=1
M18 N_12 S1 N_7 VDD mp15  l=0.13u w=0.28u m=1
M19 N_13 C VDD VDD mp15  l=0.13u w=0.42u m=1
M20 Y N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends mx03d1
* SPICE INPUT		Tue Jul 31 19:43:54 2018	mx03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx03d2
.subckt mx03d2 VDD Y A S1 GND C B S0
M1 N_3 B GND GND mn15  l=0.13u w=0.23u m=1
M2 GND B N_3 GND mn15  l=0.13u w=0.23u m=1
M3 N_5 S0 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_8 S0 N_3 GND mn15  l=0.13u w=0.37u m=1
M5 N_8 N_5 N_10 GND mn15  l=0.13u w=0.37u m=1
M6 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND S1 N_7 GND mn15  l=0.13u w=0.28u m=1
M8 GND N_14 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_14 Y GND mn15  l=0.13u w=0.46u m=1
M10 N_8 N_7 N_14 GND mn15  l=0.13u w=0.37u m=1
M11 N_15 S1 N_14 GND mn15  l=0.13u w=0.37u m=1
M12 GND C N_15 GND mn15  l=0.13u w=0.41u m=1
M13 VDD B N_3 VDD mp15  l=0.13u w=0.39u m=1
M14 N_3 B VDD VDD mp15  l=0.13u w=0.3u m=1
M15 N_5 S0 VDD VDD mp15  l=0.13u w=0.39u m=1
M16 N_3 N_5 N_8 VDD mp15  l=0.13u w=0.37u m=1
M17 N_10 S0 N_8 VDD mp15  l=0.13u w=0.37u m=1
M18 N_10 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_7 S1 VDD VDD mp15  l=0.13u w=0.39u m=1
M20 VDD N_14 Y VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_14 Y VDD mp15  l=0.13u w=0.69u m=1
M22 N_15 N_7 N_14 VDD mp15  l=0.13u w=0.37u m=1
M23 N_14 S1 N_8 VDD mp15  l=0.13u w=0.37u m=1
M24 VDD C N_15 VDD mp15  l=0.13u w=0.61u m=1
.ends mx03d2
* SPICE INPUT		Tue Jul 31 19:44:07 2018	mx03d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx03d3
.subckt mx03d3 GND Y S1 VDD C B A S0
M1 N_3 B GND GND mn15  l=0.13u w=0.23u m=1
M2 GND B N_3 GND mn15  l=0.13u w=0.23u m=1
M3 N_5 S0 GND GND mn15  l=0.13u w=0.28u m=1
M4 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_9 N_13 N_8 GND mn15  l=0.13u w=0.37u m=1
M8 GND C N_10 GND mn15  l=0.13u w=0.46u m=1
M9 N_10 S1 N_8 GND mn15  l=0.13u w=0.37u m=1
M10 N_9 S0 N_3 GND mn15  l=0.13u w=0.37u m=1
M11 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M12 N_9 N_5 N_16 GND mn15  l=0.13u w=0.37u m=1
M13 GND S1 N_13 GND mn15  l=0.13u w=0.28u m=1
M14 N_3 N_5 N_9 VDD mp15  l=0.13u w=0.37u m=1
M15 N_16 S0 N_9 VDD mp15  l=0.13u w=0.37u m=1
M16 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_13 S1 VDD VDD mp15  l=0.13u w=0.39u m=1
M18 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_10 N_13 N_8 VDD mp15  l=0.13u w=0.37u m=1
M22 N_10 C VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_8 S1 N_9 VDD mp15  l=0.13u w=0.37u m=1
M24 N_3 B VDD VDD mp15  l=0.13u w=0.3u m=1
M25 VDD B N_3 VDD mp15  l=0.13u w=0.39u m=1
M26 N_5 S0 VDD VDD mp15  l=0.13u w=0.39u m=1
.ends mx03d3
* SPICE INPUT		Tue Jul 31 19:44:19 2018	mx04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d0
.subckt mx04d0 VDD Y S1 B A D S0 GND C
M1 N_68 C GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 N_4 N_68 GND mn15  l=0.13u w=0.26u m=1
M3 N_69 D GND GND mn15  l=0.13u w=0.26u m=1
M4 N_70 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_2 N_4 N_67 GND mn15  l=0.13u w=0.26u m=1
M6 N_70 S0 N_2 GND mn15  l=0.13u w=0.26u m=1
M7 N_69 S0 N_5 GND mn15  l=0.13u w=0.26u m=1
M8 N_4 S0 GND GND mn15  l=0.13u w=0.26u m=1
M9 N_67 A GND GND mn15  l=0.13u w=0.26u m=1
M10 Y N_7 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_13 S1 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_2 N_13 N_7 GND mn15  l=0.13u w=0.26u m=1
M13 N_5 S1 N_7 GND mn15  l=0.13u w=0.26u m=1
M14 N_15 C VDD VDD mp15  l=0.13u w=0.4u m=1
M15 N_15 S0 N_5 VDD mp15  l=0.13u w=0.4u m=1
M16 N_16 N_4 N_5 VDD mp15  l=0.13u w=0.4u m=1
M17 VDD D N_16 VDD mp15  l=0.13u w=0.4u m=1
M18 VDD B N_14 VDD mp15  l=0.13u w=0.4u m=1
M19 N_2 N_4 N_14 VDD mp15  l=0.13u w=0.4u m=1
M20 N_4 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_5 N_13 N_7 VDD mp15  l=0.13u w=0.26u m=1
M22 N_2 S1 N_7 VDD mp15  l=0.13u w=0.26u m=1
M23 N_17 S0 N_2 VDD mp15  l=0.13u w=0.4u m=1
M24 N_17 A VDD VDD mp15  l=0.13u w=0.4u m=1
M25 Y N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M26 N_13 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mx04d0
* SPICE INPUT		Tue Jul 31 19:44:32 2018	mx04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d1
.subckt mx04d1 VDD Y A B S1 D S0 C GND
M1 N_69 C GND GND mn15  l=0.13u w=0.32u m=1
M2 N_69 N_4 N_5 GND mn15  l=0.13u w=0.32u m=1
M3 GND D N_70 GND mn15  l=0.13u w=0.32u m=1
M4 N_71 B GND GND mn15  l=0.13u w=0.32u m=1
M5 N_2 N_4 N_68 GND mn15  l=0.13u w=0.32u m=1
M6 N_68 A GND GND mn15  l=0.13u w=0.32u m=1
M7 N_4 S0 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_2 S0 N_71 GND mn15  l=0.13u w=0.32u m=1
M9 N_70 S0 N_5 GND mn15  l=0.13u w=0.32u m=1
M10 N_2 N_14 N_9 GND mn15  l=0.13u w=0.28u m=1
M11 N_5 S1 N_9 GND mn15  l=0.13u w=0.28u m=1
M12 Y N_9 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_14 S1 GND GND mn15  l=0.13u w=0.26u m=1
M14 N_16 C VDD VDD mp15  l=0.13u w=0.47u m=1
M15 N_16 S0 N_5 VDD mp15  l=0.13u w=0.47u m=1
M16 N_17 N_4 N_5 VDD mp15  l=0.13u w=0.47u m=1
M17 N_17 D VDD VDD mp15  l=0.13u w=0.47u m=1
M18 VDD B N_15 VDD mp15  l=0.13u w=0.47u m=1
M19 N_2 N_4 N_15 VDD mp15  l=0.13u w=0.47u m=1
M20 N_4 S0 VDD VDD mp15  l=0.13u w=0.42u m=1
M21 VDD A N_18 VDD mp15  l=0.13u w=0.47u m=1
M22 N_2 S0 N_18 VDD mp15  l=0.13u w=0.47u m=1
M23 N_5 N_14 N_9 VDD mp15  l=0.13u w=0.28u m=1
M24 N_2 S1 N_9 VDD mp15  l=0.13u w=0.28u m=1
M25 Y N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_14 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mx04d1
* SPICE INPUT		Tue Jul 31 19:44:45 2018	mx04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d2
.subckt mx04d2 GND Y VDD S1 A S0 B D C
M1 N_3 S0 GND GND mn15  l=0.13u w=0.37u m=1
M2 N_21 N_3 N_4 GND mn15  l=0.13u w=0.225u m=1
M3 N_22 C GND GND mn15  l=0.13u w=0.225u m=1
M4 N_21 C GND GND mn15  l=0.13u w=0.225u m=1
M5 GND D N_20 GND mn15  l=0.13u w=0.225u m=1
M6 N_23 D GND GND mn15  l=0.13u w=0.225u m=1
M7 N_20 S0 N_4 GND mn15  l=0.13u w=0.225u m=1
M8 N_23 S0 N_4 GND mn15  l=0.13u w=0.225u m=1
M9 N_22 N_3 N_4 GND mn15  l=0.13u w=0.225u m=1
M10 N_10 S0 N_24 GND mn15  l=0.13u w=0.45u m=1
M11 N_24 B GND GND mn15  l=0.13u w=0.45u m=1
M12 N_10 N_3 N_25 GND mn15  l=0.13u w=0.45u m=1
M13 N_25 A GND GND mn15  l=0.13u w=0.45u m=1
M14 N_10 N_18 N_13 GND mn15  l=0.13u w=0.32u m=1
M15 N_4 S1 N_13 GND mn15  l=0.13u w=0.36u m=1
M16 GND S1 N_18 GND mn15  l=0.13u w=0.26u m=1
M17 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M18 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M19 N_3 S0 VDD VDD mp15  l=0.13u w=0.55u m=1
M20 N_107 C VDD VDD mp15  l=0.13u w=0.32u m=1
M21 N_106 C VDD VDD mp15  l=0.13u w=0.33u m=1
M22 N_108 D VDD VDD mp15  l=0.13u w=0.29u m=1
M23 VDD D N_105 VDD mp15  l=0.13u w=0.36u m=1
M24 N_106 S0 N_4 VDD mp15  l=0.13u w=0.33u m=1
M25 N_107 S0 N_4 VDD mp15  l=0.13u w=0.32u m=1
M26 N_108 N_3 N_4 VDD mp15  l=0.13u w=0.29u m=1
M27 N_4 N_3 N_105 VDD mp15  l=0.13u w=0.36u m=1
M28 N_110 B VDD VDD mp15  l=0.13u w=0.31u m=1
M29 VDD B N_109 VDD mp15  l=0.13u w=0.34u m=1
M30 N_10 N_3 N_110 VDD mp15  l=0.13u w=0.31u m=1
M31 N_10 N_3 N_109 VDD mp15  l=0.13u w=0.34u m=1
M32 N_111 A VDD VDD mp15  l=0.13u w=0.31u m=1
M33 N_112 A VDD VDD mp15  l=0.13u w=0.3u m=1
M34 N_111 S0 N_10 VDD mp15  l=0.13u w=0.31u m=1
M35 N_10 S0 N_112 VDD mp15  l=0.13u w=0.3u m=1
M36 N_13 N_18 N_4 VDD mp15  l=0.13u w=0.35u m=1
M37 N_10 S1 N_13 VDD mp15  l=0.13u w=0.35u m=1
M38 N_18 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
M39 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
M40 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
.ends mx04d2
* SPICE INPUT		Tue Jul 31 19:44:58 2018	mx04d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d3
.subckt mx04d3 GND Y S0 S1 B D A VDD C
M1 N_3 S0 GND GND mn15  l=0.13u w=0.36u m=1
M2 N_21 S0 N_4 GND mn15  l=0.13u w=0.225u m=1
M3 N_24 S0 N_4 GND mn15  l=0.13u w=0.225u m=1
M4 N_22 N_3 N_4 GND mn15  l=0.13u w=0.225u m=1
M5 N_23 N_3 N_4 GND mn15  l=0.13u w=0.225u m=1
M6 N_23 C GND GND mn15  l=0.13u w=0.225u m=1
M7 N_22 C GND GND mn15  l=0.13u w=0.225u m=1
M8 GND D N_21 GND mn15  l=0.13u w=0.225u m=1
M9 N_24 D GND GND mn15  l=0.13u w=0.225u m=1
M10 N_10 S0 N_25 GND mn15  l=0.13u w=0.45u m=1
M11 N_25 B GND GND mn15  l=0.13u w=0.45u m=1
M12 N_10 N_3 N_26 GND mn15  l=0.13u w=0.45u m=1
M13 N_26 A GND GND mn15  l=0.13u w=0.45u m=1
M14 N_4 S1 N_13 GND mn15  l=0.13u w=0.45u m=1
M15 N_10 N_18 N_13 GND mn15  l=0.13u w=0.32u m=1
M16 GND S1 N_18 GND mn15  l=0.13u w=0.28u m=1
M17 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M18 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M19 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M20 N_3 S0 VDD VDD mp15  l=0.13u w=0.53u m=1
M21 N_50 S0 N_4 VDD mp15  l=0.13u w=0.33u m=1
M22 N_51 S0 N_4 VDD mp15  l=0.13u w=0.32u m=1
M23 N_52 N_3 N_4 VDD mp15  l=0.13u w=0.29u m=1
M24 N_4 N_3 N_49 VDD mp15  l=0.13u w=0.36u m=1
M25 N_51 C VDD VDD mp15  l=0.13u w=0.32u m=1
M26 N_50 C VDD VDD mp15  l=0.13u w=0.33u m=1
M27 VDD D N_49 VDD mp15  l=0.13u w=0.36u m=1
M28 N_52 D VDD VDD mp15  l=0.13u w=0.29u m=1
M29 N_54 N_3 N_10 VDD mp15  l=0.13u w=0.32u m=1
M30 N_10 N_3 N_53 VDD mp15  l=0.13u w=0.33u m=1
M31 N_54 B VDD VDD mp15  l=0.13u w=0.32u m=1
M32 VDD B N_53 VDD mp15  l=0.13u w=0.33u m=1
M33 N_56 A VDD VDD mp15  l=0.13u w=0.31u m=1
M34 N_55 A VDD VDD mp15  l=0.13u w=0.31u m=1
M35 N_10 S1 N_13 VDD mp15  l=0.13u w=0.53u m=1
M36 N_4 N_18 N_13 VDD mp15  l=0.13u w=0.53u m=1
M37 N_55 S0 N_10 VDD mp15  l=0.13u w=0.31u m=1
M38 N_10 S0 N_56 VDD mp15  l=0.13u w=0.31u m=1
M39 N_18 S1 VDD VDD mp15  l=0.13u w=0.42u m=1
M40 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M42 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends mx04d3
* SPICE INPUT		Tue Jul 31 19:45:11 2018	mx04dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04dm
.subckt mx04dm VDD Y GND A D B S1 S0 C
M1 Y N_5 GND GND mn15  l=0.13u w=0.36u m=1
M2 N_4 S1 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_69 D GND GND mn15  l=0.13u w=0.26u m=1
M4 N_70 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 N_11 N_67 GND mn15  l=0.13u w=0.26u m=1
M6 N_11 S0 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_70 S0 N_8 GND mn15  l=0.13u w=0.26u m=1
M8 N_69 S0 N_6 GND mn15  l=0.13u w=0.26u m=1
M9 N_67 A GND GND mn15  l=0.13u w=0.26u m=1
M10 N_68 C GND GND mn15  l=0.13u w=0.26u m=1
M11 N_6 N_11 N_68 GND mn15  l=0.13u w=0.26u m=1
M12 N_8 N_4 N_5 GND mn15  l=0.13u w=0.26u m=1
M13 N_6 S1 N_5 GND mn15  l=0.13u w=0.26u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.55u m=1
M15 N_4 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.26u m=1
M17 N_14 S0 N_8 VDD mp15  l=0.13u w=0.4u m=1
M18 N_8 S1 N_5 VDD mp15  l=0.13u w=0.26u m=1
M19 N_14 A VDD VDD mp15  l=0.13u w=0.4u m=1
M20 VDD D N_17 VDD mp15  l=0.13u w=0.4u m=1
M21 N_16 S0 N_6 VDD mp15  l=0.13u w=0.4u m=1
M22 VDD B N_15 VDD mp15  l=0.13u w=0.4u m=1
M23 N_8 N_11 N_15 VDD mp15  l=0.13u w=0.4u m=1
M24 N_11 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M25 N_16 C VDD VDD mp15  l=0.13u w=0.4u m=1
M26 N_17 N_11 N_6 VDD mp15  l=0.13u w=0.4u m=1
.ends mx04dm
* SPICE INPUT		Tue Jul 31 19:45:23 2018	nd02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d0
.subckt nd02d0 VDD Y GND B A
M1 GND A N_14 GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.26u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.35u m=1
M4 Y B VDD VDD mp15  l=0.13u w=0.35u m=1
.ends nd02d0
* SPICE INPUT		Tue Jul 31 19:45:36 2018	nd02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d1
.subckt nd02d1 Y VDD A B GND
M1 GND A N_14 GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.46u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
.ends nd02d1
* SPICE INPUT		Tue Jul 31 19:45:49 2018	nd02d1p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d1p5
.subckt nd02d1p5 Y VDD A B GND
M1 GND A N_14 GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.46u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
.ends nd02d1p5
* SPICE INPUT		Tue Jul 31 19:46:02 2018	nd02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d2
.subckt nd02d2 GND Y VDD A B
M1 Y B N_5 GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M5 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M6 Y B VDD VDD mp15  l=0.13u w=0.61u m=1
M7 Y A VDD VDD mp15  l=0.13u w=0.61u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.61u m=1
.ends nd02d2
* SPICE INPUT		Tue Jul 31 19:46:15 2018	nd02d2p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d2p5
.subckt nd02d2p5 GND Y A B VDD
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_5 GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M5 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nd02d2p5
* SPICE INPUT		Tue Jul 31 19:46:28 2018	nd02d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d3
.subckt nd02d3 Y GND A VDD B
M1 N_3 B Y GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B Y GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B Y GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B Y GND mn15  l=0.13u w=0.46u m=1
M5 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M8 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M9 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M10 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M11 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M12 Y B VDD VDD mp15  l=0.13u w=0.61u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.61u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
M16 Y A VDD VDD mp15  l=0.13u w=0.61u m=1
.ends nd02d3
* SPICE INPUT		Tue Jul 31 19:46:41 2018	nd02d3p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d3p5
.subckt nd02d3p5 GND Y VDD A B
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_9 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_8 GND mn15  l=0.13u w=0.46u m=1
M4 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_7 GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M8 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M11 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nd02d3p5
* SPICE INPUT		Tue Jul 31 19:46:54 2018	nd02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02dm
.subckt nd02dm Y VDD GND A B
M1 GND A N_14 GND mn15  l=0.13u w=0.36u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.36u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.45u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.45u m=1
.ends nd02dm
* SPICE INPUT		Tue Jul 31 19:47:07 2018	nd02od
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02od
.subckt nd02od VDD B GND A Y
M1 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_22 B N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_3 N_5 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_22 A GND GND mn15  l=0.13u w=0.26u m=1
M5 N_5 B VDD VDD mp15  l=0.13u w=0.35u m=1
M6 N_3 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_5 A VDD VDD mp15  l=0.13u w=0.35u m=1
.ends nd02od
* SPICE INPUT		Tue Jul 31 19:47:20 2018	nd03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d0
.subckt nd03d0 VDD Y C B A GND
M1 N_19 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_19 B N_18 GND mn15  l=0.13u w=0.26u m=1
M3 Y C N_18 GND mn15  l=0.13u w=0.26u m=1
M4 Y A VDD VDD mp15  l=0.13u w=0.31u m=1
M5 Y B VDD VDD mp15  l=0.13u w=0.31u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.31u m=1
.ends nd03d0
* SPICE INPUT		Tue Jul 31 19:47:34 2018	nd03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d1
.subckt nd03d1 VDD Y C B A GND
M1 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y C N_18 GND mn15  l=0.13u w=0.46u m=1
M3 N_19 B N_18 GND mn15  l=0.13u w=0.46u m=1
M4 Y A VDD VDD mp15  l=0.13u w=0.54u m=1
M5 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M6 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
.ends nd03d1
* SPICE INPUT		Tue Jul 31 19:47:46 2018	nd03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d2
.subckt nd03d2 GND Y B C A VDD
M1 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_8 B N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 C Y GND mn15  l=0.13u w=0.46u m=1
M5 Y C N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M8 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
M9 VDD B Y VDD mp15  l=0.13u w=0.54u m=1
M10 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M11 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.54u m=1
.ends nd03d2
* SPICE INPUT		Tue Jul 31 19:47:59 2018	nd03d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d3
.subckt nd03d3 VDD Y GND C B A
M1 N_18 B N_19 GND mn15  l=0.13u w=0.46u m=1
M2 N_19 B N_18 GND mn15  l=0.13u w=0.46u m=1
M3 N_18 B N_19 GND mn15  l=0.13u w=0.46u m=1
M4 N_18 B N_19 GND mn15  l=0.13u w=0.46u m=1
M5 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_19 GND mn15  l=0.13u w=0.46u m=1
M7 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M8 GND A N_19 GND mn15  l=0.13u w=0.46u m=1
M9 Y C N_18 GND mn15  l=0.13u w=0.46u m=1
M10 Y C N_18 GND mn15  l=0.13u w=0.46u m=1
M11 N_18 C Y GND mn15  l=0.13u w=0.46u m=1
M12 N_18 C Y GND mn15  l=0.13u w=0.46u m=1
M13 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M14 VDD B Y VDD mp15  l=0.13u w=0.54u m=1
M15 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M16 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M17 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
M18 Y A VDD VDD mp15  l=0.13u w=0.54u m=1
M19 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
M20 Y A VDD VDD mp15  l=0.13u w=0.54u m=1
M21 VDD C Y VDD mp15  l=0.13u w=0.54u m=1
M22 VDD C Y VDD mp15  l=0.13u w=0.54u m=1
M23 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M24 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
.ends nd03d3
* SPICE INPUT		Tue Jul 31 19:48:12 2018	nd03od
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03od
.subckt nd03od GND Y VDD A B C
M1 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 C N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 N_6 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 B N_7 GND mn15  l=0.13u w=0.26u m=1
M6 N_6 C VDD VDD mp15  l=0.13u w=0.31u m=1
M7 N_5 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_6 A VDD VDD mp15  l=0.13u w=0.31u m=1
M9 N_6 B VDD VDD mp15  l=0.13u w=0.31u m=1
.ends nd03od
* SPICE INPUT		Tue Jul 31 19:48:25 2018	nd04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d0
.subckt nd04d0 VDD Y GND D C B A
M1 N_17 C N_15 GND mn15  l=0.13u w=0.26u m=1
M2 Y D N_15 GND mn15  l=0.13u w=0.26u m=1
M3 N_17 B N_16 GND mn15  l=0.13u w=0.26u m=1
M4 N_16 A GND GND mn15  l=0.13u w=0.26u m=1
M5 VDD C Y VDD mp15  l=0.13u w=0.29u m=1
M6 Y D VDD VDD mp15  l=0.13u w=0.29u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.29u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.29u m=1
.ends nd04d0
* SPICE INPUT		Tue Jul 31 19:48:38 2018	nd04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d1
.subckt nd04d1 Y VDD A D C B GND
M1 Y D N_15 GND mn15  l=0.13u w=0.46u m=1
M2 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_17 B N_16 GND mn15  l=0.13u w=0.46u m=1
M4 N_17 C N_15 GND mn15  l=0.13u w=0.46u m=1
M5 VDD D Y VDD mp15  l=0.13u w=0.52u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M7 VDD B Y VDD mp15  l=0.13u w=0.52u m=1
M8 VDD C Y VDD mp15  l=0.13u w=0.52u m=1
.ends nd04d1
* SPICE INPUT		Tue Jul 31 19:48:51 2018	nd04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d2
.subckt nd04d2 VDD Y GND D C B A
M1 N_12 C N_15 GND mn15  l=0.13u w=0.46u m=1
M2 N_12 C N_15 GND mn15  l=0.13u w=0.46u m=1
M3 N_12 D Y GND mn15  l=0.13u w=0.46u m=1
M4 N_12 D Y GND mn15  l=0.13u w=0.46u m=1
M5 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_16 GND mn15  l=0.13u w=0.46u m=1
M7 N_16 B N_15 GND mn15  l=0.13u w=0.46u m=1
M8 N_16 B N_15 GND mn15  l=0.13u w=0.46u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M11 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M12 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M14 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M15 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M16 VDD D Y VDD mp15  l=0.13u w=0.52u m=1
.ends nd04d2
* SPICE INPUT		Tue Jul 31 19:49:04 2018	nd04d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d3
.subckt nd04d3 GND VDD Y D C B A
M1 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M2 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M3 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M6 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M7 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M9 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M10 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M11 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M12 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M13 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M14 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M15 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M16 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M17 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M18 VDD B Y VDD mp15  l=0.13u w=0.52u m=1
M19 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M20 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M21 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M23 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M25 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M26 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M27 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M28 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M29 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M30 VDD D Y VDD mp15  l=0.13u w=0.52u m=1
M31 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M32 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
.ends nd04d3
* SPICE INPUT		Tue Jul 31 19:49:18 2018	nd12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d0
.subckt nd12d0 Y GND B VDD AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 GND N_3 N_5 GND mn15  l=0.13u w=0.26u m=1
M3 Y B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_3 AN VDD VDD mp15  l=0.13u w=0.4u m=1
M5 VDD N_3 Y VDD mp15  l=0.13u w=0.35u m=1
M6 Y B VDD VDD mp15  l=0.13u w=0.35u m=1
.ends nd12d0
* SPICE INPUT		Tue Jul 31 19:49:31 2018	nd12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d1
.subckt nd12d1 Y GND VDD B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.3u m=1
M2 GND N_3 N_5 GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_5 GND mn15  l=0.13u w=0.46u m=1
M4 VDD AN N_3 VDD mp15  l=0.13u w=0.45u m=1
M5 VDD N_3 Y VDD mp15  l=0.13u w=0.63u m=1
M6 VDD B Y VDD mp15  l=0.13u w=0.63u m=1
.ends nd12d1
* SPICE INPUT		Tue Jul 31 19:49:43 2018	nd12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d2
.subckt nd12d2 GND Y VDD B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M4 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_3 N_6 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y N_3 VDD VDD mp15  l=0.13u w=0.63u m=1
M8 VDD B Y VDD mp15  l=0.13u w=0.63u m=1
M9 Y B VDD VDD mp15  l=0.13u w=0.63u m=1
M10 Y N_3 VDD VDD mp15  l=0.13u w=0.63u m=1
.ends nd12d2
* SPICE INPUT		Tue Jul 31 19:49:56 2018	nd12d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d3
.subckt nd12d3 GND Y VDD B AN
M1 GND AN N_4 GND mn15  l=0.13u w=0.4u m=1
M2 N_4 AN GND GND mn15  l=0.13u w=0.4u m=1
M3 N_10 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_11 B Y GND mn15  l=0.13u w=0.46u m=1
M5 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M6 Y B N_9 GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_12 GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 N_9 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_11 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M11 VDD AN N_4 VDD mp15  l=0.13u w=0.55u m=1
M12 N_4 AN VDD VDD mp15  l=0.13u w=0.55u m=1
M13 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M14 Y B VDD VDD mp15  l=0.13u w=0.61u m=1
M15 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M16 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M17 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M20 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
.ends nd12d3
* SPICE INPUT		Tue Jul 31 19:50:08 2018	nd12dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12dm
.subckt nd12dm Y GND AN VDD B
M1 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_5 GND mn15  l=0.13u w=0.36u m=1
M3 GND N_3 N_5 GND mn15  l=0.13u w=0.36u m=1
M4 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
M5 VDD B Y VDD mp15  l=0.13u w=0.45u m=1
M6 VDD N_3 Y VDD mp15  l=0.13u w=0.45u m=1
.ends nd12dm
* SPICE INPUT		Tue Jul 31 19:50:21 2018	nd13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d0
.subckt nd13d0 Y GND AN C B VDD
M1 N_6 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M2 Y C N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M5 Y N_3 VDD VDD mp15  l=0.13u w=0.31u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.31u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.31u m=1
M8 N_3 AN VDD VDD mp15  l=0.13u w=0.4u m=1
.ends nd13d0
* SPICE INPUT		Tue Jul 31 19:50:34 2018	nd13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d1
.subckt nd13d1 Y GND C VDD B AN
M1 N_6 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M2 Y C N_5 GND mn15  l=0.13u w=0.46u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.3u m=1
M4 N_6 B N_5 GND mn15  l=0.13u w=0.46u m=1
M5 Y N_3 VDD VDD mp15  l=0.13u w=0.56u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.56u m=1
M7 VDD AN N_3 VDD mp15  l=0.13u w=0.45u m=1
M8 Y B VDD VDD mp15  l=0.13u w=0.56u m=1
.ends nd13d1
* SPICE INPUT		Tue Jul 31 19:50:47 2018	nd13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d2
.subckt nd13d2 GND Y VDD B C AN
M1 N_9 B N_6 GND mn15  l=0.13u w=0.46u m=1
M2 GND N_4 N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_4 AN GND GND mn15  l=0.13u w=0.36u m=1
M4 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M5 N_7 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_9 C Y GND mn15  l=0.13u w=0.46u m=1
M7 N_8 C Y GND mn15  l=0.13u w=0.46u m=1
M8 VDD B Y VDD mp15  l=0.13u w=0.56u m=1
M9 VDD N_4 Y VDD mp15  l=0.13u w=0.56u m=1
M10 N_4 AN VDD VDD mp15  l=0.13u w=0.55u m=1
M11 Y B VDD VDD mp15  l=0.13u w=0.56u m=1
M12 Y N_4 VDD VDD mp15  l=0.13u w=0.56u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.56u m=1
M14 Y C VDD VDD mp15  l=0.13u w=0.56u m=1
.ends nd13d2
* SPICE INPUT		Tue Jul 31 19:51:00 2018	nd13d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d3
.subckt nd13d3 Y VDD AN B GND C
M1 N_5 AN GND GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 N_18 GND mn15  l=0.13u w=0.46u m=1
M3 GND N_5 N_18 GND mn15  l=0.13u w=0.46u m=1
M4 GND N_5 N_18 GND mn15  l=0.13u w=0.46u m=1
M5 N_18 N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_21 B N_18 GND mn15  l=0.13u w=0.46u m=1
M7 N_21 B N_18 GND mn15  l=0.13u w=0.46u m=1
M8 N_21 B N_18 GND mn15  l=0.13u w=0.46u m=1
M9 N_21 B N_18 GND mn15  l=0.13u w=0.46u m=1
M10 N_21 C Y GND mn15  l=0.13u w=0.46u m=1
M11 N_21 C Y GND mn15  l=0.13u w=0.46u m=1
M12 N_21 C Y GND mn15  l=0.13u w=0.46u m=1
M13 N_21 C Y GND mn15  l=0.13u w=0.46u m=1
M14 N_5 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_5 Y VDD mp15  l=0.13u w=0.54u m=1
M16 VDD N_5 Y VDD mp15  l=0.13u w=0.54u m=1
M17 VDD N_5 Y VDD mp15  l=0.13u w=0.54u m=1
M18 Y N_5 VDD VDD mp15  l=0.13u w=0.54u m=1
M19 VDD B Y VDD mp15  l=0.13u w=0.54u m=1
M20 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M21 VDD B Y VDD mp15  l=0.13u w=0.54u m=1
M22 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M23 VDD C Y VDD mp15  l=0.13u w=0.54u m=1
M24 VDD C Y VDD mp15  l=0.13u w=0.54u m=1
M25 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M26 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
.ends nd13d3
* SPICE INPUT		Tue Jul 31 19:51:13 2018	nd14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d0
.subckt nd14d0 Y GND VDD D C B AN
M1 N_7 C N_5 GND mn15  l=0.13u w=0.26u m=1
M2 Y D N_5 GND mn15  l=0.13u w=0.26u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M5 N_6 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M6 VDD C Y VDD mp15  l=0.13u w=0.29u m=1
M7 Y D VDD VDD mp15  l=0.13u w=0.29u m=1
M8 N_3 AN VDD VDD mp15  l=0.13u w=0.4u m=1
M9 Y B VDD VDD mp15  l=0.13u w=0.29u m=1
M10 Y N_3 VDD VDD mp15  l=0.13u w=0.29u m=1
.ends nd14d0
* SPICE INPUT		Tue Jul 31 19:51:27 2018	nd14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d1
.subckt nd14d1 Y GND VDD D C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.3u m=1
M2 N_7 C N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M4 Y D N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_6 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 AN VDD VDD mp15  l=0.13u w=0.45u m=1
M7 VDD C Y VDD mp15  l=0.13u w=0.52u m=1
M8 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M9 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M10 Y N_3 VDD VDD mp15  l=0.13u w=0.52u m=1
.ends nd14d1
* SPICE INPUT		Tue Jul 31 19:51:39 2018	nd14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d2
.subckt nd14d2 VDD Y GND D C B AN
M1 N_3 AN GND GND mn15  l=0.13u w=0.4u m=1
M2 N_18 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND N_3 N_18 GND mn15  l=0.13u w=0.46u m=1
M4 N_18 B N_17 GND mn15  l=0.13u w=0.46u m=1
M5 N_18 B N_17 GND mn15  l=0.13u w=0.46u m=1
M6 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M7 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_14 C N_17 GND mn15  l=0.13u w=0.46u m=1
M9 N_14 C N_17 GND mn15  l=0.13u w=0.46u m=1
M10 N_3 AN VDD VDD mp15  l=0.13u w=0.6u m=1
M11 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M12 VDD D Y VDD mp15  l=0.13u w=0.52u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M14 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M15 Y N_3 VDD VDD mp15  l=0.13u w=0.52u m=1
M16 Y N_3 VDD VDD mp15  l=0.13u w=0.52u m=1
M17 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M18 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
.ends nd14d2
* SPICE INPUT		Tue Jul 31 19:51:53 2018	nd14d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d3
.subckt nd14d3 GND VDD Y D C B AN
M1 GND AN N_12 GND mn15  l=0.13u w=0.4u m=1
M2 GND AN N_12 GND mn15  l=0.13u w=0.4u m=1
M3 N_11 N_12 GND GND mn15  l=0.13u w=0.46u m=1
M4 GND N_12 N_11 GND mn15  l=0.13u w=0.46u m=1
M5 N_11 N_12 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_12 N_11 GND mn15  l=0.13u w=0.46u m=1
M7 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M8 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M9 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M10 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M11 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M12 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M13 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M14 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M15 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M16 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M17 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M18 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M19 VDD AN N_12 VDD mp15  l=0.13u w=0.58u m=1
M20 VDD AN N_12 VDD mp15  l=0.13u w=0.58u m=1
M21 VDD N_12 Y VDD mp15  l=0.13u w=0.5u m=1
M22 Y N_12 VDD VDD mp15  l=0.13u w=0.5u m=1
M23 VDD N_12 Y VDD mp15  l=0.13u w=0.5u m=1
M24 Y N_12 VDD VDD mp15  l=0.13u w=0.5u m=1
M25 Y B VDD VDD mp15  l=0.13u w=0.5u m=1
M26 Y B VDD VDD mp15  l=0.13u w=0.5u m=1
M27 Y B VDD VDD mp15  l=0.13u w=0.5u m=1
M28 Y B VDD VDD mp15  l=0.13u w=0.5u m=1
M29 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M30 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M31 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M32 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M33 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M34 VDD D Y VDD mp15  l=0.13u w=0.5u m=1
M35 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M36 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
.ends nd14d3
* SPICE INPUT		Tue Jul 31 19:52:07 2018	nd24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d0
.subckt nd24d0 Y GND BN D AN VDD C
M1 N_9 N_5 N_8 GND mn15  l=0.13u w=0.26u m=1
M2 N_9 C N_7 GND mn15  l=0.13u w=0.26u m=1
M3 N_8 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 D Y GND mn15  l=0.13u w=0.26u m=1
M5 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M6 GND BN N_5 GND mn15  l=0.13u w=0.26u m=1
M7 N_5 BN VDD VDD mp15  l=0.13u w=0.4u m=1
M8 VDD N_5 Y VDD mp15  l=0.13u w=0.29u m=1
M9 Y C VDD VDD mp15  l=0.13u w=0.29u m=1
M10 Y N_3 VDD VDD mp15  l=0.13u w=0.29u m=1
M11 Y D VDD VDD mp15  l=0.13u w=0.29u m=1
M12 N_3 AN VDD VDD mp15  l=0.13u w=0.4u m=1
.ends nd24d0
* SPICE INPUT		Tue Jul 31 19:52:20 2018	nd24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d1
.subckt nd24d1 GND Y BN AN D C VDD
M1 GND BN N_2 GND mn15  l=0.13u w=0.3u m=1
M2 GND AN N_5 GND mn15  l=0.13u w=0.3u m=1
M3 N_8 N_5 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_9 N_2 N_8 GND mn15  l=0.13u w=0.46u m=1
M5 N_9 C N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_7 D Y GND mn15  l=0.13u w=0.46u m=1
M7 N_2 BN VDD VDD mp15  l=0.13u w=0.43u m=1
M8 VDD AN N_5 VDD mp15  l=0.13u w=0.43u m=1
M9 Y N_5 VDD VDD mp15  l=0.13u w=0.5u m=1
M10 Y N_2 VDD VDD mp15  l=0.13u w=0.5u m=1
M11 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M12 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
.ends nd24d1
* SPICE INPUT		Tue Jul 31 19:52:33 2018	nd24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d2
.subckt nd24d2 GND Y BN AN VDD D C
M1 N_3 AN GND GND mn15  l=0.13u w=0.4u m=1
M2 N_4 BN GND GND mn15  l=0.13u w=0.4u m=1
M3 N_6 N_4 N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_6 N_4 N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_6 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_3 N_6 GND mn15  l=0.13u w=0.46u m=1
M7 N_11 C N_5 GND mn15  l=0.13u w=0.46u m=1
M8 N_11 C N_5 GND mn15  l=0.13u w=0.46u m=1
M9 N_11 D Y GND mn15  l=0.13u w=0.46u m=1
M10 N_11 D Y GND mn15  l=0.13u w=0.46u m=1
M11 N_3 AN VDD VDD mp15  l=0.13u w=0.58u m=1
M12 N_4 BN VDD VDD mp15  l=0.13u w=0.58u m=1
M13 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M14 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M15 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M16 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M17 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M18 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M19 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M20 VDD D Y VDD mp15  l=0.13u w=0.5u m=1
.ends nd24d2
* SPICE INPUT		Tue Jul 31 19:52:46 2018	nd24d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d3
.subckt nd24d3 VDD Y GND D C AN BN
M1 N_4 BN GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.46u m=1
M3 N_27 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_27 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_27 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_27 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_27 N_4 N_26 GND mn15  l=0.13u w=0.46u m=1
M8 N_27 N_4 N_26 GND mn15  l=0.13u w=0.46u m=1
M9 N_27 N_4 N_26 GND mn15  l=0.13u w=0.46u m=1
M10 N_27 N_4 N_26 GND mn15  l=0.13u w=0.46u m=1
M11 N_23 C N_26 GND mn15  l=0.13u w=0.46u m=1
M12 N_23 C N_26 GND mn15  l=0.13u w=0.46u m=1
M13 N_23 C N_26 GND mn15  l=0.13u w=0.46u m=1
M14 N_23 C N_26 GND mn15  l=0.13u w=0.46u m=1
M15 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M16 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M17 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M18 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M19 N_4 BN VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_3 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M21 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M22 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M23 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M24 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M25 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M26 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M27 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M28 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M29 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M30 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M31 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M32 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M33 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M34 VDD D Y VDD mp15  l=0.13u w=0.5u m=1
M35 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M36 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
.ends nd24d3
* SPICE INPUT		Tue Jul 31 19:52:58 2018	nr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d0
.subckt nr02d0 Y GND VDD B A
M1 GND B Y GND mn15  l=0.13u w=0.26u m=1
M2 GND A Y GND mn15  l=0.13u w=0.26u m=1
M3 Y B N_8 VDD mp15  l=0.13u w=0.4u m=1
M4 VDD A N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends nr02d0
* SPICE INPUT		Tue Jul 31 19:53:11 2018	nr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d1
.subckt nr02d1 Y GND VDD B A
M1 GND B Y GND mn15  l=0.13u w=0.34u m=1
M2 GND A Y GND mn15  l=0.13u w=0.34u m=1
M3 Y B N_8 VDD mp15  l=0.13u w=0.69u m=1
M4 VDD A N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends nr02d1
* SPICE INPUT		Tue Jul 31 19:53:24 2018	nr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d2
.subckt nr02d2 VDD Y GND A B
M1 GND B Y GND mn15  l=0.13u w=0.34u m=1
M2 Y B GND GND mn15  l=0.13u w=0.34u m=1
M3 Y A GND GND mn15  l=0.13u w=0.34u m=1
M4 GND A Y GND mn15  l=0.13u w=0.34u m=1
M5 Y B N_5 VDD mp15  l=0.13u w=0.69u m=1
M6 Y B N_6 VDD mp15  l=0.13u w=0.69u m=1
M7 N_6 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends nr02d2
* SPICE INPUT		Tue Jul 31 19:53:38 2018	nr02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d4
.subckt nr02d4 Y GND VDD B A
M1 GND A Y GND mn15  l=0.13u w=0.34u m=1
M2 Y A GND GND mn15  l=0.13u w=0.34u m=1
M3 GND A Y GND mn15  l=0.13u w=0.34u m=1
M4 Y A GND GND mn15  l=0.13u w=0.34u m=1
M5 GND B Y GND mn15  l=0.13u w=0.34u m=1
M6 GND B Y GND mn15  l=0.13u w=0.34u m=1
M7 GND B Y GND mn15  l=0.13u w=0.34u m=1
M8 Y B GND GND mn15  l=0.13u w=0.34u m=1
M9 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M13 Y B N_13 VDD mp15  l=0.13u w=0.69u m=1
M14 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M16 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
.ends nr02d4
* SPICE INPUT		Tue Jul 31 19:53:50 2018	nr02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02dm
.subckt nr02dm Y GND VDD B A
M1 GND B Y GND mn15  l=0.13u w=0.27u m=1
M2 GND A Y GND mn15  l=0.13u w=0.27u m=1
M3 Y B N_8 VDD mp15  l=0.13u w=0.55u m=1
M4 VDD A N_8 VDD mp15  l=0.13u w=0.55u m=1
.ends nr02dm
* SPICE INPUT		Tue Jul 31 19:54:03 2018	nr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d0
.subckt nr03d0 GND Y VDD C B A
M1 Y C GND GND mn15  l=0.13u w=0.26u m=1
M2 Y B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y C N_16 VDD mp15  l=0.13u w=0.4u m=1
M5 N_17 B N_16 VDD mp15  l=0.13u w=0.4u m=1
M6 N_17 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends nr03d0
* SPICE INPUT		Tue Jul 31 19:54:17 2018	nr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d1
.subckt nr03d1 Y VDD GND C B A
M1 Y C GND GND mn15  l=0.13u w=0.29u m=1
M2 Y B GND GND mn15  l=0.13u w=0.29u m=1
M3 Y A GND GND mn15  l=0.13u w=0.29u m=1
M4 Y C N_4 VDD mp15  l=0.13u w=0.69u m=1
M5 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M6 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nr03d1
* SPICE INPUT		Tue Jul 31 19:54:29 2018	nr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d2
.subckt nr03d2 Y VDD GND C B A
M1 Y A GND GND mn15  l=0.13u w=0.29u m=1
M2 Y A GND GND mn15  l=0.13u w=0.29u m=1
M3 GND B Y GND mn15  l=0.13u w=0.29u m=1
M4 Y C GND GND mn15  l=0.13u w=0.29u m=1
M5 Y B GND GND mn15  l=0.13u w=0.29u m=1
M6 GND C Y GND mn15  l=0.13u w=0.29u m=1
M7 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_12 B N_9 VDD mp15  l=0.13u w=0.69u m=1
M10 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M12 Y C N_9 VDD mp15  l=0.13u w=0.69u m=1
.ends nr03d2
* SPICE INPUT		Tue Jul 31 19:54:42 2018	nr03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d4
.subckt nr03d4 Y GND VDD C B A
M1 GND A Y GND mn15  l=0.13u w=0.29u m=1
M2 GND A Y GND mn15  l=0.13u w=0.29u m=1
M3 GND A Y GND mn15  l=0.13u w=0.29u m=1
M4 Y A GND GND mn15  l=0.13u w=0.29u m=1
M5 GND C Y GND mn15  l=0.13u w=0.29u m=1
M6 GND C Y GND mn15  l=0.13u w=0.29u m=1
M7 GND C Y GND mn15  l=0.13u w=0.29u m=1
M8 Y C GND GND mn15  l=0.13u w=0.29u m=1
M9 GND B Y GND mn15  l=0.13u w=0.29u m=1
M10 Y B GND GND mn15  l=0.13u w=0.29u m=1
M11 GND B Y GND mn15  l=0.13u w=0.29u m=1
M12 Y B GND GND mn15  l=0.13u w=0.29u m=1
M13 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_18 C Y VDD mp15  l=0.13u w=0.69u m=1
M18 N_18 C Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_18 C Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y C N_18 VDD mp15  l=0.13u w=0.69u m=1
M21 N_18 B N_20 VDD mp15  l=0.13u w=0.69u m=1
M22 N_20 B N_18 VDD mp15  l=0.13u w=0.69u m=1
M23 N_18 B N_20 VDD mp15  l=0.13u w=0.69u m=1
M24 N_20 B N_18 VDD mp15  l=0.13u w=0.69u m=1
.ends nr03d4
* SPICE INPUT		Tue Jul 31 19:54:55 2018	nr04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d0
.subckt nr04d0 GND Y VDD D C B A
M1 Y A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y D GND GND mn15  l=0.13u w=0.26u m=1
M4 Y C GND GND mn15  l=0.13u w=0.26u m=1
M5 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_14 B N_13 VDD mp15  l=0.13u w=0.4u m=1
M7 Y D N_12 VDD mp15  l=0.13u w=0.4u m=1
M8 N_14 C N_12 VDD mp15  l=0.13u w=0.4u m=1
.ends nr04d0
* SPICE INPUT		Tue Jul 31 19:55:08 2018	nr04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d1
.subckt nr04d1 Y VDD GND D C B A
M1 GND D Y GND mn15  l=0.13u w=0.28u m=1
M2 Y A GND GND mn15  l=0.13u w=0.28u m=1
M3 GND B Y GND mn15  l=0.13u w=0.28u m=1
M4 GND C Y GND mn15  l=0.13u w=0.28u m=1
M5 Y D N_4 VDD mp15  l=0.13u w=0.69u m=1
M6 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_6 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_6 C N_4 VDD mp15  l=0.13u w=0.69u m=1
.ends nr04d1
* SPICE INPUT		Tue Jul 31 19:55:21 2018	nr04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d2
.subckt nr04d2 GND Y VDD D C B A
M1 Y D GND GND mn15  l=0.13u w=0.28u m=1
M2 GND D Y GND mn15  l=0.13u w=0.28u m=1
M3 Y C GND GND mn15  l=0.13u w=0.28u m=1
M4 Y C GND GND mn15  l=0.13u w=0.28u m=1
M5 Y B GND GND mn15  l=0.13u w=0.28u m=1
M6 Y B GND GND mn15  l=0.13u w=0.28u m=1
M7 Y A GND GND mn15  l=0.13u w=0.28u m=1
M8 Y A GND GND mn15  l=0.13u w=0.28u m=1
M9 N_16 B N_15 VDD mp15  l=0.13u w=0.69u m=1
M10 N_16 B N_15 VDD mp15  l=0.13u w=0.69u m=1
M11 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M13 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_12 C N_15 VDD mp15  l=0.13u w=0.69u m=1
M16 N_15 C N_12 VDD mp15  l=0.13u w=0.69u m=1
.ends nr04d2
* SPICE INPUT		Tue Jul 31 19:55:34 2018	nr04d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d4
.subckt nr04d4 VDD Y GND D C B A
M1 Y B GND GND mn15  l=0.13u w=0.28u m=1
M2 Y B GND GND mn15  l=0.13u w=0.28u m=1
M3 Y B GND GND mn15  l=0.13u w=0.28u m=1
M4 Y B GND GND mn15  l=0.13u w=0.28u m=1
M5 Y C GND GND mn15  l=0.13u w=0.28u m=1
M6 Y C GND GND mn15  l=0.13u w=0.28u m=1
M7 Y C GND GND mn15  l=0.13u w=0.28u m=1
M8 Y C GND GND mn15  l=0.13u w=0.28u m=1
M9 Y D GND GND mn15  l=0.13u w=0.28u m=1
M10 GND D Y GND mn15  l=0.13u w=0.28u m=1
M11 Y D GND GND mn15  l=0.13u w=0.28u m=1
M12 Y D GND GND mn15  l=0.13u w=0.28u m=1
M13 Y A GND GND mn15  l=0.13u w=0.28u m=1
M14 Y A GND GND mn15  l=0.13u w=0.28u m=1
M15 Y A GND GND mn15  l=0.13u w=0.28u m=1
M16 Y A GND GND mn15  l=0.13u w=0.28u m=1
M17 N_3 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M18 N_3 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M19 N_3 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M20 N_2 B N_3 VDD mp15  l=0.13u w=0.69u m=1
M21 N_3 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD A N_3 VDD mp15  l=0.13u w=0.69u m=1
M23 N_3 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 VDD A N_3 VDD mp15  l=0.13u w=0.69u m=1
M25 N_12 C N_2 VDD mp15  l=0.13u w=0.69u m=1
M26 N_2 C N_12 VDD mp15  l=0.13u w=0.69u m=1
M27 N_12 C N_2 VDD mp15  l=0.13u w=0.69u m=1
M28 N_2 C N_12 VDD mp15  l=0.13u w=0.69u m=1
M29 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M31 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y D N_12 VDD mp15  l=0.13u w=0.69u m=1
.ends nr04d4
* SPICE INPUT		Tue Jul 31 19:55:46 2018	nr12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d0
.subckt nr12d0 Y VDD GND B AN
M1 GND N_3 Y GND mn15  l=0.13u w=0.26u m=1
M2 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M3 GND B Y GND mn15  l=0.13u w=0.26u m=1
M4 VDD N_3 N_5 VDD mp15  l=0.13u w=0.4u m=1
M5 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
M6 Y B N_5 VDD mp15  l=0.13u w=0.4u m=1
.ends nr12d0
* SPICE INPUT		Tue Jul 31 19:55:59 2018	nr12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d1
.subckt nr12d1 Y VDD GND B AN
M1 GND N_3 Y GND mn15  l=0.13u w=0.34u m=1
M2 GND B Y GND mn15  l=0.13u w=0.34u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.28u m=1
M4 VDD N_3 N_5 VDD mp15  l=0.13u w=0.69u m=1
M5 Y B N_5 VDD mp15  l=0.13u w=0.69u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.42u m=1
.ends nr12d1
* SPICE INPUT		Tue Jul 31 19:56:11 2018	nr12d1p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d1p5
.subckt nr12d1p5 Y VDD GND B AN
M1 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND B Y GND mn15  l=0.13u w=0.46u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.42u m=1
M4 VDD N_3 N_5 VDD mp15  l=0.13u w=0.69u m=1
M5 Y B N_5 VDD mp15  l=0.13u w=0.69u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.52u m=1
.ends nr12d1p5
* SPICE INPUT		Tue Jul 31 19:56:24 2018	nr12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d2
.subckt nr12d2 VDD Y GND B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.34u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.34u m=1
M3 GND B Y GND mn15  l=0.13u w=0.34u m=1
M4 Y B GND GND mn15  l=0.13u w=0.34u m=1
M5 Y N_3 GND GND mn15  l=0.13u w=0.34u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.52u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y B N_6 VDD mp15  l=0.13u w=0.69u m=1
M9 Y B N_7 VDD mp15  l=0.13u w=0.69u m=1
M10 N_6 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nr12d2
* SPICE INPUT		Tue Jul 31 19:56:37 2018	nr12d2p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d2p5
.subckt nr12d2p5 VDD Y GND B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.46u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND B Y GND mn15  l=0.13u w=0.46u m=1
M4 Y B GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.69u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y B N_6 VDD mp15  l=0.13u w=0.69u m=1
M9 Y B N_7 VDD mp15  l=0.13u w=0.69u m=1
M10 N_6 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nr12d2p5
* SPICE INPUT		Tue Jul 31 19:56:51 2018	nr12d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d4
.subckt nr12d4 Y GND VDD B AN
M1 GND B Y GND mn15  l=0.13u w=0.34u m=1
M2 GND B Y GND mn15  l=0.13u w=0.34u m=1
M3 GND B Y GND mn15  l=0.13u w=0.34u m=1
M4 Y B GND GND mn15  l=0.13u w=0.34u m=1
M5 N_5 AN GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.34u m=1
M7 Y N_5 GND GND mn15  l=0.13u w=0.34u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.34u m=1
M9 Y N_5 GND GND mn15  l=0.13u w=0.34u m=1
M10 VDD AN N_5 VDD mp15  l=0.13u w=0.69u m=1
M11 Y B N_14 VDD mp15  l=0.13u w=0.69u m=1
M12 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M13 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_14 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
M17 N_14 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
.ends nr12d4
* SPICE INPUT		Tue Jul 31 19:57:05 2018	nr12dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12dm
.subckt nr12dm Y VDD GND B AN
M1 GND N_3 Y GND mn15  l=0.13u w=0.27u m=1
M2 GND B Y GND mn15  l=0.13u w=0.27u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M4 VDD N_3 N_5 VDD mp15  l=0.13u w=0.55u m=1
M5 Y B N_5 VDD mp15  l=0.13u w=0.55u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
.ends nr12dm
* SPICE INPUT		Tue Jul 31 19:57:18 2018	nr13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d0
.subckt nr13d0 Y VDD GND C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 Y B GND GND mn15  l=0.13u w=0.26u m=1
M4 Y C GND GND mn15  l=0.13u w=0.26u m=1
M5 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
M6 N_8 N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_8 B N_7 VDD mp15  l=0.13u w=0.4u m=1
M8 Y C N_7 VDD mp15  l=0.13u w=0.4u m=1
.ends nr13d0
* SPICE INPUT		Tue Jul 31 19:57:31 2018	nr13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d1
.subckt nr13d1 Y VDD GND C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.28u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.29u m=1
M3 Y B GND GND mn15  l=0.13u w=0.29u m=1
M4 Y C GND GND mn15  l=0.13u w=0.29u m=1
M5 VDD AN N_3 VDD mp15  l=0.13u w=0.42u m=1
M6 N_8 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_8 B N_7 VDD mp15  l=0.13u w=0.69u m=1
M8 Y C N_7 VDD mp15  l=0.13u w=0.69u m=1
.ends nr13d1
* SPICE INPUT		Tue Jul 31 19:57:44 2018	nr13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d2
.subckt nr13d2 Y GND VDD C B AN
M1 Y B GND GND mn15  l=0.13u w=0.29u m=1
M2 Y B GND GND mn15  l=0.13u w=0.29u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.29u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.29u m=1
M5 N_5 AN GND GND mn15  l=0.13u w=0.33u m=1
M6 GND C Y GND mn15  l=0.13u w=0.29u m=1
M7 GND C Y GND mn15  l=0.13u w=0.29u m=1
M8 N_12 B N_14 VDD mp15  l=0.13u w=0.69u m=1
M9 N_14 B N_12 VDD mp15  l=0.13u w=0.69u m=1
M10 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD AN N_5 VDD mp15  l=0.13u w=0.5u m=1
.ends nr13d2
* SPICE INPUT		Tue Jul 31 19:57:57 2018	nr13d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d4
.subckt nr13d4 Y GND VDD C B AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.29u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.29u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.29u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.29u m=1
M6 GND C Y GND mn15  l=0.13u w=0.29u m=1
M7 GND C Y GND mn15  l=0.13u w=0.29u m=1
M8 GND C Y GND mn15  l=0.13u w=0.29u m=1
M9 Y C GND GND mn15  l=0.13u w=0.29u m=1
M10 GND B Y GND mn15  l=0.13u w=0.29u m=1
M11 Y B GND GND mn15  l=0.13u w=0.29u m=1
M12 GND B Y GND mn15  l=0.13u w=0.29u m=1
M13 Y B GND GND mn15  l=0.13u w=0.29u m=1
M14 VDD AN N_5 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_5 N_21 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_5 N_21 VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_5 N_21 VDD mp15  l=0.13u w=0.69u m=1
M18 N_21 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 Y C N_19 VDD mp15  l=0.13u w=0.69u m=1
M20 N_19 C Y VDD mp15  l=0.13u w=0.69u m=1
M21 N_19 C Y VDD mp15  l=0.13u w=0.69u m=1
M22 N_19 C Y VDD mp15  l=0.13u w=0.69u m=1
M23 N_19 B N_21 VDD mp15  l=0.13u w=0.69u m=1
M24 N_21 B N_19 VDD mp15  l=0.13u w=0.69u m=1
M25 N_19 B N_21 VDD mp15  l=0.13u w=0.69u m=1
M26 N_21 B N_19 VDD mp15  l=0.13u w=0.69u m=1
.ends nr13d4
* SPICE INPUT		Tue Jul 31 19:58:10 2018	nr14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d0
.subckt nr14d0 Y VDD GND D C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND B Y GND mn15  l=0.13u w=0.26u m=1
M4 GND D Y GND mn15  l=0.13u w=0.26u m=1
M5 GND C Y GND mn15  l=0.13u w=0.26u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
M7 N_9 N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_10 B N_9 VDD mp15  l=0.13u w=0.4u m=1
M9 Y D N_8 VDD mp15  l=0.13u w=0.4u m=1
M10 N_10 C N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends nr14d0
* SPICE INPUT		Tue Jul 31 19:58:23 2018	nr14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d1
.subckt nr14d1 Y VDD GND D C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.28u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M3 GND B Y GND mn15  l=0.13u w=0.28u m=1
M4 GND D Y GND mn15  l=0.13u w=0.28u m=1
M5 GND C Y GND mn15  l=0.13u w=0.28u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.42u m=1
M7 N_9 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_10 B N_9 VDD mp15  l=0.13u w=0.69u m=1
M9 Y D N_8 VDD mp15  l=0.13u w=0.69u m=1
M10 N_10 C N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends nr14d1
* SPICE INPUT		Tue Jul 31 19:58:36 2018	nr14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d2
.subckt nr14d2 GND Y VDD D C B AN
M1 Y D GND GND mn15  l=0.13u w=0.28u m=1
M2 GND D Y GND mn15  l=0.13u w=0.28u m=1
M3 Y C GND GND mn15  l=0.13u w=0.28u m=1
M4 Y C GND GND mn15  l=0.13u w=0.28u m=1
M5 Y N_12 GND GND mn15  l=0.13u w=0.28u m=1
M6 Y N_12 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y B GND GND mn15  l=0.13u w=0.28u m=1
M8 Y B GND GND mn15  l=0.13u w=0.28u m=1
M9 N_12 AN GND GND mn15  l=0.13u w=0.33u m=1
M10 N_12 AN VDD VDD mp15  l=0.13u w=0.5u m=1
M11 N_18 N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_12 N_18 VDD mp15  l=0.13u w=0.69u m=1
M13 N_18 B N_17 VDD mp15  l=0.13u w=0.69u m=1
M14 N_18 B N_17 VDD mp15  l=0.13u w=0.69u m=1
M15 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M16 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M17 N_14 C N_17 VDD mp15  l=0.13u w=0.69u m=1
M18 N_17 C N_14 VDD mp15  l=0.13u w=0.69u m=1
.ends nr14d2
* SPICE INPUT		Tue Jul 31 19:58:49 2018	nr14d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d4
.subckt nr14d4 VDD Y GND D C B AN
M1 N_2 AN GND GND mn15  l=0.13u w=0.46u m=1
M2 Y N_2 GND GND mn15  l=0.13u w=0.28u m=1
M3 Y N_2 GND GND mn15  l=0.13u w=0.28u m=1
M4 Y N_2 GND GND mn15  l=0.13u w=0.28u m=1
M5 Y N_2 GND GND mn15  l=0.13u w=0.28u m=1
M6 Y B GND GND mn15  l=0.13u w=0.28u m=1
M7 Y B GND GND mn15  l=0.13u w=0.28u m=1
M8 Y B GND GND mn15  l=0.13u w=0.28u m=1
M9 Y B GND GND mn15  l=0.13u w=0.28u m=1
M10 Y C GND GND mn15  l=0.13u w=0.28u m=1
M11 Y C GND GND mn15  l=0.13u w=0.28u m=1
M12 Y C GND GND mn15  l=0.13u w=0.28u m=1
M13 Y C GND GND mn15  l=0.13u w=0.28u m=1
M14 Y D GND GND mn15  l=0.13u w=0.28u m=1
M15 GND D Y GND mn15  l=0.13u w=0.28u m=1
M16 Y D GND GND mn15  l=0.13u w=0.28u m=1
M17 Y D GND GND mn15  l=0.13u w=0.28u m=1
M18 VDD AN N_2 VDD mp15  l=0.13u w=0.69u m=1
M19 N_5 N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_2 N_5 VDD mp15  l=0.13u w=0.69u m=1
M21 N_5 N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_2 N_5 VDD mp15  l=0.13u w=0.69u m=1
M23 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M24 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M25 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M26 N_4 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M27 N_14 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M28 N_4 C N_14 VDD mp15  l=0.13u w=0.69u m=1
M29 N_14 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M30 N_4 C N_14 VDD mp15  l=0.13u w=0.69u m=1
M31 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M32 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M33 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M34 Y D N_14 VDD mp15  l=0.13u w=0.69u m=1
.ends nr14d4
* SPICE INPUT		Tue Jul 31 19:59:02 2018	nr24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d0
.subckt nr24d0 GND Y VDD AN C D BN
M1 N_5 AN GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_3 Y GND mn15  l=0.13u w=0.26u m=1
M4 Y C GND GND mn15  l=0.13u w=0.26u m=1
M5 Y D GND GND mn15  l=0.13u w=0.26u m=1
M6 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M7 VDD AN N_5 VDD mp15  l=0.13u w=0.4u m=1
M8 N_15 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_16 N_3 N_15 VDD mp15  l=0.13u w=0.4u m=1
M10 N_16 C N_14 VDD mp15  l=0.13u w=0.4u m=1
M11 N_14 D Y VDD mp15  l=0.13u w=0.4u m=1
M12 VDD BN N_3 VDD mp15  l=0.13u w=0.4u m=1
.ends nr24d0
* SPICE INPUT		Tue Jul 31 19:59:14 2018	nr24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d1
.subckt nr24d1 GND Y VDD AN C D BN
M1 N_5 AN GND GND mn15  l=0.13u w=0.28u m=1
M2 Y N_5 GND GND mn15  l=0.13u w=0.28u m=1
M3 GND N_3 Y GND mn15  l=0.13u w=0.28u m=1
M4 Y C GND GND mn15  l=0.13u w=0.28u m=1
M5 Y D GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 BN GND GND mn15  l=0.13u w=0.28u m=1
M7 VDD AN N_5 VDD mp15  l=0.13u w=0.42u m=1
M8 N_15 N_5 VDD VDD mp15  l=0.13u w=0.7u m=1
M9 N_16 N_3 N_15 VDD mp15  l=0.13u w=0.7u m=1
M10 N_16 C N_14 VDD mp15  l=0.13u w=0.7u m=1
M11 N_14 D Y VDD mp15  l=0.13u w=0.7u m=1
M12 VDD BN N_3 VDD mp15  l=0.13u w=0.42u m=1
.ends nr24d1
* SPICE INPUT		Tue Jul 31 19:59:27 2018	nr24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d2
.subckt nr24d2 GND Y VDD C BN AN D
M1 N_4 BN GND GND mn15  l=0.13u w=0.4u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.4u m=1
M3 Y D GND GND mn15  l=0.13u w=0.28u m=1
M4 GND D Y GND mn15  l=0.13u w=0.28u m=1
M5 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M8 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M9 Y C GND GND mn15  l=0.13u w=0.28u m=1
M10 Y C GND GND mn15  l=0.13u w=0.28u m=1
M11 N_4 BN VDD VDD mp15  l=0.13u w=0.6u m=1
M12 N_3 AN VDD VDD mp15  l=0.13u w=0.6u m=1
M13 N_21 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_3 N_21 VDD mp15  l=0.13u w=0.69u m=1
M15 N_21 N_4 N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_21 N_4 N_20 VDD mp15  l=0.13u w=0.69u m=1
M17 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M18 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_19 C N_20 VDD mp15  l=0.13u w=0.69u m=1
M20 N_20 C N_19 VDD mp15  l=0.13u w=0.69u m=1
.ends nr24d2
* SPICE INPUT		Tue Jul 31 19:59:40 2018	nr24d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d4
.subckt nr24d4 VDD Y GND D C AN BN
M1 N_4 BN GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M4 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M5 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M8 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M10 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M11 Y C GND GND mn15  l=0.13u w=0.28u m=1
M12 Y C GND GND mn15  l=0.13u w=0.28u m=1
M13 Y C GND GND mn15  l=0.13u w=0.28u m=1
M14 Y C GND GND mn15  l=0.13u w=0.28u m=1
M15 Y D GND GND mn15  l=0.13u w=0.28u m=1
M16 GND D Y GND mn15  l=0.13u w=0.28u m=1
M17 Y D GND GND mn15  l=0.13u w=0.28u m=1
M18 Y D GND GND mn15  l=0.13u w=0.28u m=1
M19 N_4 BN VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_3 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_6 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_3 N_6 VDD mp15  l=0.13u w=0.69u m=1
M23 N_6 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_3 N_6 VDD mp15  l=0.13u w=0.69u m=1
M25 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.69u m=1
M26 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.69u m=1
M27 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.69u m=1
M28 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.69u m=1
M29 N_15 C N_5 VDD mp15  l=0.13u w=0.69u m=1
M30 N_5 C N_15 VDD mp15  l=0.13u w=0.69u m=1
M31 N_15 C N_5 VDD mp15  l=0.13u w=0.69u m=1
M32 N_5 C N_15 VDD mp15  l=0.13u w=0.69u m=1
M33 N_15 D Y VDD mp15  l=0.13u w=0.69u m=1
M34 N_15 D Y VDD mp15  l=0.13u w=0.69u m=1
M35 N_15 D Y VDD mp15  l=0.13u w=0.69u m=1
M36 Y D N_15 VDD mp15  l=0.13u w=0.69u m=1
.ends nr24d4
* SPICE INPUT		Tue Jul 31 19:59:53 2018	oai211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d0
.subckt oai211d0 Y GND VDD D C B A
M1 N_4 C N_6 GND mn15  l=0.13u w=0.26u m=1
M2 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M3 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_6 D Y GND mn15  l=0.13u w=0.26u m=1
M5 Y C VDD VDD mp15  l=0.13u w=0.27u m=1
M6 N_13 B Y VDD mp15  l=0.13u w=0.4u m=1
M7 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 Y D VDD VDD mp15  l=0.13u w=0.27u m=1
.ends oai211d0
* SPICE INPUT		Tue Jul 31 20:00:06 2018	oai211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d1
.subckt oai211d1 Y GND VDD D C B A
M1 N_4 C N_6 GND mn15  l=0.13u w=0.46u m=1
M2 N_4 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M4 Y D N_6 GND mn15  l=0.13u w=0.46u m=1
M5 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M6 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M7 N_14 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oai211d1
* SPICE INPUT		Tue Jul 31 20:00:19 2018	oai211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d2
.subckt oai211d2 GND Y B A D C VDD
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_2 C N_9 GND mn15  l=0.13u w=0.46u m=1
M6 Y D N_9 GND mn15  l=0.13u w=0.46u m=1
M7 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_10 C N_2 GND mn15  l=0.13u w=0.46u m=1
M9 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_21 B Y VDD mp15  l=0.13u w=0.69u m=1
M11 Y B N_20 VDD mp15  l=0.13u w=0.69u m=1
M12 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M14 VDD D Y VDD mp15  l=0.13u w=0.48u m=1
M15 VDD D Y VDD mp15  l=0.13u w=0.48u m=1
M16 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
.ends oai211d2
* SPICE INPUT		Tue Jul 31 20:00:33 2018	oai211d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d4
.subckt oai211d4 GND VDD D Y C A B
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_10 B GND GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_10 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_10 GND mn15  l=0.13u w=0.46u m=1
M7 GND B N_10 GND mn15  l=0.13u w=0.46u m=1
M8 GND B N_10 GND mn15  l=0.13u w=0.46u m=1
M9 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M10 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M11 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M12 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M13 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M14 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M15 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M16 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M17 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_16 B Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_15 B Y VDD mp15  l=0.13u w=0.69u m=1
M20 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M23 VDD D Y VDD mp15  l=0.13u w=0.46u m=1
M24 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M25 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M26 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M28 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M29 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M30 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M31 N_18 B Y VDD mp15  l=0.13u w=0.69u m=1
M32 N_17 B Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai211d4
* SPICE INPUT		Tue Jul 31 20:00:46 2018	oai21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d0
.subckt oai21d0 Y GND VDD C B A
M1 GND A N_2 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.26u m=1
M3 Y C N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_20 A VDD VDD mp15  l=0.13u w=0.4u m=1
M5 N_20 B Y VDD mp15  l=0.13u w=0.4u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.27u m=1
.ends oai21d0
* SPICE INPUT		Tue Jul 31 20:00:59 2018	oai21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d1
.subckt oai21d1 Y GND VDD C B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 Y C N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M5 N_20 B Y VDD mp15  l=0.13u w=0.69u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oai21d1
* SPICE INPUT		Tue Jul 31 20:01:12 2018	oai21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d2
.subckt oai21d2 Y VDD GND C A B
M1 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 C Y GND mn15  l=0.13u w=0.46u m=1
M3 N_12 C Y GND mn15  l=0.13u w=0.46u m=1
M4 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND B N_12 GND mn15  l=0.13u w=0.46u m=1
M6 N_12 B GND GND mn15  l=0.13u w=0.46u m=1
M7 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 VDD C Y VDD mp15  l=0.13u w=0.46u m=1
M9 VDD C Y VDD mp15  l=0.13u w=0.46u m=1
M10 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 B Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y B N_7 VDD mp15  l=0.13u w=0.69u m=1
.ends oai21d2
* SPICE INPUT		Tue Jul 31 20:01:25 2018	oai21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d4
.subckt oai21d4 Y VDD GND C A B
M1 GND A N_20 GND mn15  l=0.13u w=0.46u m=1
M2 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M7 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M8 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M10 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M11 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M12 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M13 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M17 Y B N_13 VDD mp15  l=0.13u w=0.69u m=1
M18 N_12 B Y VDD mp15  l=0.13u w=0.69u m=1
M19 Y B N_11 VDD mp15  l=0.13u w=0.69u m=1
M20 N_14 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD C Y VDD mp15  l=0.13u w=0.46u m=1
M22 VDD C Y VDD mp15  l=0.13u w=0.46u m=1
M23 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M24 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oai21d4
* SPICE INPUT		Tue Jul 31 20:01:38 2018	oai21dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21dm
.subckt oai21dm Y GND VDD C B A
M1 GND B N_2 GND mn15  l=0.13u w=0.36u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.36u m=1
M3 Y C N_2 GND mn15  l=0.13u w=0.36u m=1
M4 N_20 B Y VDD mp15  l=0.13u w=0.55u m=1
M5 N_20 A VDD VDD mp15  l=0.13u w=0.55u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.37u m=1
.ends oai21dm
* SPICE INPUT		Tue Jul 31 20:01:51 2018	oai21md0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21md0
.subckt oai21md0 VDD Y B CN GND A
M1 N_3 CN GND GND mn15  l=0.13u w=0.26u m=1
M2 GND A N_9 GND mn15  l=0.13u w=0.26u m=1
M3 GND B N_9 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_3 N_9 GND mn15  l=0.13u w=0.26u m=1
M5 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_6 B Y VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_3 VDD VDD mp15  l=0.13u w=0.27u m=1
M8 N_3 CN VDD VDD mp15  l=0.13u w=0.4u m=1
.ends oai21md0
* SPICE INPUT		Tue Jul 31 20:02:04 2018	oai21md1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21md1
.subckt oai21md1 Y VDD GND CN B A
M1 GND A N_11 GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M3 Y N_5 N_11 GND mn15  l=0.13u w=0.46u m=1
M4 GND CN N_5 GND mn15  l=0.13u w=0.26u m=1
M5 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 N_7 B Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD N_5 Y VDD mp15  l=0.13u w=0.46u m=1
M8 VDD CN N_5 VDD mp15  l=0.13u w=0.4u m=1
.ends oai21md1
* SPICE INPUT		Tue Jul 31 20:02:18 2018	oai21md2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21md2
.subckt oai21md2 Y GND VDD CN B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_9 N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_2 N_9 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND CN N_9 GND mn15  l=0.13u w=0.3u m=1
M8 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M9 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_9 VDD VDD mp15  l=0.13u w=0.46u m=1
M13 Y N_9 VDD VDD mp15  l=0.13u w=0.46u m=1
M14 N_9 CN VDD VDD mp15  l=0.13u w=0.43u m=1
.ends oai21md2
* SPICE INPUT		Tue Jul 31 20:02:31 2018	oai21md4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21md4
.subckt oai21md4 Y GND VDD CN B A
M1 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 N_15 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_3 N_15 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_3 N_15 Y GND mn15  l=0.13u w=0.46u m=1
M8 N_3 N_15 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M10 GND B N_3 GND mn15  l=0.13u w=0.46u m=1
M11 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M12 GND B N_3 GND mn15  l=0.13u w=0.46u m=1
M13 GND CN N_15 GND mn15  l=0.13u w=0.46u m=1
M14 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_15 VDD VDD mp15  l=0.13u w=0.46u m=1
M19 VDD N_15 Y VDD mp15  l=0.13u w=0.46u m=1
M20 Y N_15 VDD VDD mp15  l=0.13u w=0.46u m=1
M21 Y N_15 VDD VDD mp15  l=0.13u w=0.46u m=1
M22 Y B N_20 VDD mp15  l=0.13u w=0.55u m=1
M23 N_20 B Y VDD mp15  l=0.13u w=0.55u m=1
M24 Y B N_20 VDD mp15  l=0.13u w=0.55u m=1
M25 Y B N_20 VDD mp15  l=0.13u w=0.55u m=1
M26 Y B N_20 VDD mp15  l=0.13u w=0.56u m=1
M27 VDD CN N_15 VDD mp15  l=0.13u w=0.69u m=1
.ends oai21md4
* SPICE INPUT		Tue Jul 31 20:02:44 2018	oai221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d0
.subckt oai221d0 VDD Y GND E C D B A
M1 GND B N_14 GND mn15  l=0.13u w=0.26u m=1
M2 GND A N_14 GND mn15  l=0.13u w=0.26u m=1
M3 N_13 D N_14 GND mn15  l=0.13u w=0.26u m=1
M4 N_14 C N_13 GND mn15  l=0.13u w=0.26u m=1
M5 Y E N_13 GND mn15  l=0.13u w=0.26u m=1
M6 Y B N_8 VDD mp15  l=0.13u w=0.4u m=1
M7 Y D N_7 VDD mp15  l=0.13u w=0.4u m=1
M8 N_7 C VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y E VDD VDD mp15  l=0.13u w=0.27u m=1
.ends oai221d0
* SPICE INPUT		Tue Jul 31 20:02:57 2018	oai221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d1
.subckt oai221d1 GND Y VDD E C D B A
M1 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 Y E N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 C N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_5 D N_2 GND mn15  l=0.13u w=0.46u m=1
M6 Y B N_18 VDD mp15  l=0.13u w=0.69u m=1
M7 N_17 C VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y D N_17 VDD mp15  l=0.13u w=0.69u m=1
M9 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y E VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oai221d1
* SPICE INPUT		Tue Jul 31 20:03:10 2018	oai221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d2
.subckt oai221d2 Y VDD GND E C D A B
M1 N_20 C N_22 GND mn15  l=0.13u w=0.46u m=1
M2 N_20 D N_22 GND mn15  l=0.13u w=0.46u m=1
M3 N_20 D N_22 GND mn15  l=0.13u w=0.46u m=1
M4 N_20 C N_22 GND mn15  l=0.13u w=0.46u m=1
M5 N_20 E Y GND mn15  l=0.13u w=0.46u m=1
M6 N_20 E Y GND mn15  l=0.13u w=0.46u m=1
M7 GND B N_22 GND mn15  l=0.13u w=0.46u m=1
M8 N_22 B GND GND mn15  l=0.13u w=0.46u m=1
M9 GND A N_22 GND mn15  l=0.13u w=0.46u m=1
M10 N_22 A GND GND mn15  l=0.13u w=0.46u m=1
M11 N_11 C VDD VDD mp15  l=0.13u w=0.595u m=1
M12 N_11 D Y VDD mp15  l=0.13u w=0.595u m=1
M13 Y D N_10 VDD mp15  l=0.13u w=0.595u m=1
M14 N_10 C VDD VDD mp15  l=0.13u w=0.595u m=1
M15 VDD E Y VDD mp15  l=0.13u w=0.46u m=1
M16 VDD E Y VDD mp15  l=0.13u w=0.46u m=1
M17 Y B N_12 VDD mp15  l=0.13u w=0.69u m=1
M18 Y B N_13 VDD mp15  l=0.13u w=0.69u m=1
M19 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends oai221d2
* SPICE INPUT		Tue Jul 31 20:03:23 2018	oai221d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d4
.subckt oai221d4 Y D C A B GND VDD E
M1 N_10 C N_11 GND mn15  l=0.13u w=0.46u m=1
M2 N_10 C N_11 GND mn15  l=0.13u w=0.46u m=1
M3 N_10 C N_11 GND mn15  l=0.13u w=0.46u m=1
M4 N_10 D N_11 GND mn15  l=0.13u w=0.46u m=1
M5 N_10 D N_11 GND mn15  l=0.13u w=0.46u m=1
M6 N_10 D N_11 GND mn15  l=0.13u w=0.46u m=1
M7 N_10 D N_11 GND mn15  l=0.13u w=0.46u m=1
M8 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M9 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M10 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M11 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M12 N_10 C N_11 GND mn15  l=0.13u w=0.46u m=1
M13 N_11 B GND GND mn15  l=0.13u w=0.46u m=1
M14 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M15 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M16 GND A N_11 GND mn15  l=0.13u w=0.46u m=1
M17 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M18 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M19 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M20 GND A N_11 GND mn15  l=0.13u w=0.46u m=1
M21 N_21 B Y VDD mp15  l=0.13u w=0.69u m=1
M22 N_20 B Y VDD mp15  l=0.13u w=0.69u m=1
M23 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_22 B Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_23 B Y VDD mp15  l=0.13u w=0.69u m=1
M28 N_24 C VDD VDD mp15  l=0.13u w=0.595u m=1
M29 N_24 D Y VDD mp15  l=0.13u w=0.595u m=1
M30 N_23 A VDD VDD mp15  l=0.13u w=0.69u m=1
M31 N_26 C VDD VDD mp15  l=0.13u w=0.595u m=1
M32 N_25 C VDD VDD mp15  l=0.13u w=0.595u m=1
M33 N_25 D Y VDD mp15  l=0.13u w=0.595u m=1
M34 N_26 D Y VDD mp15  l=0.13u w=0.595u m=1
M35 N_27 D Y VDD mp15  l=0.13u w=0.595u m=1
M36 VDD E Y VDD mp15  l=0.13u w=0.46u m=1
M37 VDD E Y VDD mp15  l=0.13u w=0.46u m=1
M38 Y E VDD VDD mp15  l=0.13u w=0.46u m=1
M39 Y E VDD VDD mp15  l=0.13u w=0.46u m=1
M40 N_27 C VDD VDD mp15  l=0.13u w=0.595u m=1
.ends oai221d4
* SPICE INPUT		Tue Jul 31 20:03:37 2018	oai222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d0
.subckt oai222d0 Y VDD GND F E C D B A
M1 N_14 E Y GND mn15  l=0.13u w=0.26u m=1
M2 N_14 F Y GND mn15  l=0.13u w=0.26u m=1
M3 N_14 C N_16 GND mn15  l=0.13u w=0.26u m=1
M4 GND A N_16 GND mn15  l=0.13u w=0.26u m=1
M5 N_16 B GND GND mn15  l=0.13u w=0.26u m=1
M6 N_16 D N_14 GND mn15  l=0.13u w=0.26u m=1
M7 VDD C N_11 VDD mp15  l=0.13u w=0.4u m=1
M8 VDD E N_9 VDD mp15  l=0.13u w=0.4u m=1
M9 Y F N_9 VDD mp15  l=0.13u w=0.4u m=1
M10 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M11 Y B N_10 VDD mp15  l=0.13u w=0.4u m=1
M12 N_11 D Y VDD mp15  l=0.13u w=0.4u m=1
.ends oai222d0
* SPICE INPUT		Tue Jul 31 20:03:50 2018	oai222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d1
.subckt oai222d1 GND Y VDD E F C D B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 D N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M5 Y E N_3 GND mn15  l=0.13u w=0.46u m=1
M6 Y F N_3 GND mn15  l=0.13u w=0.46u m=1
M7 VDD E N_21 VDD mp15  l=0.13u w=0.69u m=1
M8 Y F N_21 VDD mp15  l=0.13u w=0.69u m=1
M9 N_23 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_23 B Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_24 D Y VDD mp15  l=0.13u w=0.36u m=1
M12 VDD C N_24 VDD mp15  l=0.13u w=0.36u m=1
M13 VDD C N_22 VDD mp15  l=0.13u w=0.35u m=1
M14 Y D N_22 VDD mp15  l=0.13u w=0.35u m=1
.ends oai222d1
* SPICE INPUT		Tue Jul 31 20:04:02 2018	oai222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d2
.subckt oai222d2 Y GND VDD A B D F E C
M1 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M2 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M3 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M4 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_7 C N_3 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 D N_7 GND mn15  l=0.13u w=0.46u m=1
M8 N_3 D N_7 GND mn15  l=0.13u w=0.46u m=1
M9 N_7 B GND GND mn15  l=0.13u w=0.46u m=1
M10 GND A N_7 GND mn15  l=0.13u w=0.46u m=1
M11 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M12 N_7 B GND GND mn15  l=0.13u w=0.46u m=1
M13 N_21 E VDD VDD mp15  l=0.13u w=0.46u m=1
M14 N_21 E VDD VDD mp15  l=0.13u w=0.46u m=1
M15 N_21 E VDD VDD mp15  l=0.13u w=0.46u m=1
M16 N_20 C VDD VDD mp15  l=0.13u w=0.46u m=1
M17 VDD C N_20 VDD mp15  l=0.13u w=0.46u m=1
M18 N_20 C VDD VDD mp15  l=0.13u w=0.46u m=1
M19 N_20 D Y VDD mp15  l=0.13u w=0.46u m=1
M20 N_20 D Y VDD mp15  l=0.13u w=0.46u m=1
M21 N_20 D Y VDD mp15  l=0.13u w=0.46u m=1
M22 N_28 B Y VDD mp15  l=0.13u w=0.69u m=1
M23 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_27 B Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_21 F Y VDD mp15  l=0.13u w=0.46u m=1
M27 Y F N_21 VDD mp15  l=0.13u w=0.46u m=1
M28 Y F N_21 VDD mp15  l=0.13u w=0.46u m=1
.ends oai222d2
* SPICE INPUT		Tue Jul 31 20:04:15 2018	oai222d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d4
.subckt oai222d4 GND Y F C VDD E A D B
M1 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 C N_3 GND mn15  l=0.13u w=0.46u m=1
M5 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M7 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M8 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M9 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M10 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M11 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M12 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M13 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M14 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M15 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M16 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M17 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M18 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M19 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M20 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M21 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M22 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M23 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M24 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M25 N_37 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD A N_37 VDD mp15  l=0.13u w=0.69u m=1
M27 N_37 A VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD A N_37 VDD mp15  l=0.13u w=0.69u m=1
M29 N_37 B Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y B N_37 VDD mp15  l=0.13u w=0.69u m=1
M31 N_37 B Y VDD mp15  l=0.13u w=0.69u m=1
M32 N_37 B Y VDD mp15  l=0.13u w=0.69u m=1
M33 Y F N_31 VDD mp15  l=0.13u w=0.565u m=1
M34 Y F N_31 VDD mp15  l=0.13u w=0.565u m=1
M35 Y F N_31 VDD mp15  l=0.13u w=0.565u m=1
M36 N_31 F Y VDD mp15  l=0.13u w=0.565u m=1
M37 Y F N_31 VDD mp15  l=0.13u w=0.5u m=1
M38 VDD C N_33 VDD mp15  l=0.13u w=0.56u m=1
M39 N_33 C VDD VDD mp15  l=0.13u w=0.55u m=1
M40 N_33 C VDD VDD mp15  l=0.13u w=0.55u m=1
M41 VDD C N_33 VDD mp15  l=0.13u w=0.55u m=1
M42 N_33 C VDD VDD mp15  l=0.13u w=0.55u m=1
M43 Y D N_33 VDD mp15  l=0.13u w=0.565u m=1
M44 Y D N_33 VDD mp15  l=0.13u w=0.565u m=1
M45 Y D N_33 VDD mp15  l=0.13u w=0.565u m=1
M46 N_33 D Y VDD mp15  l=0.13u w=0.565u m=1
M47 N_33 D Y VDD mp15  l=0.13u w=0.5u m=1
M48 N_31 E VDD VDD mp15  l=0.13u w=0.56u m=1
M49 VDD E N_31 VDD mp15  l=0.13u w=0.55u m=1
M50 N_31 E VDD VDD mp15  l=0.13u w=0.55u m=1
M51 N_31 E VDD VDD mp15  l=0.13u w=0.55u m=1
M52 N_31 E VDD VDD mp15  l=0.13u w=0.55u m=1
.ends oai222d4
* SPICE INPUT		Tue Jul 31 20:04:28 2018	oai22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d0
.subckt oai22d0 VDD Y GND A C B D
M1 N_12 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_12 D Y GND mn15  l=0.13u w=0.26u m=1
M3 N_12 B GND GND mn15  l=0.13u w=0.26u m=1
M4 N_12 C Y GND mn15  l=0.13u w=0.26u m=1
M5 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y D N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 Y B N_8 VDD mp15  l=0.13u w=0.4u m=1
M8 VDD C N_7 VDD mp15  l=0.13u w=0.4u m=1
.ends oai22d0
* SPICE INPUT		Tue Jul 31 20:04:41 2018	oai22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d1
.subckt oai22d1 VDD Y GND A C B D
M1 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 D Y GND mn15  l=0.13u w=0.46u m=1
M3 N_12 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_12 C Y GND mn15  l=0.13u w=0.46u m=1
M5 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y D N_7 VDD mp15  l=0.13u w=0.595u m=1
M7 N_8 B Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD C N_7 VDD mp15  l=0.13u w=0.595u m=1
.ends oai22d1
* SPICE INPUT		Tue Jul 31 20:04:54 2018	oai22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d2
.subckt oai22d2 VDD Y GND D A B C
M1 GND B N_20 GND mn15  l=0.13u w=0.46u m=1
M2 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M5 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M7 N_20 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_20 D Y GND mn15  l=0.13u w=0.46u m=1
M9 N_9 B Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y B N_8 VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD C N_7 VDD mp15  l=0.13u w=0.595u m=1
M13 N_9 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_10 C VDD VDD mp15  l=0.13u w=0.595u m=1
M15 Y D N_7 VDD mp15  l=0.13u w=0.595u m=1
M16 Y D N_10 VDD mp15  l=0.13u w=0.595u m=1
.ends oai22d2
* SPICE INPUT		Tue Jul 31 20:05:07 2018	oai22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d4
.subckt oai22d4 VDD Y A B D GND C
M1 GND B N_30 GND mn15  l=0.13u w=0.46u m=1
M2 N_30 B GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_30 GND mn15  l=0.13u w=0.46u m=1
M4 N_30 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_30 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_30 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_30 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_30 C Y GND mn15  l=0.13u w=0.46u m=1
M9 N_30 A GND GND mn15  l=0.13u w=0.46u m=1
M10 N_30 C Y GND mn15  l=0.13u w=0.46u m=1
M11 N_30 D Y GND mn15  l=0.13u w=0.46u m=1
M12 N_30 D Y GND mn15  l=0.13u w=0.46u m=1
M13 N_30 C Y GND mn15  l=0.13u w=0.46u m=1
M14 N_30 C Y GND mn15  l=0.13u w=0.46u m=1
M15 N_30 D Y GND mn15  l=0.13u w=0.46u m=1
M16 N_30 D Y GND mn15  l=0.13u w=0.46u m=1
M17 N_15 B Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y B N_14 VDD mp15  l=0.13u w=0.69u m=1
M19 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M21 Y B N_12 VDD mp15  l=0.13u w=0.69u m=1
M22 N_14 A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_16 C VDD VDD mp15  l=0.13u w=0.595u m=1
M25 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD C N_11 VDD mp15  l=0.13u w=0.595u m=1
M27 Y D N_11 VDD mp15  l=0.13u w=0.595u m=1
M28 Y D N_18 VDD mp15  l=0.13u w=0.595u m=1
M29 N_18 C VDD VDD mp15  l=0.13u w=0.595u m=1
M30 N_17 C VDD VDD mp15  l=0.13u w=0.595u m=1
M31 N_17 D Y VDD mp15  l=0.13u w=0.595u m=1
M32 Y D N_16 VDD mp15  l=0.13u w=0.595u m=1
.ends oai22d4
* SPICE INPUT		Tue Jul 31 20:05:20 2018	oai22dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22dm
.subckt oai22dm VDD Y GND A C B D
M1 N_12 A GND GND mn15  l=0.13u w=0.36u m=1
M2 N_12 D Y GND mn15  l=0.13u w=0.36u m=1
M3 N_12 B GND GND mn15  l=0.13u w=0.36u m=1
M4 N_12 C Y GND mn15  l=0.13u w=0.36u m=1
M5 N_8 A VDD VDD mp15  l=0.13u w=0.55u m=1
M6 Y D N_7 VDD mp15  l=0.13u w=0.55u m=1
M7 Y B N_8 VDD mp15  l=0.13u w=0.55u m=1
M8 VDD C N_7 VDD mp15  l=0.13u w=0.55u m=1
.ends oai22dm
* SPICE INPUT		Tue Jul 31 20:05:32 2018	oai2m1d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai2m1d0
.subckt oai2m1d0 VDD Y GND C A BN
M1 Y C N_11 GND mn15  l=0.13u w=0.26u m=1
M2 N_11 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND A N_11 GND mn15  l=0.13u w=0.26u m=1
M4 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M5 N_3 BN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.27u m=1
M7 N_7 N_3 Y VDD mp15  l=0.13u w=0.4u m=1
M8 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends oai2m1d0
* SPICE INPUT		Tue Jul 31 20:05:45 2018	oai2m1d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai2m1d1
.subckt oai2m1d1 GND Y VDD C A BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 Y C N_4 GND mn15  l=0.13u w=0.46u m=1
M3 N_4 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 BN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M7 N_26 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M8 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends oai2m1d1
* SPICE INPUT		Tue Jul 31 20:05:57 2018	oai2m1d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai2m1d2
.subckt oai2m1d2 GND Y VDD C A BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.46u m=1
M2 N_5 C Y GND mn15  l=0.13u w=0.46u m=1
M3 N_5 C Y GND mn15  l=0.13u w=0.46u m=1
M4 N_5 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_5 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_3 BN VDD VDD mp15  l=0.13u w=0.69u m=1
M9 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M10 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M11 N_39 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M12 N_39 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_38 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_38 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai2m1d2
* SPICE INPUT		Tue Jul 31 20:06:10 2018	oai2m1d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai2m1d4
.subckt oai2m1d4 GND Y VDD C A BN
M1 GND BN N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND BN N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M6 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M7 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M8 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M9 N_6 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_6 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_6 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M13 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M14 N_6 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M15 VDD BN N_2 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD BN N_2 VDD mp15  l=0.13u w=0.69u m=1
M17 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_29 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M20 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M21 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M22 VDD C Y VDD mp15  l=0.13u w=0.48u m=1
M23 N_29 N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M24 N_28 N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M25 N_27 N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M28 N_26 N_2 Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai2m1d4
* SPICE INPUT		Tue Jul 31 20:06:23 2018	oai31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d0
.subckt oai31d0 VDD Y GND D A B C
M1 N_11 C GND GND mn15  l=0.13u w=0.26u m=1
M2 N_11 B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y D N_11 GND mn15  l=0.13u w=0.26u m=1
M4 GND A N_11 GND mn15  l=0.13u w=0.26u m=1
M5 N_7 C Y VDD mp15  l=0.13u w=0.4u m=1
M6 N_8 B N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 Y D VDD VDD mp15  l=0.13u w=0.27u m=1
M8 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends oai31d0
* SPICE INPUT		Tue Jul 31 20:06:36 2018	oai31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d1
.subckt oai31d1 Y GND VDD D A B C
M1 Y D N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 C GND GND mn15  l=0.13u w=0.46u m=1
M5 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M6 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_15 B N_14 VDD mp15  l=0.13u w=0.69u m=1
M8 N_14 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai31d1
* SPICE INPUT		Tue Jul 31 20:06:50 2018	oai31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d2
.subckt oai31d2 Y VDD GND D A B C
M1 GND A N_17 GND mn15  l=0.13u w=0.46u m=1
M2 N_17 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_17 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_17 D Y GND mn15  l=0.13u w=0.46u m=1
M7 N_17 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_17 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_9 B N_8 VDD mp15  l=0.13u w=0.69u m=1
M11 N_9 C Y VDD mp15  l=0.13u w=0.69u m=1
M12 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
M13 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD D Y VDD mp15  l=0.13u w=0.46u m=1
M15 VDD D Y VDD mp15  l=0.13u w=0.46u m=1
M16 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends oai31d2
* SPICE INPUT		Tue Jul 31 20:07:03 2018	oai31d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d4
.subckt oai31d4 GND VDD Y D C B A
M1 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M2 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M3 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M4 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M5 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_9 B GND GND mn15  l=0.13u w=0.46u m=1
M10 N_9 B GND GND mn15  l=0.13u w=0.46u m=1
M11 N_9 B GND GND mn15  l=0.13u w=0.46u m=1
M12 N_9 B GND GND mn15  l=0.13u w=0.46u m=1
M13 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M14 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M15 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M16 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M17 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 VDD A N_11 VDD mp15  l=0.13u w=0.69u m=1
M19 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_11 VDD mp15  l=0.13u w=0.69u m=1
M21 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M22 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M23 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M24 N_10 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M25 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M26 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M27 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M28 VDD D Y VDD mp15  l=0.13u w=0.46u m=1
M29 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
M31 Y C N_10 VDD mp15  l=0.13u w=0.69u m=1
M32 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai31d4
* SPICE INPUT		Tue Jul 31 20:07:16 2018	oai32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d0
.subckt oai32d0 Y VDD GND E D A B C
M1 N_12 D Y GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_12 GND mn15  l=0.13u w=0.26u m=1
M3 N_12 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_12 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y E N_12 GND mn15  l=0.13u w=0.26u m=1
M6 VDD D N_8 VDD mp15  l=0.13u w=0.4u m=1
M7 N_10 B N_9 VDD mp15  l=0.13u w=0.4u m=1
M8 N_9 C Y VDD mp15  l=0.13u w=0.4u m=1
M9 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y E N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends oai32d0
* SPICE INPUT		Tue Jul 31 20:07:29 2018	oai32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d1
.subckt oai32d1 Y GND VDD D E A B C
M1 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M2 N_3 D Y GND mn15  l=0.13u w=0.46u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_14 D VDD VDD mp15  l=0.13u w=0.345u m=1
M7 Y E N_14 VDD mp15  l=0.13u w=0.345u m=1
M8 Y E N_17 VDD mp15  l=0.13u w=0.345u m=1
M9 N_17 D VDD VDD mp15  l=0.13u w=0.345u m=1
M10 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_16 B N_15 VDD mp15  l=0.13u w=0.69u m=1
M12 N_15 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai32d1
* SPICE INPUT		Tue Jul 31 20:07:42 2018	oai32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d2
.subckt oai32d2 Y GND VDD E D A B C
M1 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 D Y GND mn15  l=0.13u w=0.46u m=1
M6 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M7 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_3 D Y GND mn15  l=0.13u w=0.46u m=1
M9 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M10 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M11 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_27 B N_26 VDD mp15  l=0.13u w=0.69u m=1
M13 N_27 C Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_29 C Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD D N_28 VDD mp15  l=0.13u w=0.455u m=1
M16 N_32 D VDD VDD mp15  l=0.13u w=0.455u m=1
M17 N_30 B N_29 VDD mp15  l=0.13u w=0.69u m=1
M18 Y E N_28 VDD mp15  l=0.13u w=0.455u m=1
M19 N_30 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_31 D VDD VDD mp15  l=0.13u w=0.455u m=1
M21 N_32 E Y VDD mp15  l=0.13u w=0.455u m=1
M22 Y E N_31 VDD mp15  l=0.13u w=0.455u m=1
.ends oai32d2
* SPICE INPUT		Tue Jul 31 20:07:55 2018	oai32d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d4
.subckt oai32d4 D GND VDD Y E C B A
M1 N_10 B GND GND mn15  l=0.13u w=0.46u m=1
M2 N_10 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_10 B GND GND mn15  l=0.13u w=0.46u m=1
M4 GND B N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M6 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M7 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M9 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M10 N_10 C GND GND mn15  l=0.13u w=0.46u m=1
M11 N_10 C GND GND mn15  l=0.13u w=0.46u m=1
M12 N_10 C GND GND mn15  l=0.13u w=0.46u m=1
M13 GND C N_10 GND mn15  l=0.13u w=0.46u m=1
M14 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M15 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M16 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M17 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M18 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M19 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M20 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M21 N_12 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M22 N_12 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M23 N_12 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M24 N_11 B N_12 VDD mp15  l=0.13u w=0.69u m=1
M25 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M27 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M29 N_37 D VDD VDD mp15  l=0.13u w=0.47u m=1
M30 N_38 E Y VDD mp15  l=0.13u w=0.47u m=1
M31 N_39 D VDD VDD mp15  l=0.13u w=0.47u m=1
M32 VDD D N_38 VDD mp15  l=0.13u w=0.47u m=1
M33 N_41 D VDD VDD mp15  l=0.13u w=0.47u m=1
M34 VDD D N_40 VDD mp15  l=0.13u w=0.47u m=1
M35 N_11 C Y VDD mp15  l=0.13u w=0.69u m=1
M36 N_11 C Y VDD mp15  l=0.13u w=0.69u m=1
M37 Y C N_11 VDD mp15  l=0.13u w=0.69u m=1
M38 N_11 C Y VDD mp15  l=0.13u w=0.69u m=1
M39 N_40 E Y VDD mp15  l=0.13u w=0.47u m=1
M40 Y E N_39 VDD mp15  l=0.13u w=0.47u m=1
M41 Y E N_37 VDD mp15  l=0.13u w=0.47u m=1
M42 Y E N_41 VDD mp15  l=0.13u w=0.47u m=1
.ends oai32d4
* SPICE INPUT		Tue Jul 31 20:08:09 2018	oai33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d0
.subckt oai33d0 VDD Y GND D E F C B A
M1 Y D N_15 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_15 GND mn15  l=0.13u w=0.26u m=1
M3 Y E N_15 GND mn15  l=0.13u w=0.26u m=1
M4 N_15 F Y GND mn15  l=0.13u w=0.26u m=1
M5 N_15 C GND GND mn15  l=0.13u w=0.26u m=1
M6 N_15 A GND GND mn15  l=0.13u w=0.26u m=1
M7 VDD D N_9 VDD mp15  l=0.13u w=0.4u m=1
M8 N_11 B N_10 VDD mp15  l=0.13u w=0.4u m=1
M9 N_12 E N_9 VDD mp15  l=0.13u w=0.4u m=1
M10 N_12 F Y VDD mp15  l=0.13u w=0.4u m=1
M11 Y C N_11 VDD mp15  l=0.13u w=0.4u m=1
M12 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends oai33d0
* SPICE INPUT		Tue Jul 31 20:08:22 2018	oai33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d1
.subckt oai33d1 Y GND VDD D E F C B A
M1 GND C N_2 GND mn15  l=0.13u w=0.46u m=1
M2 Y F N_2 GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M5 Y D N_2 GND mn15  l=0.13u w=0.46u m=1
M6 Y E N_2 GND mn15  l=0.13u w=0.46u m=1
M7 Y C N_42 VDD mp15  l=0.13u w=0.69u m=1
M8 Y F N_13 VDD mp15  l=0.13u w=0.69u m=1
M9 N_42 B N_41 VDD mp15  l=0.13u w=0.69u m=1
M10 N_41 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 E N_12 VDD mp15  l=0.13u w=0.35u m=1
M12 N_12 E N_13 VDD mp15  l=0.13u w=0.34u m=1
M13 VDD D N_12 VDD mp15  l=0.13u w=0.69u m=1
.ends oai33d1
* SPICE INPUT		Tue Jul 31 20:08:35 2018	oai33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d2
.subckt oai33d2 Y GND VDD E F D B C A
M1 GND A N_3 GND mn15  l=0.13u w=0.35u m=1
M2 GND B N_3 GND mn15  l=0.13u w=0.34u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.35u m=1
M4 N_3 A GND GND mn15  l=0.13u w=0.34u m=1
M5 N_3 C GND GND mn15  l=0.13u w=0.35u m=1
M6 N_3 C GND GND mn15  l=0.13u w=0.34u m=1
M7 N_3 E Y GND mn15  l=0.13u w=0.35u m=1
M8 N_3 E Y GND mn15  l=0.13u w=0.34u m=1
M9 N_3 D Y GND mn15  l=0.13u w=0.34u m=1
M10 N_3 D Y GND mn15  l=0.13u w=0.35u m=1
M11 N_3 F Y GND mn15  l=0.13u w=0.34u m=1
M12 N_3 F Y GND mn15  l=0.13u w=0.35u m=1
M13 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_15 B N_27 VDD mp15  l=0.13u w=0.69u m=1
M15 N_15 B N_28 VDD mp15  l=0.13u w=0.69u m=1
M16 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_15 C Y VDD mp15  l=0.13u w=0.69u m=1
M18 N_15 C Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_23 E N_20 VDD mp15  l=0.13u w=0.46u m=1
M20 N_20 E N_23 VDD mp15  l=0.13u w=0.46u m=1
M21 N_23 E N_20 VDD mp15  l=0.13u w=0.46u m=1
M22 N_23 D VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_23 D VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_20 F Y VDD mp15  l=0.13u w=0.46u m=1
M25 N_20 F Y VDD mp15  l=0.13u w=0.46u m=1
M26 Y F N_20 VDD mp15  l=0.13u w=0.46u m=1
.ends oai33d2
* SPICE INPUT		Tue Jul 31 20:08:48 2018	oai33d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d4
.subckt oai33d4 GND F Y D C E VDD B A
M1 N_14 F Y GND mn15  l=0.13u w=0.56u m=1
M2 Y F N_14 GND mn15  l=0.13u w=0.56u m=1
M3 Y F N_14 GND mn15  l=0.13u w=0.56u m=1
M4 Y F N_14 GND mn15  l=0.13u w=0.16u m=1
M5 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_14 B GND GND mn15  l=0.13u w=0.46u m=1
M10 N_14 B GND GND mn15  l=0.13u w=0.46u m=1
M11 N_14 B GND GND mn15  l=0.13u w=0.46u m=1
M12 N_14 B GND GND mn15  l=0.13u w=0.46u m=1
M13 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M14 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M15 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M16 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M17 N_14 E Y GND mn15  l=0.13u w=0.46u m=1
M18 N_14 E Y GND mn15  l=0.13u w=0.46u m=1
M19 N_14 E Y GND mn15  l=0.13u w=0.46u m=1
M20 Y E N_14 GND mn15  l=0.13u w=0.46u m=1
M21 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M22 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M23 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M24 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M25 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M27 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M29 N_13 B N_12 VDD mp15  l=0.13u w=0.69u m=1
M30 N_12 B N_13 VDD mp15  l=0.13u w=0.69u m=1
M31 N_12 B N_13 VDD mp15  l=0.13u w=0.69u m=1
M32 N_12 B N_13 VDD mp15  l=0.13u w=0.69u m=1
M33 Y F N_15 VDD mp15  l=0.13u w=0.6u m=1
M34 Y F N_15 VDD mp15  l=0.13u w=0.6u m=1
M35 Y F N_15 VDD mp15  l=0.13u w=0.6u m=1
M36 N_15 F Y VDD mp15  l=0.13u w=0.6u m=1
M37 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
M38 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
M39 Y C N_13 VDD mp15  l=0.13u w=0.69u m=1
M40 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
M41 N_11 E N_15 VDD mp15  l=0.13u w=0.6u m=1
M42 N_15 E N_11 VDD mp15  l=0.13u w=0.6u m=1
M43 N_11 E N_15 VDD mp15  l=0.13u w=0.6u m=1
M44 N_15 E N_11 VDD mp15  l=0.13u w=0.6u m=1
M45 N_11 D VDD VDD mp15  l=0.13u w=0.6u m=1
M46 N_11 D VDD VDD mp15  l=0.13u w=0.6u m=1
M47 N_11 D VDD VDD mp15  l=0.13u w=0.6u m=1
M48 VDD D N_11 VDD mp15  l=0.13u w=0.6u m=1
.ends oai33d4
* SPICE INPUT		Tue Jul 31 20:09:01 2018	oaim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d0
.subckt oaim21d0 Y GND VDD C AN BN
M1 N_6 BN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 N_5 GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 AN GND GND mn15  l=0.13u w=0.26u m=1
M5 N_3 BN VDD VDD mp15  l=0.13u w=0.35u m=1
M6 Y N_3 VDD VDD mp15  l=0.13u w=0.35u m=1
M7 VDD C Y VDD mp15  l=0.13u w=0.35u m=1
M8 N_3 AN VDD VDD mp15  l=0.13u w=0.35u m=1
.ends oaim21d0
* SPICE INPUT		Tue Jul 31 20:09:14 2018	oaim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d1
.subckt oaim21d1 Y GND VDD C AN BN
M1 Y N_3 N_5 GND mn15  l=0.13u w=0.46u m=1
M2 GND C N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 AN GND GND mn15  l=0.13u w=0.29u m=1
M4 N_6 BN N_3 GND mn15  l=0.13u w=0.29u m=1
M5 VDD N_3 Y VDD mp15  l=0.13u w=0.61u m=1
M6 VDD C Y VDD mp15  l=0.13u w=0.61u m=1
M7 N_3 AN VDD VDD mp15  l=0.13u w=0.35u m=1
M8 N_3 BN VDD VDD mp15  l=0.13u w=0.35u m=1
.ends oaim21d1
* SPICE INPUT		Tue Jul 31 20:09:27 2018	oaim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d2
.subckt oaim21d2 GND Y VDD C AN BN
M1 Y N_3 N_6 GND mn15  l=0.13u w=0.46u m=1
M2 Y N_3 N_8 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_8 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_7 AN GND GND mn15  l=0.13u w=0.37u m=1
M6 N_7 BN N_3 GND mn15  l=0.13u w=0.37u m=1
M7 VDD N_3 Y VDD mp15  l=0.13u w=0.61u m=1
M8 VDD N_3 Y VDD mp15  l=0.13u w=0.61u m=1
M9 VDD C Y VDD mp15  l=0.13u w=0.61u m=1
M10 Y C VDD VDD mp15  l=0.13u w=0.61u m=1
M11 VDD AN N_3 VDD mp15  l=0.13u w=0.46u m=1
M12 N_3 BN VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oaim21d2
* SPICE INPUT		Tue Jul 31 20:09:40 2018	oaim21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d4
.subckt oaim21d4 GND Y C VDD AN BN
M1 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 C GND GND mn15  l=0.13u w=0.46u m=1
M3 N_13 N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_4 N_12 GND mn15  l=0.13u w=0.46u m=1
M5 N_12 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_11 AN GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_4 N_9 GND mn15  l=0.13u w=0.46u m=1
M8 Y N_4 N_14 GND mn15  l=0.13u w=0.46u m=1
M9 N_11 BN N_4 GND mn15  l=0.13u w=0.46u m=1
M10 N_4 BN N_10 GND mn15  l=0.13u w=0.46u m=1
M11 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M12 N_10 AN GND GND mn15  l=0.13u w=0.46u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.61u m=1
M14 Y C VDD VDD mp15  l=0.13u w=0.61u m=1
M15 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M16 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M17 Y C VDD VDD mp15  l=0.13u w=0.61u m=1
M18 VDD AN N_4 VDD mp15  l=0.13u w=0.57u m=1
M19 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M21 N_4 BN VDD VDD mp15  l=0.13u w=0.57u m=1
M22 N_4 BN VDD VDD mp15  l=0.13u w=0.57u m=1
M23 VDD C Y VDD mp15  l=0.13u w=0.61u m=1
M24 N_4 AN VDD VDD mp15  l=0.13u w=0.57u m=1
.ends oaim21d4
* SPICE INPUT		Tue Jul 31 20:09:53 2018	oaim21dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21dm
.subckt oaim21dm Y GND VDD C AN BN
M1 Y N_3 N_5 GND mn15  l=0.13u w=0.36u m=1
M2 N_6 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 BN N_3 GND mn15  l=0.13u w=0.26u m=1
M4 GND C N_5 GND mn15  l=0.13u w=0.36u m=1
M5 VDD N_3 Y VDD mp15  l=0.13u w=0.45u m=1
M6 N_3 AN VDD VDD mp15  l=0.13u w=0.35u m=1
M7 N_3 BN VDD VDD mp15  l=0.13u w=0.35u m=1
M8 VDD C Y VDD mp15  l=0.13u w=0.45u m=1
.ends oaim21dm
* SPICE INPUT		Tue Jul 31 20:10:06 2018	oaim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d0
.subckt oaim22d0 VDD Y GND D C AN BN
M1 Y N_6 N_10 GND mn15  l=0.13u w=0.26u m=1
M2 N_15 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 N_10 D GND GND mn15  l=0.13u w=0.26u m=1
M4 GND C N_10 GND mn15  l=0.13u w=0.26u m=1
M5 N_15 BN N_6 GND mn15  l=0.13u w=0.26u m=1
M6 N_6 AN VDD VDD mp15  l=0.13u w=0.35u m=1
M7 Y N_6 VDD VDD mp15  l=0.13u w=0.27u m=1
M8 N_7 D Y VDD mp15  l=0.13u w=0.4u m=1
M9 N_7 C VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_6 BN VDD VDD mp15  l=0.13u w=0.35u m=1
.ends oaim22d0
* SPICE INPUT		Tue Jul 31 20:10:19 2018	oaim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d1
.subckt oaim22d1 VDD Y GND D C AN BN
M1 Y N_6 N_10 GND mn15  l=0.13u w=0.46u m=1
M2 N_15 AN GND GND mn15  l=0.13u w=0.29u m=1
M3 N_10 D GND GND mn15  l=0.13u w=0.46u m=1
M4 GND C N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_15 BN N_6 GND mn15  l=0.13u w=0.29u m=1
M6 N_6 AN VDD VDD mp15  l=0.13u w=0.37u m=1
M7 Y N_6 VDD VDD mp15  l=0.13u w=0.48u m=1
M8 N_7 D Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_7 C VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_6 BN VDD VDD mp15  l=0.13u w=0.37u m=1
.ends oaim22d1
* SPICE INPUT		Tue Jul 31 20:10:32 2018	oaim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d2
.subckt oaim22d2 VDD Y GND C D BN AN
M1 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M2 N_14 D GND GND mn15  l=0.13u w=0.46u m=1
M3 N_14 D GND GND mn15  l=0.13u w=0.46u m=1
M4 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_14 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_14 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_5 BN N_19 GND mn15  l=0.13u w=0.46u m=1
M8 GND AN N_19 GND mn15  l=0.13u w=0.46u m=1
M9 VDD C N_9 VDD mp15  l=0.13u w=0.69u m=1
M10 Y D N_9 VDD mp15  l=0.13u w=0.69u m=1
M11 Y D N_10 VDD mp15  l=0.13u w=0.69u m=1
M12 N_10 C VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y N_5 VDD VDD mp15  l=0.13u w=0.47u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.46u m=1
M15 N_5 BN VDD VDD mp15  l=0.13u w=0.6u m=1
M16 N_5 AN VDD VDD mp15  l=0.13u w=0.6u m=1
.ends oaim22d2
* SPICE INPUT		Tue Jul 31 20:10:45 2018	oaim22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d4
.subckt oaim22d4 VDD Y AN BN D GND C
M1 N_27 D GND GND mn15  l=0.13u w=0.46u m=1
M2 N_27 D GND GND mn15  l=0.13u w=0.46u m=1
M3 N_27 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_27 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M5 N_27 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_27 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_27 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 N_27 C GND GND mn15  l=0.13u w=0.46u m=1
M9 N_27 C GND GND mn15  l=0.13u w=0.46u m=1
M10 N_27 D GND GND mn15  l=0.13u w=0.46u m=1
M11 N_27 D GND GND mn15  l=0.13u w=0.46u m=1
M12 N_27 C GND GND mn15  l=0.13u w=0.46u m=1
M13 N_5 BN N_29 GND mn15  l=0.13u w=0.46u m=1
M14 N_5 BN N_30 GND mn15  l=0.13u w=0.46u m=1
M15 N_30 AN GND GND mn15  l=0.13u w=0.46u m=1
M16 GND AN N_29 GND mn15  l=0.13u w=0.46u m=1
M17 N_5 BN VDD VDD mp15  l=0.13u w=0.55u m=1
M18 N_5 BN VDD VDD mp15  l=0.13u w=0.55u m=1
M19 N_5 AN VDD VDD mp15  l=0.13u w=0.55u m=1
M20 N_17 D Y VDD mp15  l=0.13u w=0.69u m=1
M21 Y D N_16 VDD mp15  l=0.13u w=0.69u m=1
M22 N_16 C VDD VDD mp15  l=0.13u w=0.69u m=1
M23 Y N_5 VDD VDD mp15  l=0.13u w=0.46u m=1
M24 Y N_5 VDD VDD mp15  l=0.13u w=0.46u m=1
M25 VDD N_5 Y VDD mp15  l=0.13u w=0.46u m=1
M26 Y N_5 VDD VDD mp15  l=0.13u w=0.46u m=1
M27 N_5 AN VDD VDD mp15  l=0.13u w=0.55u m=1
M28 N_18 C VDD VDD mp15  l=0.13u w=0.69u m=1
M29 N_17 C VDD VDD mp15  l=0.13u w=0.69u m=1
M30 Y D N_15 VDD mp15  l=0.13u w=0.69u m=1
M31 Y D N_18 VDD mp15  l=0.13u w=0.69u m=1
M32 VDD C N_15 VDD mp15  l=0.13u w=0.69u m=1
.ends oaim22d4
* SPICE INPUT		Tue Jul 31 20:10:58 2018	oaim22dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22dm
.subckt oaim22dm VDD Y GND D C AN BN
M1 GND C N_10 GND mn15  l=0.13u w=0.36u m=1
M2 N_15 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 N_15 BN N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_10 D GND GND mn15  l=0.13u w=0.36u m=1
M5 Y N_6 N_10 GND mn15  l=0.13u w=0.36u m=1
M6 Y N_6 VDD VDD mp15  l=0.13u w=0.38u m=1
M7 N_7 C VDD VDD mp15  l=0.13u w=0.55u m=1
M8 N_6 AN VDD VDD mp15  l=0.13u w=0.35u m=1
M9 N_6 BN VDD VDD mp15  l=0.13u w=0.35u m=1
M10 N_7 D Y VDD mp15  l=0.13u w=0.55u m=1
.ends oaim22dm
* SPICE INPUT		Tue Jul 31 20:11:11 2018	or02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d0
.subckt or02d0 VDD Y GND A B
M1 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_5 B N_4 VDD mp15  l=0.13u w=0.4u m=1
M5 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends or02d0
* SPICE INPUT		Tue Jul 31 20:11:24 2018	or02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d1
.subckt or02d1 VDD Y GND A B
M1 N_4 B GND GND mn15  l=0.13u w=0.29u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.29u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 B N_4 VDD mp15  l=0.13u w=0.58u m=1
M5 N_5 A VDD VDD mp15  l=0.13u w=0.58u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or02d1
* SPICE INPUT		Tue Jul 31 20:11:37 2018	or02d1p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d1p5
.subckt or02d1p5 VDD Y A B GND
M1 N_4 B GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M5 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or02d1p5
* SPICE INPUT		Tue Jul 31 20:11:50 2018	or02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d2
.subckt or02d2 Y GND VDD A B
M1 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.35u m=1
M4 N_5 B GND GND mn15  l=0.13u w=0.35u m=1
M5 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M6 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M7 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_11 B N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends or02d2
* SPICE INPUT		Tue Jul 31 20:12:04 2018	or02d2p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d2p5
.subckt or02d2p5 Y VDD GND A B
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_8 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M9 N_5 B N_7 VDD mp15  l=0.13u w=0.69u m=1
M10 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
.ends or02d2p5
* SPICE INPUT		Tue Jul 31 20:12:17 2018	or02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d4
.subckt or02d4 Y GND VDD A B
M1 N_6 A GND GND mn15  l=0.13u w=0.29u m=1
M2 N_6 B GND GND mn15  l=0.13u w=0.29u m=1
M3 N_6 B GND GND mn15  l=0.13u w=0.29u m=1
M4 N_6 A GND GND mn15  l=0.13u w=0.29u m=1
M5 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_16 A VDD VDD mp15  l=0.13u w=0.67u m=1
M10 N_17 B N_6 VDD mp15  l=0.13u w=0.67u m=1
M11 N_6 B N_16 VDD mp15  l=0.13u w=0.67u m=1
M12 N_17 A VDD VDD mp15  l=0.13u w=0.67u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or02d4
* SPICE INPUT		Tue Jul 31 20:12:31 2018	or02d4p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d4p5
.subckt or02d4p5 Y GND VDD A B
M1 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_15 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M12 N_5 B N_15 VDD mp15  l=0.13u w=0.69u m=1
M13 N_15 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_15 VDD mp15  l=0.13u w=0.69u m=1
M15 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or02d4p5
* SPICE INPUT		Tue Jul 31 20:12:44 2018	or02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02dm
.subckt or02dm VDD Y GND A B
M1 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M4 N_5 B N_4 VDD mp15  l=0.13u w=0.4u m=1
M5 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends or02dm
* SPICE INPUT		Tue Jul 31 20:12:57 2018	or02od
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02od
.subckt or02od B A GND VDD Y
M1 N_2 A GND GND mn15  l=0.13u w=0.3u m=1
M2 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M4 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M5 GND B N_2 GND mn15  l=0.13u w=0.3u m=1
M6 VDD A N_18 VDD mp15  l=0.13u w=0.6u m=1
M7 N_2 B N_18 VDD mp15  l=0.13u w=0.6u m=1
.ends or02od
* SPICE INPUT		Tue Jul 31 20:13:10 2018	or03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d0
.subckt or03d0 VDD Y GND A B C
M1 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_4 C GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 B N_7 VDD mp15  l=0.13u w=0.4u m=1
M6 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_7 C N_4 VDD mp15  l=0.13u w=0.4u m=1
.ends or03d0
* SPICE INPUT		Tue Jul 31 20:13:24 2018	or03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d1
.subckt or03d1 VDD Y GND A B C
M1 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.28u m=1
M3 N_4 B GND GND mn15  l=0.13u w=0.28u m=1
M4 N_4 C GND GND mn15  l=0.13u w=0.28u m=1
M5 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M6 N_6 A VDD VDD mp15  l=0.13u w=0.66u m=1
M7 N_6 B N_5 VDD mp15  l=0.13u w=0.66u m=1
M8 N_5 C N_4 VDD mp15  l=0.13u w=0.66u m=1
.ends or03d1
* SPICE INPUT		Tue Jul 31 20:13:37 2018	or03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d2
.subckt or03d2 Y VDD GND A B C
M1 N_4 A GND GND mn15  l=0.13u w=0.34u m=1
M2 N_4 C GND GND mn15  l=0.13u w=0.34u m=1
M3 N_4 B GND GND mn15  l=0.13u w=0.34u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 VDD A N_7 VDD mp15  l=0.13u w=0.69u m=1
M7 N_6 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M8 N_7 B N_6 VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends or03d2
* SPICE INPUT		Tue Jul 31 20:13:50 2018	or03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d4
.subckt or03d4 Y VDD B C A GND
M1 N_5 A GND GND mn15  l=0.13u w=0.32u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND C N_5 GND mn15  l=0.13u w=0.33u m=1
M7 N_5 C GND GND mn15  l=0.13u w=0.33u m=1
M8 GND A N_5 GND mn15  l=0.13u w=0.34u m=1
M9 N_5 B GND GND mn15  l=0.13u w=0.32u m=1
M10 N_5 B GND GND mn15  l=0.13u w=0.34u m=1
M11 VDD A N_9 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M15 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_12 C N_5 VDD mp15  l=0.13u w=0.77u m=1
M17 N_5 C N_10 VDD mp15  l=0.13u w=0.61u m=1
M18 VDD A N_11 VDD mp15  l=0.13u w=0.69u m=1
M19 N_10 B N_9 VDD mp15  l=0.13u w=0.61u m=1
M20 N_12 B N_11 VDD mp15  l=0.13u w=0.77u m=1
.ends or03d4
* SPICE INPUT		Tue Jul 31 20:14:03 2018	or03dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03dm
.subckt or03dm VDD Y GND A B C
M1 N_4 C GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M4 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_7 C N_4 VDD mp15  l=0.13u w=0.4u m=1
M6 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
M8 N_8 B N_7 VDD mp15  l=0.13u w=0.4u m=1
.ends or03dm
* SPICE INPUT		Tue Jul 31 20:14:16 2018	or04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d0
.subckt or04d0 VDD Y GND A B C D
M1 GND C N_4 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_4 D GND GND mn15  l=0.13u w=0.26u m=1
M5 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M6 N_9 C N_8 VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_8 D N_4 VDD mp15  l=0.13u w=0.4u m=1
M10 N_10 B N_9 VDD mp15  l=0.13u w=0.4u m=1
.ends or04d0
* SPICE INPUT		Tue Jul 31 20:14:28 2018	or04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d1
.subckt or04d1 VDD Y GND A B C D
M1 N_4 D GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND C N_4 GND mn15  l=0.13u w=0.26u m=1
M4 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M6 N_8 D N_4 VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_9 C N_8 VDD mp15  l=0.13u w=0.4u m=1
M9 N_10 B N_9 VDD mp15  l=0.13u w=0.4u m=1
M10 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends or04d1
* SPICE INPUT		Tue Jul 31 20:14:41 2018	or04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d2
.subckt or04d2 Y VDD GND A B C D
M1 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_4 D GND GND mn15  l=0.13u w=0.28u m=1
M4 GND C N_4 GND mn15  l=0.13u w=0.28u m=1
M5 N_4 B GND GND mn15  l=0.13u w=0.28u m=1
M6 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_6 D N_4 VDD mp15  l=0.13u w=0.69u m=1
M10 N_7 C N_6 VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 B N_7 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends or04d2
* SPICE INPUT		Tue Jul 31 20:14:54 2018	or04d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d4
.subckt or04d4 Y GND VDD A B C D
M1 N_6 D GND GND mn15  l=0.13u w=0.29u m=1
M2 N_6 D GND GND mn15  l=0.13u w=0.29u m=1
M3 N_6 C GND GND mn15  l=0.13u w=0.29u m=1
M4 N_6 C GND GND mn15  l=0.13u w=0.29u m=1
M5 N_6 A GND GND mn15  l=0.13u w=0.29u m=1
M6 N_6 B GND GND mn15  l=0.13u w=0.29u m=1
M7 N_6 B GND GND mn15  l=0.13u w=0.29u m=1
M8 N_6 A GND GND mn15  l=0.13u w=0.29u m=1
M9 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M13 N_19 D N_6 VDD mp15  l=0.13u w=0.69u m=1
M14 N_6 D N_19 VDD mp15  l=0.13u w=0.69u m=1
M15 N_19 C N_18 VDD mp15  l=0.13u w=0.69u m=1
M16 N_19 C N_18 VDD mp15  l=0.13u w=0.69u m=1
M17 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_25 B N_18 VDD mp15  l=0.13u w=0.69u m=1
M19 N_18 B N_24 VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_25 VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or04d4
* SPICE INPUT		Tue Jul 31 20:15:07 2018	ora211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d0
.subckt ora211d0 VDD Y GND A B C D
M1 N_11 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_11 B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_11 C N_15 GND mn15  l=0.13u w=0.26u m=1
M5 N_15 D N_4 GND mn15  l=0.13u w=0.26u m=1
M6 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_7 B N_4 VDD mp15  l=0.13u w=0.4u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_4 C VDD VDD mp15  l=0.13u w=0.27u m=1
M10 VDD D N_4 VDD mp15  l=0.13u w=0.27u m=1
.ends ora211d0
* SPICE INPUT		Tue Jul 31 20:15:20 2018	ora211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d1
.subckt ora211d1 VDD Y GND A B C D
M1 N_11 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_11 B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_11 C N_15 GND mn15  l=0.13u w=0.26u m=1
M5 N_15 D N_4 GND mn15  l=0.13u w=0.26u m=1
M6 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_7 B N_4 VDD mp15  l=0.13u w=0.4u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_4 C VDD VDD mp15  l=0.13u w=0.27u m=1
M10 VDD D N_4 VDD mp15  l=0.13u w=0.27u m=1
.ends ora211d1
* SPICE INPUT		Tue Jul 31 20:15:33 2018	ora211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d2
.subckt ora211d2 Y GND VDD D C B A
M1 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_6 C N_9 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_6 GND mn15  l=0.13u w=0.46u m=1
M5 N_6 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_5 D N_9 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 C VDD VDD mp15  l=0.13u w=0.48u m=1
M8 N_36 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_36 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 D VDD VDD mp15  l=0.13u w=0.48u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ora211d2
* SPICE INPUT		Tue Jul 31 20:15:46 2018	ora211d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d4
.subckt ora211d4 GND Y VDD C D A B
M1 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_15 D N_8 GND mn15  l=0.13u w=0.46u m=1
M6 N_8 D N_14 GND mn15  l=0.13u w=0.46u m=1
M7 N_15 C N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_2 C N_14 GND mn15  l=0.13u w=0.46u m=1
M9 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M13 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_25 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_26 B N_8 VDD mp15  l=0.13u w=0.69u m=1
M19 N_8 B N_25 VDD mp15  l=0.13u w=0.69u m=1
M20 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_8 D VDD VDD mp15  l=0.13u w=0.46u m=1
M22 N_8 D VDD VDD mp15  l=0.13u w=0.46u m=1
M23 VDD C N_8 VDD mp15  l=0.13u w=0.46u m=1
M24 N_8 C VDD VDD mp15  l=0.13u w=0.46u m=1
.ends ora211d4
* SPICE INPUT		Tue Jul 31 20:15:58 2018	ora21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d0
.subckt ora21d0 VDD Y GND C B A
M1 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_10 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C N_10 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_6 B N_5 VDD mp15  l=0.13u w=0.4u m=1
M8 N_5 C VDD VDD mp15  l=0.13u w=0.27u m=1
.ends ora21d0
* SPICE INPUT		Tue Jul 31 20:16:12 2018	ora21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d1
.subckt ora21d1 VDD Y GND C B A
M1 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_10 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C N_10 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_6 B N_5 VDD mp15  l=0.13u w=0.4u m=1
M7 N_5 C VDD VDD mp15  l=0.13u w=0.27u m=1
M8 Y N_5 VDD VDD mp15  l=0.13u w=0.34u m=1
M9 Y N_5 VDD VDD mp15  l=0.13u w=0.34u m=1
.ends ora21d1
* SPICE INPUT		Tue Jul 31 20:16:24 2018	ora21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d2
.subckt ora21d2 GND Y VDD C B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M4 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_30 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_30 B N_3 VDD mp15  l=0.13u w=0.69u m=1
M8 VDD C N_3 VDD mp15  l=0.13u w=0.48u m=1
M9 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ora21d2
* SPICE INPUT		Tue Jul 31 20:16:38 2018	ora21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d4
.subckt ora21d4 GND Y VDD C A B
M1 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M7 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M10 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M11 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_21 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M13 N_2 B N_20 VDD mp15  l=0.13u w=0.69u m=1
M14 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD C N_2 VDD mp15  l=0.13u w=0.48u m=1
M16 VDD C N_2 VDD mp15  l=0.13u w=0.48u m=1
M17 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora21d4
* SPICE INPUT		Tue Jul 31 20:16:51 2018	ora221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora221d0
.subckt ora221d0 VDD Y GND E D C A B
M1 GND A N_16 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_16 GND mn15  l=0.13u w=0.26u m=1
M3 N_14 C N_16 GND mn15  l=0.13u w=0.26u m=1
M4 N_14 D N_16 GND mn15  l=0.13u w=0.26u m=1
M5 N_3 E N_14 GND mn15  l=0.13u w=0.26u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_8 B N_3 VDD mp15  l=0.13u w=0.4u m=1
M9 N_9 C VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_9 D N_3 VDD mp15  l=0.13u w=0.4u m=1
M11 N_3 E VDD VDD mp15  l=0.13u w=0.27u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ora221d0
* SPICE INPUT		Tue Jul 31 20:17:05 2018	ora221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora221d1
.subckt ora221d1 VDD Y GND E D C A B
M1 GND B N_16 GND mn15  l=0.13u w=0.26u m=1
M2 GND A N_16 GND mn15  l=0.13u w=0.26u m=1
M3 N_14 C N_16 GND mn15  l=0.13u w=0.26u m=1
M4 N_14 D N_16 GND mn15  l=0.13u w=0.26u m=1
M5 N_3 E N_14 GND mn15  l=0.13u w=0.26u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_8 B N_3 VDD mp15  l=0.13u w=0.4u m=1
M8 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_9 C VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_9 D N_3 VDD mp15  l=0.13u w=0.4u m=1
M11 N_3 E VDD VDD mp15  l=0.13u w=0.27u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora221d1
* SPICE INPUT		Tue Jul 31 20:17:18 2018	ora221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora221d2
.subckt ora221d2 Y GND VDD E D C A B
M1 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_6 C N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_10 E N_6 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 D N_6 GND mn15  l=0.13u w=0.46u m=1
M8 VDD E N_10 VDD mp15  l=0.13u w=0.48u m=1
M9 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_15 D N_10 VDD mp15  l=0.13u w=0.35u m=1
M12 N_15 D N_10 VDD mp15  l=0.13u w=0.34u m=1
M13 VDD A N_44 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD C N_15 VDD mp15  l=0.13u w=0.69u m=1
M15 N_44 B N_10 VDD mp15  l=0.13u w=0.69u m=1
.ends ora221d2
* SPICE INPUT		Tue Jul 31 20:17:32 2018	ora221d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora221d4
.subckt ora221d4 GND Y VDD E D C A B
M1 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M2 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_2 C N_3 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M7 N_2 D N_3 GND mn15  l=0.13u w=0.565u m=1
M8 N_3 D N_2 GND mn15  l=0.13u w=0.355u m=1
M9 GND N_16 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_16 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_16 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_16 Y GND mn15  l=0.13u w=0.46u m=1
M13 N_3 E N_16 GND mn15  l=0.13u w=0.565u m=1
M14 N_3 E N_16 GND mn15  l=0.13u w=0.355u m=1
M15 N_16 B N_28 VDD mp15  l=0.13u w=0.69u m=1
M16 N_16 B N_24 VDD mp15  l=0.13u w=0.69u m=1
M17 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_19 C VDD VDD mp15  l=0.13u w=0.46u m=1
M20 VDD C N_19 VDD mp15  l=0.13u w=0.46u m=1
M21 N_19 C VDD VDD mp15  l=0.13u w=0.46u m=1
M22 N_16 D N_19 VDD mp15  l=0.13u w=0.56u m=1
M23 N_16 D N_19 VDD mp15  l=0.13u w=0.56u m=1
M24 N_16 D N_19 VDD mp15  l=0.13u w=0.26u m=1
M25 N_16 E VDD VDD mp15  l=0.13u w=0.6u m=1
M26 N_16 E VDD VDD mp15  l=0.13u w=0.36u m=1
M27 VDD N_16 Y VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_16 Y VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_16 Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora221d4
* SPICE INPUT		Tue Jul 31 20:17:45 2018	ora222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora222d0
.subckt ora222d0 VDD Y GND F E C D B A
M1 GND A N_19 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_19 GND mn15  l=0.13u w=0.26u m=1
M3 N_17 D N_19 GND mn15  l=0.13u w=0.26u m=1
M4 N_19 C N_17 GND mn15  l=0.13u w=0.26u m=1
M5 N_2 E N_17 GND mn15  l=0.13u w=0.26u m=1
M6 N_2 F N_17 GND mn15  l=0.13u w=0.26u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_2 B N_12 VDD mp15  l=0.13u w=0.4u m=1
M10 N_13 D N_2 VDD mp15  l=0.13u w=0.4u m=1
M11 N_13 C VDD VDD mp15  l=0.13u w=0.4u m=1
M12 VDD E N_11 VDD mp15  l=0.13u w=0.4u m=1
M13 N_2 F N_11 VDD mp15  l=0.13u w=0.4u m=1
M14 Y N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ora222d0
* SPICE INPUT		Tue Jul 31 20:17:58 2018	ora222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora222d1
.subckt ora222d1 VDD Y GND F E C D B A
M1 GND A N_19 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_19 GND mn15  l=0.13u w=0.26u m=1
M3 N_17 D N_19 GND mn15  l=0.13u w=0.26u m=1
M4 N_19 C N_17 GND mn15  l=0.13u w=0.26u m=1
M5 N_2 E N_17 GND mn15  l=0.13u w=0.26u m=1
M6 N_2 F N_17 GND mn15  l=0.13u w=0.26u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_2 B N_12 VDD mp15  l=0.13u w=0.4u m=1
M10 N_13 D N_2 VDD mp15  l=0.13u w=0.4u m=1
M11 N_13 C VDD VDD mp15  l=0.13u w=0.4u m=1
M12 VDD E N_11 VDD mp15  l=0.13u w=0.4u m=1
M13 N_2 F N_11 VDD mp15  l=0.13u w=0.4u m=1
M14 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora222d1
* SPICE INPUT		Tue Jul 31 20:18:11 2018	ora222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora222d2
.subckt ora222d2 GND Y VDD E F C D B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 D N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 E N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 F N_7 GND mn15  l=0.13u w=0.46u m=1
M7 GND N_7 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_7 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_7 D N_24 VDD mp15  l=0.13u w=0.34u m=1
M10 N_25 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_25 B N_7 VDD mp15  l=0.13u w=0.69u m=1
M12 N_26 D N_7 VDD mp15  l=0.13u w=0.35u m=1
M13 N_26 C VDD VDD mp15  l=0.13u w=0.35u m=1
M14 VDD C N_24 VDD mp15  l=0.13u w=0.34u m=1
M15 VDD N_7 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_7 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD E N_27 VDD mp15  l=0.13u w=0.69u m=1
M18 N_27 F N_7 VDD mp15  l=0.13u w=0.69u m=1
.ends ora222d2
* SPICE INPUT		Tue Jul 31 20:18:24 2018	ora222d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora222d4
.subckt ora222d4 GND Y F VDD E C D B A
M1 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 D N_2 GND mn15  l=0.13u w=0.45u m=1
M6 N_2 C N_3 GND mn15  l=0.13u w=0.56u m=1
M7 N_2 C N_3 GND mn15  l=0.13u w=0.36u m=1
M8 N_3 D N_2 GND mn15  l=0.13u w=0.47u m=1
M9 N_3 F N_11 GND mn15  l=0.13u w=0.565u m=1
M10 N_3 F N_11 GND mn15  l=0.13u w=0.355u m=1
M11 N_3 E N_11 GND mn15  l=0.13u w=0.565u m=1
M12 N_3 E N_11 GND mn15  l=0.13u w=0.355u m=1
M13 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_11 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M16 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M17 N_37 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M18 N_38 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_37 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_11 B N_38 VDD mp15  l=0.13u w=0.69u m=1
M21 N_11 F N_36 VDD mp15  l=0.13u w=0.55u m=1
M22 N_42 E VDD VDD mp15  l=0.13u w=0.42u m=1
M23 VDD E N_36 VDD mp15  l=0.13u w=0.55u m=1
M24 VDD E N_43 VDD mp15  l=0.13u w=0.41u m=1
M25 N_11 D N_39 VDD mp15  l=0.13u w=0.69u m=1
M26 N_40 C VDD VDD mp15  l=0.13u w=0.27u m=1
M27 VDD C N_39 VDD mp15  l=0.13u w=0.605u m=1
M28 N_40 D N_11 VDD mp15  l=0.13u w=0.27u m=1
M29 N_41 D N_11 VDD mp15  l=0.13u w=0.42u m=1
M30 N_41 C VDD VDD mp15  l=0.13u w=0.505u m=1
M31 N_43 F N_11 VDD mp15  l=0.13u w=0.41u m=1
M32 N_11 F N_42 VDD mp15  l=0.13u w=0.42u m=1
M33 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
M34 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
M36 Y N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora222d4
* SPICE INPUT		Tue Jul 31 20:18:37 2018	ora22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora22d0
.subckt ora22d0 VDD Y GND C D B A
M1 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_13 D N_4 GND mn15  l=0.13u w=0.26u m=1
M3 N_13 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_13 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_13 C N_4 GND mn15  l=0.13u w=0.26u m=1
M6 N_4 D N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_4 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M9 VDD C N_7 VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ora22d0
* SPICE INPUT		Tue Jul 31 20:18:51 2018	ora22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora22d1
.subckt ora22d1 VDD Y GND C D B A
M1 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 D N_4 GND mn15  l=0.13u w=0.26u m=1
M3 N_13 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_13 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_13 C N_4 GND mn15  l=0.13u w=0.26u m=1
M6 N_4 D N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_4 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M9 VDD C N_7 VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora22d1
* SPICE INPUT		Tue Jul 31 20:19:03 2018	ora22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora22d2
.subckt ora22d2 Y GND VDD C D B A
M1 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_6 C N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_6 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 D N_5 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_6 GND mn15  l=0.13u w=0.46u m=1
M7 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_12 C VDD VDD mp15  l=0.13u w=0.345u m=1
M10 N_12 C VDD VDD mp15  l=0.13u w=0.345u m=1
M11 N_5 B N_17 VDD mp15  l=0.13u w=0.69u m=1
M12 N_5 D N_12 VDD mp15  l=0.13u w=0.69u m=1
M13 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora22d2
* SPICE INPUT		Tue Jul 31 20:19:16 2018	ora22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora22d4
.subckt ora22d4 GND Y VDD C D A B
M1 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M9 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M13 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_27 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M15 N_2 B N_26 VDD mp15  l=0.13u w=0.69u m=1
M16 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_2 D N_25 VDD mp15  l=0.13u w=0.6u m=1
M18 N_2 D N_28 VDD mp15  l=0.13u w=0.6u m=1
M19 N_25 C VDD VDD mp15  l=0.13u w=0.6u m=1
M20 N_28 C VDD VDD mp15  l=0.13u w=0.6u m=1
M21 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora22d4
* SPICE INPUT		Tue Jul 31 20:19:29 2018	ora31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d0
.subckt ora31d0 VDD Y A B C GND D
M1 N_11 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_11 B GND GND mn15  l=0.13u w=0.26u m=1
M3 N_11 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_11 D N_5 GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_9 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_9 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M8 N_8 C N_5 VDD mp15  l=0.13u w=0.4u m=1
M9 N_5 D VDD VDD mp15  l=0.13u w=0.27u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ora31d0
* SPICE INPUT		Tue Jul 31 20:19:42 2018	ora31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d1
.subckt ora31d1 VDD Y GND A B C D
M1 N_12 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_12 D N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_12 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_12 B GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_9 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_5 D VDD VDD mp15  l=0.13u w=0.27u m=1
M8 N_8 C N_5 VDD mp15  l=0.13u w=0.4u m=1
M9 N_9 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora31d1
* SPICE INPUT		Tue Jul 31 20:19:55 2018	ora31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d2
.subckt ora31d2 Y GND VDD A B C D
M1 N_6 D N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_6 C GND GND mn15  l=0.13u w=0.46u m=1
M3 N_6 B GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_6 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_4 D VDD VDD mp15  l=0.13u w=0.48u m=1
M8 N_31 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M9 N_32 B N_31 VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_32 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ora31d2
* SPICE INPUT		Tue Jul 31 20:20:08 2018	ora31d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d4
.subckt ora31d4 GND Y D VDD C B A
M1 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M7 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M8 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M13 VDD D N_2 VDD mp15  l=0.13u w=0.48u m=1
M14 VDD D N_2 VDD mp15  l=0.13u w=0.48u m=1
M15 N_60 C N_2 VDD mp15  l=0.13u w=0.69u m=1
M16 N_61 B N_60 VDD mp15  l=0.13u w=0.69u m=1
M17 N_61 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_62 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_63 C N_2 VDD mp15  l=0.13u w=0.69u m=1
M20 N_63 B N_62 VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora31d4



* SPICE INPUT		Tue Jul 31 20:36:45 2018	xn02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d0
.subckt xn02d0 GND Y VDD B A
M1 N_7 B GND GND mn15  l=0.13u w=0.3u m=1
M2 N_8 N_7 GND GND mn15  l=0.13u w=0.23u m=1
M3 N_7 A N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_8 N_5 N_6 GND mn15  l=0.13u w=0.23u m=1
M7 N_7 B VDD VDD mp15  l=0.13u w=0.45u m=1
M8 N_14 N_7 VDD VDD mp15  l=0.13u w=0.33u m=1
M9 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_6 A N_14 VDD mp15  l=0.13u w=0.33u m=1
M11 Y N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M12 N_7 N_5 N_6 VDD mp15  l=0.13u w=0.26u m=1
.ends xn02d0
* SPICE INPUT		Tue Jul 31 20:36:59 2018	xn02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d1
.subckt xn02d1 GND Y VDD B A
M1 N_8 N_7 GND GND mn15  l=0.13u w=0.3u m=1
M2 N_8 N_4 N_6 GND mn15  l=0.13u w=0.3u m=1
M3 N_7 A N_6 GND mn15  l=0.13u w=0.3u m=1
M4 GND A N_4 GND mn15  l=0.13u w=0.26u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.33u m=1
M6 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_32 N_7 VDD VDD mp15  l=0.13u w=0.45u m=1
M8 N_7 N_4 N_6 VDD mp15  l=0.13u w=0.3u m=1
M9 N_6 A N_32 VDD mp15  l=0.13u w=0.45u m=1
M10 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M11 N_7 B VDD VDD mp15  l=0.13u w=0.5u m=1
M12 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends xn02d1
* SPICE INPUT		Tue Jul 31 20:37:12 2018	xn02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d2
.subckt xn02d2 GND Y VDD A B
M1 GND B N_2 GND mn15  l=0.13u w=0.41u m=1
M2 N_10 N_2 GND GND mn15  l=0.13u w=0.41u m=1
M3 N_10 N_8 N_3 GND mn15  l=0.13u w=0.41u m=1
M4 N_3 A N_2 GND mn15  l=0.13u w=0.39u m=1
M5 GND A N_8 GND mn15  l=0.13u w=0.26u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M8 VDD B N_2 VDD mp15  l=0.13u w=0.63u m=1
M9 N_16 N_2 VDD VDD mp15  l=0.13u w=0.63u m=1
M10 N_2 N_8 N_3 VDD mp15  l=0.13u w=0.31u m=1
M11 N_16 A N_3 VDD mp15  l=0.13u w=0.63u m=1
M12 VDD A N_8 VDD mp15  l=0.13u w=0.4u m=1
M13 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
.ends xn02d2
* SPICE INPUT		Tue Jul 31 20:37:25 2018	xn02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d4
.subckt xn02d4 Y GND VDD B A
M1 N_4 A N_2 GND mn15  l=0.13u w=0.37u m=1
M2 N_4 A N_2 GND mn15  l=0.13u w=0.37u m=1
M3 GND A N_8 GND mn15  l=0.13u w=0.19u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.19u m=1
M5 N_10 N_8 N_2 GND mn15  l=0.13u w=0.53u m=1
M6 N_2 N_8 N_10 GND mn15  l=0.13u w=0.27u m=1
M7 N_10 N_4 GND GND mn15  l=0.13u w=0.35u m=1
M8 GND N_4 N_10 GND mn15  l=0.13u w=0.45u m=1
M9 GND B N_4 GND mn15  l=0.13u w=0.42u m=1
M10 N_4 B GND GND mn15  l=0.13u w=0.42u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M14 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M15 N_4 N_8 N_2 VDD mp15  l=0.13u w=0.46u m=1
M16 N_4 N_8 N_2 VDD mp15  l=0.13u w=0.46u m=1
M17 N_8 A VDD VDD mp15  l=0.13u w=0.6u m=1
M18 N_2 A N_20 VDD mp15  l=0.13u w=0.62u m=1
M19 N_2 A N_20 VDD mp15  l=0.13u w=0.62u m=1
M20 N_20 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_4 N_20 VDD mp15  l=0.13u w=0.55u m=1
M22 N_4 B VDD VDD mp15  l=0.13u w=0.63u m=1
M23 N_4 B VDD VDD mp15  l=0.13u w=0.63u m=1
M24 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M26 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M27 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends xn02d4
* SPICE INPUT		Tue Jul 31 20:37:39 2018	xn02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02dm
.subckt xn02dm GND Y VDD B A
M1 N_8 N_7 GND GND mn15  l=0.13u w=0.23u m=1
M2 N_7 A N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 B GND GND mn15  l=0.13u w=0.3u m=1
M5 Y N_6 GND GND mn15  l=0.13u w=0.36u m=1
M6 N_8 N_5 N_6 GND mn15  l=0.13u w=0.23u m=1
M7 N_14 N_7 VDD VDD mp15  l=0.13u w=0.33u m=1
M8 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_6 A N_14 VDD mp15  l=0.13u w=0.33u m=1
M10 N_7 B VDD VDD mp15  l=0.13u w=0.45u m=1
M11 Y N_6 VDD VDD mp15  l=0.13u w=0.55u m=1
M12 N_7 N_5 N_6 VDD mp15  l=0.13u w=0.26u m=1
.ends xn02dm
* SPICE INPUT		Tue Jul 31 20:37:52 2018	xn03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d0
.subckt xn03d0 GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_13 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_13 A N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_11 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_12 C GND GND mn15  l=0.13u w=0.28u m=1
M9 N_14 N_12 GND GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 N_11 GND mn15  l=0.13u w=0.28u m=1
M11 N_12 N_3 N_11 GND mn15  l=0.13u w=0.28u m=1
M12 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M13 N_23 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_7 A N_6 VDD mp15  l=0.13u w=0.28u m=1
M15 N_23 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_3 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 Y N_11 VDD VDD mp15  l=0.13u w=0.4u m=1
M19 N_12 C VDD VDD mp15  l=0.13u w=0.4u m=1
M20 N_12 N_6 N_11 VDD mp15  l=0.13u w=0.28u m=1
M21 N_24 N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 N_24 N_3 N_11 VDD mp15  l=0.13u w=0.4u m=1
.ends xn03d0
* SPICE INPUT		Tue Jul 31 20:38:05 2018	xn03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d1
.subckt xn03d1 GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_13 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_13 A N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_11 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_12 C GND GND mn15  l=0.13u w=0.28u m=1
M9 N_14 N_12 GND GND mn15  l=0.13u w=0.3u m=1
M10 N_14 N_6 N_11 GND mn15  l=0.13u w=0.3u m=1
M11 N_12 N_3 N_11 GND mn15  l=0.13u w=0.28u m=1
M12 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M13 N_23 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_7 A N_6 VDD mp15  l=0.13u w=0.28u m=1
M15 N_23 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_3 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 Y N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_12 C VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_12 N_6 N_11 VDD mp15  l=0.13u w=0.28u m=1
M21 N_24 N_12 VDD VDD mp15  l=0.13u w=0.45u m=1
M22 N_24 N_3 N_11 VDD mp15  l=0.13u w=0.45u m=1
.ends xn03d1
* SPICE INPUT		Tue Jul 31 20:38:18 2018	xn03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d2
.subckt xn03d2 GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_14 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_14 A N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M7 N_15 N_12 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_15 N_6 N_11 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 N_3 N_11 GND mn15  l=0.13u w=0.45u m=1
M10 GND C N_12 GND mn15  l=0.13u w=0.42u m=1
M11 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M13 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M14 N_60 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M15 N_7 A N_6 VDD mp15  l=0.13u w=0.36u m=1
M16 N_60 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M17 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_3 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M19 N_61 N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_61 N_3 N_11 VDD mp15  l=0.13u w=0.69u m=1
M21 N_12 N_6 N_11 VDD mp15  l=0.13u w=0.57u m=1
M22 N_12 C VDD VDD mp15  l=0.13u w=0.62u m=1
M23 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
.ends xn03d2
* SPICE INPUT		Tue Jul 31 20:38:31 2018	xn03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d4
.subckt xn03d4 GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_18 N_7 GND GND mn15  l=0.13u w=0.38u m=1
M3 N_18 A N_6 GND mn15  l=0.13u w=0.38u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.38u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.33u m=1
M7 N_10 N_6 N_19 GND mn15  l=0.13u w=0.32u m=1
M8 N_10 N_6 N_20 GND mn15  l=0.13u w=0.32u m=1
M9 GND N_14 N_20 GND mn15  l=0.13u w=0.44u m=1
M10 N_19 N_14 GND GND mn15  l=0.13u w=0.2u m=1
M11 N_14 N_3 N_10 GND mn15  l=0.13u w=0.5u m=1
M12 GND C N_14 GND mn15  l=0.13u w=0.46u m=1
M13 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M14 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M15 Y N_10 GND GND mn15  l=0.13u w=0.46u m=1
M16 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M17 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M18 N_79 N_7 VDD VDD mp15  l=0.13u w=0.57u m=1
M19 N_79 N_4 N_6 VDD mp15  l=0.13u w=0.57u m=1
M20 N_7 A N_6 VDD mp15  l=0.13u w=0.38u m=1
M21 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M22 N_3 N_6 VDD VDD mp15  l=0.13u w=0.52u m=1
M23 N_81 N_3 N_10 VDD mp15  l=0.13u w=0.425u m=1
M24 N_10 N_3 N_80 VDD mp15  l=0.13u w=0.425u m=1
M25 N_80 N_14 VDD VDD mp15  l=0.13u w=0.53u m=1
M26 N_81 N_14 VDD VDD mp15  l=0.13u w=0.32u m=1
M27 N_14 N_6 N_10 VDD mp15  l=0.13u w=0.5u m=1
M28 N_14 C VDD VDD mp15  l=0.13u w=0.66u m=1
M29 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends xn03d4
* SPICE INPUT		Tue Jul 31 20:38:44 2018	xn03dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03dm
.subckt xn03dm GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_13 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_13 A N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_11 GND GND mn15  l=0.13u w=0.36u m=1
M8 N_12 C GND GND mn15  l=0.13u w=0.28u m=1
M9 N_14 N_12 GND GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 N_11 GND mn15  l=0.13u w=0.28u m=1
M11 N_12 N_3 N_11 GND mn15  l=0.13u w=0.28u m=1
M12 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M13 N_23 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_7 A N_6 VDD mp15  l=0.13u w=0.28u m=1
M15 N_23 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_3 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 Y N_11 VDD VDD mp15  l=0.13u w=0.55u m=1
M19 N_12 C VDD VDD mp15  l=0.13u w=0.4u m=1
M20 N_12 N_6 N_11 VDD mp15  l=0.13u w=0.28u m=1
M21 N_24 N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 N_24 N_3 N_11 VDD mp15  l=0.13u w=0.4u m=1
.ends xn03dm
* SPICE INPUT		Tue Jul 31 20:38:58 2018	xr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d0
.subckt xr02d0 GND Y A VDD B
M1 GND B N_3 GND mn15  l=0.13u w=0.28u m=1
M2 N_9 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_3 N_8 N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_9 A N_2 GND mn15  l=0.13u w=0.26u m=1
M5 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M6 Y N_2 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_3 B VDD VDD mp15  l=0.13u w=0.42u m=1
M8 N_15 N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_15 N_8 N_2 VDD mp15  l=0.13u w=0.4u m=1
M10 N_2 A N_3 VDD mp15  l=0.13u w=0.26u m=1
M11 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M12 Y N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr02d0
* SPICE INPUT		Tue Jul 31 20:39:12 2018	xr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d1
.subckt xr02d1 GND Y A VDD B
M1 GND B N_3 GND mn15  l=0.13u w=0.32u m=1
M2 N_9 N_3 GND GND mn15  l=0.13u w=0.32u m=1
M3 N_3 N_8 N_2 GND mn15  l=0.13u w=0.28u m=1
M4 N_9 A N_2 GND mn15  l=0.13u w=0.32u m=1
M5 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M7 VDD B N_3 VDD mp15  l=0.13u w=0.52u m=1
M8 N_34 N_3 VDD VDD mp15  l=0.13u w=0.52u m=1
M9 N_34 N_8 N_2 VDD mp15  l=0.13u w=0.52u m=1
M10 N_2 A N_3 VDD mp15  l=0.13u w=0.42u m=1
M11 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr02d1
* SPICE INPUT		Tue Jul 31 20:39:24 2018	xr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d2
.subckt xr02d2 Y GND VDD A B
M1 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.26u m=1
M4 GND B N_7 GND mn15  l=0.13u w=0.41u m=1
M5 N_10 N_7 GND GND mn15  l=0.13u w=0.39u m=1
M6 N_7 N_4 N_6 GND mn15  l=0.13u w=0.32u m=1
M7 N_10 A N_6 GND mn15  l=0.13u w=0.39u m=1
M8 N_7 B VDD VDD mp15  l=0.13u w=0.63u m=1
M9 N_38 N_7 VDD VDD mp15  l=0.13u w=0.54u m=1
M10 N_38 N_4 N_6 VDD mp15  l=0.13u w=0.54u m=1
M11 N_6 A N_7 VDD mp15  l=0.13u w=0.46u m=1
M12 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr02d2
* SPICE INPUT		Tue Jul 31 20:39:37 2018	xr02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d4
.subckt xr02d4 GND Y VDD A B
M1 N_5 B GND GND mn15  l=0.13u w=0.42u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.42u m=1
M3 N_17 N_5 GND GND mn15  l=0.13u w=0.51u m=1
M4 N_18 N_5 GND GND mn15  l=0.13u w=0.27u m=1
M5 N_17 A N_6 GND mn15  l=0.13u w=0.51u m=1
M6 N_18 A N_6 GND mn15  l=0.13u w=0.27u m=1
M7 N_6 N_13 N_5 GND mn15  l=0.13u w=0.26u m=1
M8 N_5 N_13 N_6 GND mn15  l=0.13u w=0.26u m=1
M9 N_5 N_13 N_6 GND mn15  l=0.13u w=0.24u m=1
M10 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M11 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M14 GND A N_13 GND mn15  l=0.13u w=0.41u m=1
M15 VDD B N_5 VDD mp15  l=0.13u w=0.66u m=1
M16 VDD B N_5 VDD mp15  l=0.13u w=0.59u m=1
M17 VDD N_5 N_23 VDD mp15  l=0.13u w=0.59u m=1
M18 VDD N_5 N_23 VDD mp15  l=0.13u w=0.59u m=1
M19 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_13 A VDD VDD mp15  l=0.13u w=0.61u m=1
M24 N_23 N_13 N_6 VDD mp15  l=0.13u w=0.59u m=1
M25 N_23 N_13 N_6 VDD mp15  l=0.13u w=0.59u m=1
M26 N_6 A N_5 VDD mp15  l=0.13u w=0.52u m=1
M27 N_6 A N_5 VDD mp15  l=0.13u w=0.42u m=1
.ends xr02d4
* SPICE INPUT		Tue Jul 31 20:39:49 2018	xr02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02dm
.subckt xr02dm VDD Y GND A B
M1 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.36u m=1
M3 GND B N_2 GND mn15  l=0.13u w=0.28u m=1
M4 N_14 N_2 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_3 N_8 N_2 GND mn15  l=0.13u w=0.3u m=1
M6 N_14 A N_3 GND mn15  l=0.13u w=0.26u m=1
M7 N_2 B VDD VDD mp15  l=0.13u w=0.42u m=1
M8 N_9 N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_9 N_8 N_3 VDD mp15  l=0.13u w=0.4u m=1
M10 N_3 A N_2 VDD mp15  l=0.13u w=0.3u m=1
M11 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends xr02dm
* SPICE INPUT		Tue Jul 31 20:40:02 2018	xr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d0
.subckt xr03d0 GND Y VDD B A C
M1 N_3 A GND GND mn15  l=0.13u w=0.28u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.28u m=1
M3 N_15 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_15 N_3 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_5 A N_6 GND mn15  l=0.13u w=0.28u m=1
M6 GND C N_9 GND mn15  l=0.13u w=0.28u m=1
M7 N_16 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_9 N_14 N_8 GND mn15  l=0.13u w=0.28u m=1
M9 N_16 N_6 N_8 GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M11 Y N_8 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_58 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.28u m=1
M15 N_58 A N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 VDD C N_9 VDD mp15  l=0.13u w=0.4u m=1
M17 N_59 N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_59 N_14 N_8 VDD mp15  l=0.13u w=0.4u m=1
M19 N_9 N_6 N_8 VDD mp15  l=0.13u w=0.28u m=1
M20 N_3 A VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_14 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 Y N_8 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr03d0
* SPICE INPUT		Tue Jul 31 20:40:15 2018	xr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d1
.subckt xr03d1 GND Y VDD B A C
M1 N_3 A GND GND mn15  l=0.13u w=0.28u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.28u m=1
M3 N_15 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_15 N_3 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_5 A N_6 GND mn15  l=0.13u w=0.28u m=1
M6 GND C N_9 GND mn15  l=0.13u w=0.28u m=1
M7 N_16 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_9 N_14 N_8 GND mn15  l=0.13u w=0.28u m=1
M9 N_16 N_6 N_8 GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M11 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_60 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.28u m=1
M15 N_60 A N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 VDD C N_9 VDD mp15  l=0.13u w=0.4u m=1
M17 N_61 N_9 VDD VDD mp15  l=0.13u w=0.42u m=1
M18 N_61 N_14 N_8 VDD mp15  l=0.13u w=0.42u m=1
M19 N_9 N_6 N_8 VDD mp15  l=0.13u w=0.28u m=1
M20 N_3 A VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_14 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends xr03d1
* SPICE INPUT		Tue Jul 31 20:40:28 2018	xr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d2
.subckt xr03d2 VDD Y GND B A C
M1 N_3 A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_23 N_11 N_4 GND mn15  l=0.13u w=0.28u m=1
M3 N_23 N_3 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_3 B GND GND mn15  l=0.13u w=0.28u m=1
M5 GND N_4 N_13 GND mn15  l=0.13u w=0.28u m=1
M6 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_11 A GND GND mn15  l=0.13u w=0.28u m=1
M9 GND C N_7 GND mn15  l=0.13u w=0.42u m=1
M10 N_24 N_7 GND GND mn15  l=0.13u w=0.45u m=1
M11 N_7 N_13 N_6 GND mn15  l=0.13u w=0.21u m=1
M12 N_6 N_13 N_7 GND mn15  l=0.13u w=0.2u m=1
M13 N_24 N_4 N_6 GND mn15  l=0.13u w=0.45u m=1
M14 N_15 A N_4 VDD mp15  l=0.13u w=0.4u m=1
M15 N_3 N_11 N_4 VDD mp15  l=0.13u w=0.33u m=1
M16 N_15 N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M18 VDD C N_7 VDD mp15  l=0.13u w=0.62u m=1
M19 N_16 N_7 VDD VDD mp15  l=0.13u w=0.67u m=1
M20 N_16 N_13 N_6 VDD mp15  l=0.13u w=0.67u m=1
M21 N_7 N_4 N_6 VDD mp15  l=0.13u w=0.56u m=1
M22 N_13 N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M23 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_11 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr03d2
* SPICE INPUT		Tue Jul 31 20:40:41 2018	xr03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d4
.subckt xr03d4 VDD Y C A B GND
M1 N_3 B GND GND mn15  l=0.13u w=0.28u m=1
M2 N_80 N_3 GND GND mn15  l=0.13u w=0.38u m=1
M3 N_80 N_7 N_5 GND mn15  l=0.13u w=0.38u m=1
M4 N_3 A N_5 GND mn15  l=0.13u w=0.36u m=1
M5 N_7 A GND GND mn15  l=0.13u w=0.28u m=1
M6 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M10 GND N_5 N_9 GND mn15  l=0.13u w=0.34u m=1
M11 N_14 N_9 N_13 GND mn15  l=0.13u w=0.23u m=1
M12 N_13 N_9 N_14 GND mn15  l=0.13u w=0.23u m=1
M13 N_82 N_5 N_13 GND mn15  l=0.13u w=0.43u m=1
M14 N_13 N_5 N_81 GND mn15  l=0.13u w=0.23u m=1
M15 N_81 N_14 GND GND mn15  l=0.13u w=0.23u m=1
M16 N_82 N_14 GND GND mn15  l=0.13u w=0.43u m=1
M17 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M18 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M19 N_19 N_3 VDD VDD mp15  l=0.13u w=0.58u m=1
M20 N_5 N_7 N_3 VDD mp15  l=0.13u w=0.33u m=1
M21 N_19 A N_5 VDD mp15  l=0.13u w=0.58u m=1
M22 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M23 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_9 N_5 VDD VDD mp15  l=0.13u w=0.52u m=1
M28 N_14 N_5 N_13 VDD mp15  l=0.13u w=0.46u m=1
M29 VDD N_14 N_20 VDD mp15  l=0.13u w=0.31u m=1
M30 N_21 N_14 VDD VDD mp15  l=0.13u w=0.62u m=1
M31 N_14 C VDD VDD mp15  l=0.13u w=0.66u m=1
M32 N_21 N_9 N_13 VDD mp15  l=0.13u w=0.62u m=1
M33 N_13 N_9 N_20 VDD mp15  l=0.13u w=0.31u m=1
.ends xr03d4
* SPICE INPUT		Tue Jul 31 20:40:54 2018	xr03dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03dm
.subckt xr03dm GND Y VDD B A C
M1 N_3 A GND GND mn15  l=0.13u w=0.28u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.28u m=1
M3 N_15 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_15 N_3 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_5 A N_6 GND mn15  l=0.13u w=0.3u m=1
M6 GND C N_9 GND mn15  l=0.13u w=0.28u m=1
M7 N_16 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_9 N_14 N_8 GND mn15  l=0.13u w=0.28u m=1
M9 N_16 N_6 N_8 GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M11 Y N_8 GND GND mn15  l=0.13u w=0.36u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_58 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.3u m=1
M15 N_58 A N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 VDD C N_9 VDD mp15  l=0.13u w=0.4u m=1
M17 N_59 N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_59 N_14 N_8 VDD mp15  l=0.13u w=0.4u m=1
M19 N_9 N_6 N_8 VDD mp15  l=0.13u w=0.28u m=1
M20 N_3 A VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_14 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 Y N_8 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends xr03dm
