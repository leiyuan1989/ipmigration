* SPICE INPUT		Wed Jul 10 13:34:20 2019	dfbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb1
.subckt dfbfb1 VDD QN Q GND RN SN CKN D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_26 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_6 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CKN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_6 N_28 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M18 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_6 N_5 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_4 N_5 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_4 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_6 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M38 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfbfb1
* SPICE INPUT		Wed Jul 10 13:34:27 2019	dfbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb2
.subckt dfbfb2 VDD QN Q GND RN SN CKN D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_26 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_6 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CKN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_6 N_28 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M20 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_6 N_5 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_4 N_5 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_4 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_6 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M40 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfbfb2
* SPICE INPUT		Wed Jul 10 13:34:34 2019	dfbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb1
.subckt dfbrb1 VDD QN Q GND RN SN CK D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_6 N_26 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CK GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_6 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_8 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M13 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M14 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M17 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_6 N_5 VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_6 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M34 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M37 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfbrb1
* SPICE INPUT		Wed Jul 10 13:34:42 2019	dfbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb2
.subckt dfbrb2 VDD QN Q GND RN SN CK D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_6 N_26 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CK GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_6 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_8 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M20 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_6 N_5 VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_6 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M40 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfbrb2
* SPICE INPUT		Wed Jul 10 13:34:49 2019	dfbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq1
.subckt dfbrq1 VDD Q GND RN D SN CK
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 SN GND GND mn5  l=0.5u w=0.58u m=1
M3 N_26 N_3 Q GND mn5  l=0.5u w=0.58u m=1
M4 N_26 N_8 Q GND mn5  l=0.5u w=0.58u m=1
M5 N_25 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_3 N_25 GND mn5  l=0.5u w=0.5u m=1
M7 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_5 N_30 GND mn5  l=0.5u w=0.5u m=1
M10 N_31 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M13 N_21 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_21 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_29 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M17 N_6 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M18 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M21 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M23 Q N_3 N_18 VDD mp5  l=0.42u w=0.76u m=1
M24 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_18 N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.5u m=1
M27 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M31 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M34 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M36 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M37 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M38 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfbrq1
* SPICE INPUT		Wed Jul 10 13:34:56 2019	dfbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq2
.subckt dfbrq2 VDD Q GND SN D RN CK
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_24 SN GND GND mn5  l=0.5u w=0.72u m=1
M6 N_24 N_3 Q GND mn5  l=0.5u w=0.72u m=1
M7 Q N_8 N_24 GND mn5  l=0.5u w=0.72u m=1
M8 N_23 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_3 N_23 GND mn5  l=0.5u w=0.5u m=1
M10 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M11 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_8 N_5 N_30 GND mn5  l=0.5u w=0.5u m=1
M13 N_31 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M14 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_19 SN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_19 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_19 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M18 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_29 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M20 N_6 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M21 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M26 Q N_3 N_18 VDD mp5  l=0.42u w=0.96u m=1
M27 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_18 N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.5u m=1
M30 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M34 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M40 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
.ends dfbrq2
* SPICE INPUT		Wed Jul 10 13:35:03 2019	dfcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb1
.subckt dfcfb1 GND QN Q VDD RN D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_14 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_15 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_8 N_4 N_16 GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M18 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M19 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_22 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M23 N_21 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M24 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M29 N_25 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M33 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M36 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfcfb1
* SPICE INPUT		Wed Jul 10 13:35:11 2019	dfcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb2
.subckt dfcfb2 GND QN Q VDD RN D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_14 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_15 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_8 N_4 N_16 GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M18 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M19 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_22 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M23 N_21 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M24 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M29 N_25 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M33 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M36 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfcfb2
* SPICE INPUT		Wed Jul 10 13:35:18 2019	dfcfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfq1
.subckt dfcfq1 GND Q VDD CKN D RN
M1 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_16 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_16 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_15 GND mn5  l=0.5u w=0.5u m=1
M9 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_14 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_13 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_25 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_24 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 N_24 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_25 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_23 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_22 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_22 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_21 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_20 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_20 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcfq1
* SPICE INPUT		Wed Jul 10 13:35:25 2019	dfcfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfq2
.subckt dfcfq2 GND Q VDD CKN D RN
M1 N_16 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_16 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 N_4 N_15 GND mn5  l=0.5u w=0.5u m=1
M5 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M7 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_14 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_13 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_35 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_35 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_34 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M21 N_36 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M22 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M24 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M25 N_34 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_33 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_33 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_32 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_31 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M30 N_32 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M31 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_36 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfcfq2
* SPICE INPUT		Wed Jul 10 13:35:32 2019	dfcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb1
.subckt dfcrb1 VDD QN Q GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_26 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_26 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M10 N_25 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_24 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_24 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_23 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_23 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M27 N_17 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_14 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M33 N_15 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M34 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrb1
* SPICE INPUT		Wed Jul 10 13:35:39 2019	dfcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb2
.subckt dfcrb2 GND QN Q VDD CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_17 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_5 N_16 GND mn5  l=0.5u w=0.5u m=1
M10 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_25 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M27 N_24 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_21 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M33 N_22 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M34 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrb2
* SPICE INPUT		Wed Jul 10 13:35:47 2019	dfcrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrn1
.subckt dfcrn1 VDD QN GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_34 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_34 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_33 GND mn5  l=0.5u w=0.5u m=1
M8 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_17 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrn1
* SPICE INPUT		Wed Jul 10 13:35:54 2019	dfcrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrn2
.subckt dfcrn2 VDD QN GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_23 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_22 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_22 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_21 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_21 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_17 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrn2
* SPICE INPUT		Wed Jul 10 13:36:01 2019	dfcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq1
.subckt dfcrq1 VDD Q GND CK D RN
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 Q N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_9 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_18 N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.52u m=1
M21 N_18 N_3 Q VDD mp5  l=0.42u w=0.76u m=1
M22 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrq1
* SPICE INPUT		Wed Jul 10 13:36:08 2019	dfcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq2
.subckt dfcrq2 VDD Q GND RN D CK
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_18 N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_18 N_3 Q VDD mp5  l=0.42u w=0.96u m=1
M21 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrq2
* SPICE INPUT		Wed Jul 10 13:36:15 2019	dfnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb1
.subckt dfnfb1 VDD QN Q GND D CKN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_5 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnfb1
* SPICE INPUT		Wed Jul 10 13:36:22 2019	dfnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb2
.subckt dfnfb2 VDD QN Q GND CKN D
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_5 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M15 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M18 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfnfb2
* SPICE INPUT		Wed Jul 10 13:36:30 2019	dfnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb1
.subckt dfnrb1 VDD QN Q GND CK D
M1 QN N_10 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_10 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_32 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_31 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_30 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M11 N_6 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_10 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_10 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 VDD N_10 N_16 VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M20 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M21 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M25 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M26 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfnrb1
* SPICE INPUT		Wed Jul 10 13:36:37 2019	dfnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb2
.subckt dfnrb2 VDD QN Q GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M17 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfnrb2
* SPICE INPUT		Wed Jul 10 13:36:44 2019	dfnrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrn1
.subckt dfnrn1 VDD QN GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrn1
* SPICE INPUT		Wed Jul 10 13:36:51 2019	dfnrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrn2
.subckt dfnrn2 VDD QN GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrn2
* SPICE INPUT		Wed Jul 10 13:36:58 2019	dfnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq1
.subckt dfnrq1 VDD Q GND CK D
M1 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrq1
* SPICE INPUT		Wed Jul 10 13:37:05 2019	dfnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq2
.subckt dfnrq2 VDD Q GND CK D
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrq2
* SPICE INPUT		Wed Jul 10 13:37:13 2019	dfpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb1
.subckt dfpfb1 VDD Q QN GND CKN D SN
M1 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_36 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_36 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_33 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_33 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfpfb1
* SPICE INPUT		Wed Jul 10 13:37:20 2019	dfpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb2
.subckt dfpfb2 VDD Q QN GND CKN D SN
M1 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_36 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_36 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M10 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_33 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M32 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M33 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfpfb2
* SPICE INPUT		Wed Jul 10 13:37:27 2019	dfprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb1
.subckt dfprb1 VDD Q QN GND SN D CK
M1 N_4 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_33 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_33 N_12 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_34 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_34 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_10 GND GND mn5  l=0.5u w=0.58u m=1
M7 QN N_8 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_10 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_35 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_35 SN N_6 GND mn5  l=0.5u w=0.5u m=1
M11 N_38 N_7 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_36 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_4 N_36 GND mn5  l=0.5u w=0.5u m=1
M14 N_37 N_12 N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_37 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_38 SN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_12 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_4 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_15 N_12 N_5 VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 Q N_10 VDD VDD mp5  l=0.42u w=0.76u m=1
M24 QN N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M25 N_10 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_6 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_6 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_12 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_17 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M32 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_8 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_12 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprb1
* SPICE INPUT		Wed Jul 10 13:37:34 2019	dfprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb2
.subckt dfprb2 VDD Q QN GND SN D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_34 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_34 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M10 N_35 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_4 N_35 GND mn5  l=0.5u w=0.5u m=1
M12 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M13 N_36 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M14 N_36 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_37 SN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_37 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_4 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_7 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_7 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M30 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M32 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfprb2
* SPICE INPUT		Wed Jul 10 13:37:41 2019	dfprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq1
.subckt dfprq1 VDD Q GND CK D SN
M1 Q N_8 N_27 GND mn5  l=0.5u w=0.58u m=1
M2 N_27 SN GND GND mn5  l=0.5u w=0.58u m=1
M3 N_33 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 N_33 GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_32 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_31 GND mn5  l=0.5u w=0.5u m=1
M8 N_31 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_30 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_30 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M19 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_9 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_14 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_7 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_7 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_11 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprq1
* SPICE INPUT		Wed Jul 10 13:37:48 2019	dfprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq2
.subckt dfprq2 VDD Q GND CK D SN
M1 Q N_10 N_29 GND mn5  l=0.5u w=0.72u m=1
M2 N_29 SN GND GND mn5  l=0.5u w=0.72u m=1
M3 N_35 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_34 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 N_10 N_35 GND mn5  l=0.5u w=0.5u m=1
M6 N_34 N_5 N_10 GND mn5  l=0.5u w=0.5u m=1
M7 N_10 N_4 N_33 GND mn5  l=0.5u w=0.5u m=1
M8 N_33 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_32 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_32 N_7 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M13 N_30 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_30 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_11 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_16 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_11 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_15 N_5 N_10 VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_9 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_13 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_5 N_7 VDD mp5  l=0.42u w=0.5u m=1
M29 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_4 N_10 VDD mp5  l=0.42u w=0.5u m=1
M31 VDD N_5 N_4 VDD mp5  l=0.42u w=0.5u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprq2