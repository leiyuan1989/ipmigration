

.SUBCKT TLATNCAX12MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_3 XI14_n1__3 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_3 nmin c XI14_n1__3 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_4 nmin c XI14_n1__4 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_4 XI14_n1__4 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_5 XI14_n1__5 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_5 nmin c XI14_n1__5 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=2.9e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=2.9e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_2 ECK nmin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_3 ECK nmin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=7.9e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_3 XI14_p1__3 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPOEN_3 nmin cn XI14_p1__3 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPOEN_4 nmin cn XI14_p1__4 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_4 XI14_p1__4 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_5 XI14_p1__5 E VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPOEN_5 nmin cn XI14_p1__5 VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK nmin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK nmin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK nmin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX16MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_3 XI14_n1__3 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_3 nmin c XI14_n1__3 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_4 nmin c XI14_n1__4 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_4 XI14_n1__4 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_5 XI14_n1__5 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_5 nmin c XI14_n1__5 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_2 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_3 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=8.1e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_3 XI14_p1__3 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPOEN_3 nmin cn XI14_p1__3 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPOEN_4 nmin cn XI14_p1__4 VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_4 XI14_p1__4 E VDD VNW p12 l=1.3e-07 w=7.2e-07
mXI14_MXPA1_5 XI14_p1__5 E VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPOEN_5 nmin cn XI14_p1__5 VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.7e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK nmin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK nmin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK nmin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 ECK nmin XI1_p1__7 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_7 XI1_p1__7 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_8 XI1_p1__8 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 ECK nmin XI1_p1__8 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX20MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_3 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_4 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_5 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1_3 XI14_n1__3 E VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNOE_3 nmin c XI14_n1__3 VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNOE_4 nmin c XI14_n1__4 VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1_4 XI14_n1__4 E VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1_5 XI14_n1__5 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_5 nmin c XI14_n1__5 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_6 nmin c XI14_n1__6 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_6 XI14_n1__6 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1_7 XI14_n1__7 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_7 nmin c XI14_n1__7 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_2 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_3 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA2_4 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_4 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_4 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_5 c CK VDD VNW p12 l=1.3e-07 w=8.1e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPA1_3 XI14_p1__3 E VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPOEN_3 nmin cn XI14_p1__3 VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPOEN_4 nmin cn XI14_p1__4 VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPA1_4 XI14_p1__4 E VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI14_MXPA1_5 XI14_p1__5 E VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI14_MXPOEN_5 nmin cn XI14_p1__5 VNW p12 l=1.3e-07 w=7.1e-07
mXI14_MXPOEN_6 nmin cn XI14_p1__6 VNW p12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1_6 XI14_p1__6 E VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1_7 XI14_p1__7 E VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI14_MXPOEN_7 nmin cn XI14_p1__7 VNW p12 l=1.3e-07 w=6.8e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.8e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK nmin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK nmin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK nmin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 ECK nmin XI1_p1__7 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_7 XI1_p1__7 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_8 XI1_p1__8 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 ECK nmin XI1_p1__8 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_9 ECK nmin XI1_p1__9 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_9 XI1_p1__9 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_10 XI1_p1__10 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_10 ECK nmin XI1_p1__10 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX2MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX3MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.8e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX4MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=3e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=4.3e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=4.3e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=5.9e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=5.9e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX6MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=5.6e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNCAX8MTR ECK VDD VNW VPW VSS CK E
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI14_MXNA1_2 XI14_n1__2 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE_2 nmin c XI14_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNOE nmin c XI14_n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI14_MXNA1 XI14_n1 E VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNOE nmin cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK nmin VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1_2 ECK nmin VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI14_MXPA1_2 XI14_p1__2 E VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPOEN_2 nmin cn XI14_p1__2 VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPOEN nmin cn XI14_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPA1 XI14_p1 E VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI13_MXPOEN nmin c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m nmin VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK nmin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK nmin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK nmin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK nmin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNSRX1MTR Q QN VDD VNW VPW VSS D GN RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=4e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=3.7e-07
MXN7 net048 D VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN6 net052 RN net048 VPW n12 l=1.3e-07 w=5.3e-07
MX_t13 pm c net052 VPW n12 l=1.3e-07 w=5.3e-07
MX_t2 pm cn net98 VPW n12 l=1.3e-07 w=2.8e-07
MXN8 net98 RN net101 VPW n12 l=1.3e-07 w=2.8e-07
MXN9 VSS m net101 VPW n12 l=1.3e-07 w=2.8e-07
mX_g4_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 c GN VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI47_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI46_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP11 pm nms net61 VNW p12 l=1.3e-07 w=6.3e-07
MX_t14 net61 RN VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t9 net083 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP9 net075 nms net083 VNW p12 l=1.3e-07 w=6.4e-07
MXP10 pm cn net075 VNW p12 l=1.3e-07 w=6.4e-07
MXP13 pm c net70 VNW p12 l=1.3e-07 w=3.2e-07
MXP12 net70 nms net67 VNW p12 l=1.3e-07 w=3.2e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3.2e-07
mX_g4_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 c GN VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI47_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI46_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TLATNSRX2MTR Q QN VDD VNW VPW VSS D GN RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=6.2e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN7_2 net048__2 D VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN6_2 net052__2 RN net048__2 VPW n12 l=1.3e-07 w=5.3e-07
MX_t13_2 pm c net052__2 VPW n12 l=1.3e-07 w=5e-07
MX_t13 pm c net052 VPW n12 l=1.3e-07 w=4.1e-07
MXN6 net052 RN net048 VPW n12 l=1.3e-07 w=2.6e-07
MXN7 net048 D VSS VPW n12 l=1.3e-07 w=3.7e-07
MX_t2 pm cn net98 VPW n12 l=1.3e-07 w=2.8e-07
MXN8 net98 RN net101 VPW n12 l=1.3e-07 w=2.8e-07
MXN9 VSS m net101 VPW n12 l=1.3e-07 w=2.8e-07
mX_g4_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g5_MXNA1 c GN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI48_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI46_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=7.5e-07
MXP18 pm nms net61 VNW p12 l=1.3e-07 w=8.8e-07
MX_t14 net61 RN VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t9_2 net083__2 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP16_2 net075__2 nms net083__2 VNW p12 l=1.3e-07 w=6.4e-07
MXP17_2 pm cn net075__2 VNW p12 l=1.3e-07 w=6.4e-07
MXP17 pm cn net075 VNW p12 l=1.3e-07 w=6.4e-07
MXP16 net075 nms net083 VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 net083 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 pm c net70 VNW p12 l=1.3e-07 w=3.2e-07
MXP12 net70 nms net67 VNW p12 l=1.3e-07 w=3.2e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3.2e-07
mX_g4_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g5_MXPA1 c GN VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.4e-07
mXI48_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI46_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNSRX4MTR Q QN VDD VNW VPW VSS D GN RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=5.9e-07
mX_g3_MXNA1_2 nms SN VSS VPW n12 l=1.3e-07 w=5.8e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t6_2 pm nms VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN7_2 net048__2 D VSS VPW n12 l=1.3e-07 w=5.1e-07
MXN6_2 net052__2 RN net048__2 VPW n12 l=1.3e-07 w=5.1e-07
MX_t13_2 pm c net052__2 VPW n12 l=1.3e-07 w=5e-07
MX_t13 pm c net052 VPW n12 l=1.3e-07 w=4.1e-07
MXN6 net052 RN net048 VPW n12 l=1.3e-07 w=2.6e-07
MXN7 net048 D VSS VPW n12 l=1.3e-07 w=3.9e-07
MX_t2 pm cn net98 VPW n12 l=1.3e-07 w=2.8e-07
MXN8 net98 RN net101 VPW n12 l=1.3e-07 w=2.8e-07
MXN9 VSS m net101 VPW n12 l=1.3e-07 w=2.8e-07
mX_g4_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g5_MXNA1 c GN VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI50_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI50_MXNA1_2 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI49_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI49_MXNA1_2 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1_2 nms SN VDD VNW p12 l=1.3e-07 w=7.2e-07
MXP18 pm nms net61 VNW p12 l=1.3e-07 w=8.8e-07
MX_t14 net61 RN VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t9_2 net083__2 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP16_2 net075__2 nms net083__2 VNW p12 l=1.3e-07 w=6.4e-07
MXP17_2 pm cn net075__2 VNW p12 l=1.3e-07 w=6.4e-07
MXP17 pm cn net075 VNW p12 l=1.3e-07 w=6.4e-07
MXP16 net075 nms net083 VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 net083 D VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 pm c net70 VNW p12 l=1.3e-07 w=3.2e-07
MXP12 net70 nms net67 VNW p12 l=1.3e-07 w=3.2e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3.2e-07
mX_g4_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g5_MXPA1 c GN VDD VNW p12 l=1.3e-07 w=8.2e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI50_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI50_MXPA1_2 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI49_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI49_MXPA1_2 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX12MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g6_MXNA1_3 c CK VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g6_MXNA1_4 c CK VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g7_MXNA1_2 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_4 X_g3_n1__4 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_4 csetin c X_g3_n1__4 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_5 csetin c X_g3_n1__5 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_5 X_g3_n1__5 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_6 X_g3_n1__6 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_6 csetin c X_g3_n1__6 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1_4 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=7.9e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=8.7e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g7_MXPA1_2 setin nmsetin VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1_4 X_g3_p1__4 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_4 csetin cn X_g3_p1__4 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_5 csetin cn X_g3_p1__5 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1_5 X_g3_p1__5 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1_6 X_g3_p1__6 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN_6 csetin cn X_g3_p1__6 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.8e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.8e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK csetin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK csetin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX16MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_3 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_4 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_5 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g5_MXNA1_2 cn c VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g8_MXNA1_2 nmsetin E VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g8_MXNA2_2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g7_MXNA1_2 setin nmsetin VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g7_MXNA1_3 setin nmsetin VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=4.95e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=4.95e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=4.95e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=4.95e-07
mX_g3_MXNA1_4 X_g3_n1__4 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_4 csetin c X_g3_n1__4 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_5 csetin c X_g3_n1__5 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1_5 X_g3_n1__5 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1_6 X_g3_n1__6 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_6 csetin c X_g3_n1__6 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_7 csetin c X_g3_n1__7 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1_7 X_g3_n1__7 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1_8 X_g3_n1__8 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE_8 csetin c X_g3_n1__8 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.85e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.85e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=5e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_3 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_4 ECK csetin VSS VPW n12 l=1.3e-07 w=2e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g6_MXPA1_4 c CK VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g6_MXPA1_5 c CK VDD VNW p12 l=1.3e-07 w=7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g5_MXPA1_2 cn c VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g8_MXPA2_2 X_g8_p1__2 SE VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1_2 nmsetin E X_g8_p1__2 VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g7_MXPA1_2 setin nmsetin VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g7_MXPA1_3 setin nmsetin VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=4.65e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=4.65e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=4.65e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=4.65e-07
mX_g3_MXPA1_4 X_g3_p1__4 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_4 csetin cn X_g3_p1__4 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_5 csetin cn X_g3_p1__5 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1_5 X_g3_p1__5 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1_6 X_g3_p1__6 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_6 csetin cn X_g3_p1__6 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_7 csetin cn X_g3_p1__7 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1_7 X_g3_p1__7 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1_8 X_g3_p1__8 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN_8 csetin cn X_g3_p1__8 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=4.95e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=4.95e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK csetin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK csetin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK csetin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 ECK csetin XI1_p1__7 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_7 XI1_p1__7 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX20MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_3 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_4 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_5 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g5_MXNA1_2 cn c VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g8_MXNA1_2 nmsetin E VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g8_MXNA2_2 nmsetin SE VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g7_MXNA1_2 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g7_MXNA1_3 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=7.2e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=7.2e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNOE_4 csetin c X_g3_n1__4 VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_4 X_g3_n1__4 setin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_5 X_g3_n1__5 setin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNOE_5 csetin c X_g3_n1__5 VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNOE_6 csetin c X_g3_n1__6 VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_6 X_g3_n1__6 setin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_7 X_g3_n1__7 setin VSS VPW n12 l=1.3e-07 w=4.4e-07
mX_g3_MXNOE_7 csetin c X_g3_n1__7 VPW n12 l=1.3e-07 w=4.4e-07
mX_g3_MXNOE_8 csetin c X_g3_n1__8 VPW n12 l=1.3e-07 w=4.4e-07
mX_g3_MXNA1_8 X_g3_n1__8 setin VSS VPW n12 l=1.3e-07 w=4.4e-07
mX_g3_MXNA1_9 X_g3_n1__9 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_9 csetin c X_g3_n1__9 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA2_3 ECK c VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA1_3 ECK csetin VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_3 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_4 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_5 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g5_MXPA1_2 cn c VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g8_MXPA2_2 X_g8_p1__2 SE VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1_2 nmsetin E X_g8_p1__2 VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=8.1e-07
mX_g7_MXPA1_2 setin nmsetin VDD VNW p12 l=1.3e-07 w=8.1e-07
mX_g7_MXPA1_3 setin nmsetin VDD VNW p12 l=1.3e-07 w=8e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=8e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=8e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_4 csetin cn X_g3_p1__4 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_4 X_g3_p1__4 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_5 X_g3_p1__5 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_5 csetin cn X_g3_p1__5 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_6 csetin cn X_g3_p1__6 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_6 X_g3_p1__6 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_7 X_g3_p1__7 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_7 csetin cn X_g3_p1__7 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_8 csetin cn X_g3_p1__8 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_8 X_g3_p1__8 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1_9 X_g3_p1__9 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN_9 csetin cn X_g3_p1__9 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 ECK csetin XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 ECK csetin XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 ECK csetin XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_7 XI1_p1__7 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 ECK csetin XI1_p1__7 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 ECK csetin XI1_p1__8 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_8 XI1_p1__8 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_9 XI1_p1__9 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_9 ECK csetin XI1_p1__9 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX2MTR ECK VDD VNW VPW VSS CK E SE
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=3e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=3e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX3MTR ECK VDD VNW VPW VSS CK E SE
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=3e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=3e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX4MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=3e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=3e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=3.2e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX6MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=6e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=3e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=3e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=4.4e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=4.6e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.3e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.3e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.9e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=8.8e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNTSCAX8MTR ECK VDD VNW VPW VSS CK E SE
mX_g6_MXNA1 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXNA1_2 c CK VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXNA1 cn c VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g8_MXNA1 nmsetin E VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g8_MXNA2 nmsetin SE VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g7_MXNA1 setin nmsetin VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g7_MXNA1_2 setin nmsetin VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g3_MXNA1_2 X_g3_n1__2 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_2 csetin c X_g3_n1__2 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_3 csetin c X_g3_n1__3 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_3 X_g3_n1__3 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1_4 X_g3_n1__4 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE_4 csetin c X_g3_n1__4 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNOE csetin c X_g3_n1 VPW n12 l=1.3e-07 w=4.3e-07
mX_g3_MXNA1 X_g3_n1 setin VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g2_MXNA1 m csetin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNOE csetin cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 ECK c VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI1_MXNA1 ECK csetin VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI1_MXNA1_2 ECK csetin VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI1_MXNA2_2 ECK c VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g6_MXPA1 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1_2 c CK VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g5_MXPA1 cn c VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g8_MXPA1 nmsetin E X_g8_p1 VNW p12 l=1.3e-07 w=5.9e-07
mX_g8_MXPA2 X_g8_p1 SE VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g7_MXPA1 setin nmsetin VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g7_MXPA1_2 setin nmsetin VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1_2 X_g3_p1__2 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN_2 csetin cn X_g3_p1__2 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN_3 csetin cn X_g3_p1__3 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPA1_3 X_g3_p1__3 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPA1_4 X_g3_p1__4 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN_4 csetin cn X_g3_p1__4 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPOEN csetin cn X_g3_p1 VNW p12 l=1.3e-07 w=5.9e-07
mX_g3_MXPA1 X_g3_p1 setin VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g2_MXPA1 m csetin VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN csetin c XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2_2 XI1_p1__2 c VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 ECK csetin XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 ECK csetin XI1_p1__3 VNW p12 l=1.3e-07 w=9e-07
mXI1_MXPA2_3 XI1_p1__3 c VDD VNW p12 l=1.3e-07 w=9e-07
mXI1_MXPA2_4 XI1_p1__4 c VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI1_MXPA1_4 ECK csetin XI1_p1__4 VNW p12 l=1.3e-07 w=8.8e-07
mXI1_MXPA1 ECK csetin XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 c VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNX1MTR Q QN VDD VNW VPW VSS D GN
mX_g5_MXNA1 cn GN VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 D VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI1_MXNOE pm cn XI1_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI21_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1 cn GN VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI1_MXPOEN pm c XI1_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI21_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TLATNX2MTR Q QN VDD VNW VPW VSS D GN
mX_g5_MXNA1 cn GN VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI1_MXNA1 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNOE pm cn XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI22_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 cn GN VDD VNW p12 l=1.3e-07 w=3.8e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI1_MXPA1 XI1_p1 D VDD VNW p12 l=1.3e-07 w=7e-07
mXI1_MXPOEN pm c XI1_p1 VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI22_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATNX4MTR Q QN VDD VNW VPW VSS D GN
mX_g5_MXNA1 cn GN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI1_MXNA1 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNOE pm cn XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI24_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_2 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 cn GN VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 D VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI1_MXPOEN pm c XI1_p1 VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI24_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_2 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATSRX1MTR Q QN VDD VNW VPW VSS D G RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=3.1e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN1 net84 D VSS VPW n12 l=1.3e-07 w=3.9e-07
MXN0 net80 RN net84 VPW n12 l=1.3e-07 w=3.9e-07
MX_t13 pm c net80 VPW n12 l=1.3e-07 w=3.9e-07
MX_t2 pm cn net100 VPW n12 l=1.3e-07 w=2.6e-07
MXN2 net100 RN net105 VPW n12 l=1.3e-07 w=2.6e-07
MXN3 VSS m net105 VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3e-07
mX_g0_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP1 pm cn net47 VNW p12 l=1.3e-07 w=5.2e-07
MXP0 net47 nms net55 VNW p12 l=1.3e-07 w=5.2e-07
MX_t9 net55 D VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t14 net63 RN VDD VNW p12 l=1.3e-07 w=4.7e-07
MXP2 pm nms net63 VNW p12 l=1.3e-07 w=4.7e-07
MXP4 pm c net71 VNW p12 l=1.3e-07 w=3.2e-07
MXP3 net71 nms net67 VNW p12 l=1.3e-07 w=3.2e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3.2e-07
mX_g5_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g0_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TLATSRX2MTR Q QN VDD VNW VPW VSS D G RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=4.5e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=4e-07
MXN5 net84 D VSS VPW n12 l=1.3e-07 w=4.1e-07
MXN4 net80 RN net84 VPW n12 l=1.3e-07 w=4.1e-07
MX_t13 pm c net80 VPW n12 l=1.3e-07 w=4.1e-07
MX_t2 pm cn net100 VPW n12 l=1.3e-07 w=2.6e-07
MXN2 net100 RN net105 VPW n12 l=1.3e-07 w=2.6e-07
MXN3 VSS m net105 VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=2e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3e-07
mXI46_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP1 pm cn net47 VNW p12 l=1.3e-07 w=5.7e-07
MXP5 net47 nms net55 VNW p12 l=1.3e-07 w=8.6e-07
MX_t9 net55 D VDD VNW p12 l=1.3e-07 w=8.6e-07
MX_t14 net63 RN VDD VNW p12 l=1.3e-07 w=7.3e-07
MXP6 pm nms net63 VNW p12 l=1.3e-07 w=7.3e-07
MXP8 pm c net71 VNW p12 l=1.3e-07 w=3e-07
MXP7 net71 nms net67 VNW p12 l=1.3e-07 w=3e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI46_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATSRX4MTR Q QN VDD VNW VPW VSS D G RN SN
mX_g3_MXNA1 nms SN VSS VPW n12 l=1.3e-07 w=6.3e-07
MX_t6 pm nms VSS VPW n12 l=1.3e-07 w=4e-07
MXN5 net84 D VSS VPW n12 l=1.3e-07 w=4.1e-07
MXN4 net80 RN net84 VPW n12 l=1.3e-07 w=4.1e-07
MX_t13 pm c net80 VPW n12 l=1.3e-07 w=4.1e-07
MX_t2 pm cn net100 VPW n12 l=1.3e-07 w=2.6e-07
MXN2 net100 RN net105 VPW n12 l=1.3e-07 w=2.6e-07
MXN3 VSS m net105 VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g4_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=3.4e-07
mX_g2_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI46_MXNA1 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI46_MXNA1_2 Q pm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 nms SN VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP1 pm cn net47 VNW p12 l=1.3e-07 w=5.7e-07
MXP5 net47 nms net55 VNW p12 l=1.3e-07 w=8.6e-07
MX_t9 net55 D VDD VNW p12 l=1.3e-07 w=8.6e-07
MX_t14 net63 RN VDD VNW p12 l=1.3e-07 w=7.3e-07
MXP6 pm nms net63 VNW p12 l=1.3e-07 w=7.3e-07
MXP8 pm c net71 VNW p12 l=1.3e-07 w=3e-07
MXP7 net71 nms net67 VNW p12 l=1.3e-07 w=3e-07
MX_t5 VDD m net67 VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g4_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=4.2e-07
mX_g2_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI46_MXPA1 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI46_MXPA1_2 Q pm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATX1MTR Q QN VDD VNW VPW VSS D G
mX_g6_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g5_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g3_MXNOE net52 c X_g3_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI5_MXNOE net52 cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m net52 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI25_MXNA1 Q net52 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g5_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g3_MXPOEN net52 cn X_g3_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI5_MXPOEN net52 c XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 m net52 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI25_MXPA1 Q net52 VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TLATX2MTR Q QN VDD VNW VPW VSS D G
mX_g6_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=6.5e-07
mX_g3_MXNOE net52 c X_g3_n1 VPW n12 l=1.3e-07 w=6.5e-07
mXI5_MXNOE net52 cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m net52 VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI25_MXNA1 Q net52 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=8e-07
mX_g3_MXPOEN net52 cn X_g3_p1 VNW p12 l=1.3e-07 w=8e-07
mXI5_MXPOEN net52 c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 m net52 VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI25_MXPA1 Q net52 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TLATX4MTR Q QN VDD VNW VPW VSS D G
mX_g6_MXNA1 cn G VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g5_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNOE net52 c X_g3_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI5_MXNOE net52 cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 m net52 VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI26_MXNA1 Q net52 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI26_MXNA1_2 Q net52 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN m VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g6_MXPA1 cn G VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g3_MXPOEN net52 cn X_g3_p1 VNW p12 l=1.3e-07 w=6.9e-07
mXI5_MXPOEN net52 c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 m net52 VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI26_MXPA1 Q net52 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI26_MXPA1_2 Q net52 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN m VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


***********************************************************



.SUBCKT DFFHQNX1MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFHQNX2MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQNX4MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=6.1e-07
.ends


.SUBCKT DFFHQNX8MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_3 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_4 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_3 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_4 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQX1MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=3.4e-07
MXN3 net87 cn VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP4 net061 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm nmin net62 VNW p12 l=1.3e-07 w=4.1e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.4e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFHQX2MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=4.8e-07
MXN4 net87 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP6 net061 c cn VNW p12 l=1.3e-07 w=4.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP7 pm nmin net62 VNW p12 l=1.3e-07 w=5.9e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.4e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQX4MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net87 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP8 net061 c cn VNW p12 l=1.3e-07 w=7.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP9 pm nmin net62 VNW p12 l=1.3e-07 w=8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI36_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQX8MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=4.4e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net87 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=7.3e-07
MXP10 net061 c cn VNW p12 l=1.3e-07 w=7.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=8.5e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP9 pm nmin net62 VNW p12 l=1.3e-07 w=8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI36_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=7.3e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHX1MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net42 cn VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP5 net63 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP2 net53 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP6 pm nmin net53 VNW p12 l=1.3e-07 w=4.4e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.9e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFHX2MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=5.1e-07
MXN4 net42 cn VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP7 net63 c cn VNW p12 l=1.3e-07 w=4.6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8e-07
MXP8 net53 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP10 pm nmin net53 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI32_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.1e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT DFFHX4MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=7e-07
MXN5 net42 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP11 net63 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP8 net53 c VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP12 pm nmin net53 VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI32_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT DFFHX8MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=7e-07
MXN5 net42 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP11 net63 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP8 net53 c VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP12 pm nmin net53 VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI32_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT DFFNHX1MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=4.3e-07
MXN2 net67 cn VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net56 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=6.8e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP3 pm net150 net42 VNW p12 l=1.3e-07 w=3.3e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.8e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNHX2MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=6.1e-07
MXN3 net67 cn VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net56 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1_2 cn nckn VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP4 pm net150 net42 VNW p12 l=1.3e-07 w=4.6e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNHX4MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=5.4e-07
MXN3 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN3_2 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 pm net150 net67 VPW n12 l=1.3e-07 w=5.4e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI37_MXNOE_2 bm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP5 net56 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=6.6e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g10_MXPA1_2 cn nckn VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 pm net150 net42 VNW p12 l=1.3e-07 w=6.9e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI37_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mXI52_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNHX8MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=5e-07
mX_g13_MXNA1_2 net150 D VSS VPW n12 l=1.3e-07 w=5e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=7.4e-07
MXN3 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN3_2 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 pm net150 net67 VPW n12 l=1.3e-07 w=5.7e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI37_MXNOE_2 bm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP7 net56 cn c VNW p12 l=1.3e-07 w=6.4e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g13_MXPA1_2 net150 D VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g10_MXPA1_2 cn nckn VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 pm net150 net42 VNW p12 l=1.3e-07 w=6.9e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI37_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mXI52_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI52_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI52_MXPA1_5 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNSRHX1MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS SN net68 VPW n12 l=1.3e-07 w=4.3e-07
MXN11 net68 cn net72 VPW n12 l=1.3e-07 w=4.3e-07
MXN0 pm nmin net72 VPW n12 l=1.3e-07 w=4.3e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 m pm net80 VPW n12 l=1.3e-07 w=4.5e-07
MXN13 VSS RN net80 VPW n12 l=1.3e-07 w=4.5e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
MXN7 bm cn net91 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net91 RN net88 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net88 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net152 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP13 net152 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmin net118 VNW p12 l=1.3e-07 w=3.3e-07
MXP9 net118 c VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=4.8e-07
MXP1 net142 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net142 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.8e-07
MXP16 bm nmset net154 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net154 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP18 bm c net110 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net110 nmset net114 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net114 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT DFFNSRHX2MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS SN net70 VPW n12 l=1.3e-07 w=6e-07
MXN16 net70 cn net66 VPW n12 l=1.3e-07 w=6e-07
MXN0 pm nmin net66 VPW n12 l=1.3e-07 w=6e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 m pm net78 VPW n12 l=1.3e-07 w=6.3e-07
MXN18 VSS RN net78 VPW n12 l=1.3e-07 w=6.3e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.6e-07
MXN7 bm cn net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net89 RN net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net154 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP13 net154 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 pm nmin net120 VNW p12 l=1.3e-07 w=4.6e-07
MXP9 net120 c VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP1 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP20 bm nmset net104 VNW p12 l=1.3e-07 w=2.8e-07
MXP4 net104 RN VDD VNW p12 l=1.3e-07 w=2.8e-07
MXP18 bm c net112 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net112 nmset net116 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net116 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFNSRHX4MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=3e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN20 VSS SN net67 VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net67 cn net71 VPW n12 l=1.3e-07 w=7.5e-07
MXN0 pm nmin net71 VPW n12 l=1.3e-07 w=7.5e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 m pm net79 VPW n12 l=1.3e-07 w=8.4e-07
MXN21 VSS RN net79 VPW n12 l=1.3e-07 w=8.4e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN7 bm cn net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net90 RN net87 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net87 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net155 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP21 net155 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.6e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP22 pm nmin net121 VNW p12 l=1.3e-07 w=6.9e-07
MXP9 net121 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP11_2 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP1 net145 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net145 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP23 bm nmset net105 VNW p12 l=1.3e-07 w=3.6e-07
MXP4 net105 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP18 bm c net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net113 nmset net117 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net117 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFNSRHX8MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g10_MXNA1_2 cn nck VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN20 VSS SN net66 VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net66 cn net70 VPW n12 l=1.3e-07 w=7.5e-07
MXN0 pm nmin net70 VPW n12 l=1.3e-07 w=7.5e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=2.5e-07
MXN4 m pm net78 VPW n12 l=1.3e-07 w=8.7e-07
MXN22 VSS RN net78 VPW n12 l=1.3e-07 w=8.7e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN7 bm cn net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net89 RN net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=3e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP2 net154 CKN VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP24 net154 cn c VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g10_MXPA1_2 cn nck VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=1.03e-06
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP22 pm nmin net120 VNW p12 l=1.3e-07 w=6.9e-07
MXP9 net120 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP11_2 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP1 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP25 bm nmset net104 VNW p12 l=1.3e-07 w=3.5e-07
MXP4 net104 RN VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP18 bm c net112 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net112 nmset net116 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net116 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQNX1MTR QN VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE nm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE nm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN nm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN nm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFQNX2MTR QN VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE nm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE nm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN nm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN nm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQNX4MTR QN VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE nm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE nm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN nm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN nm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQX1MTR Q VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI6_MXNOE ns c XI6_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI7_MXNOE ns cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI6_MXPOEN ns cn XI6_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI7_MXPOEN ns c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFQX2MTR Q VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI6_MXNOE ns c XI6_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI7_MXNOE ns cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI6_MXPOEN ns cn XI6_p1 VNW p12 l=1.3e-07 w=4.9e-07
mXI7_MXPOEN ns c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g1_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQX4MTR Q VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI6_MXNOE ns c XI6_n1 VPW n12 l=1.3e-07 w=4.2e-07
mXI7_MXNOE ns cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI6_MXPOEN ns cn XI6_p1 VNW p12 l=1.3e-07 w=6.1e-07
mXI7_MXPOEN ns c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g1_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRHQX1MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net89 cn VSS VPW n12 l=1.3e-07 w=3.5e-07
MXN2 pm nmin net89 VPW n12 l=1.3e-07 w=3.5e-07
MXN3 pm c net66 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net66 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net73 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
MXN11 m pm net73 VPW n12 l=1.3e-07 w=4.9e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=3.7e-07
MXN7 bm cn net85 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net85 RN net82 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net82 VPW n12 l=1.3e-07 w=1.5e-07
mXI52_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net126 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP11 net126 c cn VNW p12 l=1.3e-07 w=4.2e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP2 net134 c VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP12 pm nmin net134 VNW p12 l=1.3e-07 w=4.2e-07
MXP14 pm cn net104 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 VDD m net104 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.3e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP16 bm c net120 VNW p12 l=1.3e-07 w=2.3e-07
MXP15 VDD s net120 VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFRHQX2MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net90 cn VSS VPW n12 l=1.3e-07 w=5.1e-07
MXN2 pm nmin net90 VPW n12 l=1.3e-07 w=5.1e-07
MXN3 pm c net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 net74 RN VSS VPW n12 l=1.3e-07 w=6.8e-07
MXN11 m pm net74 VPW n12 l=1.3e-07 w=6.8e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.4e-07
MXN7 bm cn net86 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net86 RN net83 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net83 VPW n12 l=1.3e-07 w=1.5e-07
mXI50_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI51_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net131 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP18 net131 c cn VNW p12 l=1.3e-07 w=4.5e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP19 pm nmin net105 VNW p12 l=1.3e-07 w=6.2e-07
MXP20 pm cn net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP5 VDD m net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=8.5e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.1e-07
mXI58_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=5.3e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=2.7e-07
MXP21 bm c net125 VNW p12 l=1.3e-07 w=1.5e-07
MXP15 VDD s net125 VNW p12 l=1.3e-07 w=1.5e-07
mXI50_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRHQX4MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MXN15 net90 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm nmin net90 VPW n12 l=1.3e-07 w=5.1e-07
MXN3 pm c net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net74 RN VSS VPW n12 l=1.3e-07 w=5.9e-07
MXN11 m pm net74 VPW n12 l=1.3e-07 w=5.9e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MXN7 bm cn net86 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net86 RN net83 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net83 VPW n12 l=1.3e-07 w=1.5e-07
mXI50_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net131 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP18 net131 c cn VNW p12 l=1.3e-07 w=4.5e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
MXP2 net105 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP19 pm nmin net105 VNW p12 l=1.3e-07 w=6.2e-07
MXP20 pm cn net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP5 VDD m net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP6_2 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI58_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=3e-07
MXP21 bm c net125 VNW p12 l=1.3e-07 w=1.5e-07
MXP15 VDD s net125 VNW p12 l=1.3e-07 w=1.5e-07
mXI50_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRHQX8MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MXN15 net90 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm nmin net90 VPW n12 l=1.3e-07 w=5.1e-07
MXN3 pm c net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net74 RN VSS VPW n12 l=1.3e-07 w=5.9e-07
MXN11 m pm net74 VPW n12 l=1.3e-07 w=5.9e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MXN7 bm cn net86 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net86 RN net83 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net83 VPW n12 l=1.3e-07 w=1.5e-07
mXI50_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net131 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP18 net131 c cn VNW p12 l=1.3e-07 w=4.5e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
MXP2 net105 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP19 pm nmin net105 VNW p12 l=1.3e-07 w=6.2e-07
MXP20 pm cn net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP5 VDD m net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP6_2 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI58_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=3e-07
MXP21 bm c net125 VNW p12 l=1.3e-07 w=1.5e-07
MXP15 VDD s net125 VNW p12 l=1.3e-07 w=1.5e-07
mXI50_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRQX1MTR Q VDD VNW VPW VSS CK D RN
MXN5 net86 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net78 D net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 pm cn net78 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 pm c net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net66 m net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net66 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI37_MXNOE net119 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE net119 cn XI4_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 s net119 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP4 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 D VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP6 pm c net105 VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI37_MXPOEN net119 cn m VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN net119 c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 s net119 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFRQX2MTR Q VDD VNW VPW VSS CK D RN
MXN5 net86 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net78 D net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 pm cn net78 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 pm c net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net66 m net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net66 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI37_MXNOE net119 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE net119 cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 s net119 XI0_n1 VPW n12 l=1.3e-07 w=2.7e-07
mXI0_MXNA2 XI0_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 D VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP6 pm c net105 VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3e-07
mXI37_MXPOEN net119 cn m VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN net119 c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 s net119 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRQX4MTR Q VDD VNW VPW VSS CK D RN
MXN5 net86 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net78 D net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 pm cn net78 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 pm c net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net66 m net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net66 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI37_MXNOE net119 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE net119 cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 s net119 XI0_n1 VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA2 XI0_n1 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 D VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP6 pm c net105 VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3e-07
mXI37_MXPOEN net119 cn m VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN net119 c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 s net119 VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRX1MTR Q QN VDD VNW VPW VSS CK D RN
MXN2 pm cn net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net45 D net53 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net53 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 pm c net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net61 m net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net61 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE bm cn XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 net90 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 net90 bm XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI45_MXNA1 Q net90 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP2 net68 D VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm c net68 VNW p12 l=1.3e-07 w=4.1e-07
MXP1 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MXP7 pm cn net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD m net72 VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI40_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI5_MXPOEN bm c XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 net90 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 net90 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 net90 bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI45_MXPA1 Q net90 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFRX2MTR Q QN VDD VNW VPW VSS CK D RN
MXN2 pm cn net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net45 D net53 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net53 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 pm c net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net61 m net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net61 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE bm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 net90 VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1 net90 bm XI1_n1 VPW n12 l=1.3e-07 w=2.7e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI45_MXNA1 Q net90 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP2 net68 D VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm c net68 VNW p12 l=1.3e-07 w=4.1e-07
MXP1 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 pm cn net72 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 VDD m net72 VNW p12 l=1.3e-07 w=2.2e-07
mXI43_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI40_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI5_MXPOEN bm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 net90 VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 net90 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 net90 bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI45_MXPA1 Q net90 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRX4MTR Q QN VDD VNW VPW VSS CK D RN
MXN2 pm cn net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net45 D net53 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net53 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 pm c net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net61 m net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net61 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE bm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 net90 VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1 net90 bm XI1_n1 VPW n12 l=1.3e-07 w=4.9e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI46_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI45_MXNA1 Q net90 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI45_MXNA1_2 Q net90 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP2 net68 D VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm c net68 VNW p12 l=1.3e-07 w=4.1e-07
MXP1 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 pm cn net72 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 VDD m net72 VNW p12 l=1.3e-07 w=2.2e-07
mXI43_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI40_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI5_MXPOEN bm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 net90 VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 net90 RN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 net90 bm VDD VNW p12 l=1.3e-07 w=3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI46_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI45_MXPA1 Q net90 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI45_MXPA1_2 Q net90 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSHQX1MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 VSS SN net92 VPW n12 l=1.3e-07 w=4.5e-07
MXN7 net92 cn net89 VPW n12 l=1.3e-07 w=4.5e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP7 net099 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 pm nmin net091 VNW p12 l=1.3e-07 w=3.7e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT DFFSHQX2MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS SN net92 VPW n12 l=1.3e-07 w=6.4e-07
MXN11 net92 cn net89 VPW n12 l=1.3e-07 w=6.4e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=6.4e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP13 net099 c cn VNW p12 l=1.3e-07 w=4.9e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmin net091 VNW p12 l=1.3e-07 w=5.4e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSHQX4MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN14 VSS SN net92 VPW n12 l=1.3e-07 w=7.5e-07
MXN13 net92 cn net89 VPW n12 l=1.3e-07 w=7.5e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=7.5e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP15 net099 c cn VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP16 pm nmin net091 VNW p12 l=1.3e-07 w=6.9e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSHQX8MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN14 VSS SN net92 VPW n12 l=1.3e-07 w=7.5e-07
MXN13 net92 cn net89 VPW n12 l=1.3e-07 w=7.5e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=7.5e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP15 net099 c cn VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP16 pm nmin net091 VNW p12 l=1.3e-07 w=6.9e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSQX1MTR Q VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN2 bm cn net84 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 NSN s net84 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI34_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm c net62 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD s net62 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSQX2MTR Q VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN2 bm cn net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 NSN s net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN1 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI34_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 bm c net53 VNW p12 l=1.3e-07 w=1.5e-07
MXP7 VDD s net53 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSQX4MTR Q VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN2 bm cn net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 NSN s net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN1 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI34_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 bm c net53 VNW p12 l=1.3e-07 w=1.5e-07
MXP7 VDD s net53 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRHQX1MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 VSS SN net62 VPW n12 l=1.3e-07 w=4.1e-07
MXN12 net62 cn net82 VPW n12 l=1.3e-07 w=4.1e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=4.1e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=4.3e-07
MXN14 VSS RN net70 VPW n12 l=1.3e-07 w=4.3e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net122 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 pm nmin net128 VNW p12 l=1.3e-07 w=3.1e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP17 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.6e-07
MXP23 bm nmset net112 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSRHQX2MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN21 VSS SN net62 VPW n12 l=1.3e-07 w=5.8e-07
MXN20 net62 cn net82 VPW n12 l=1.3e-07 w=5.8e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=5.8e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=6.1e-07
MXN22 VSS RN net70 VPW n12 l=1.3e-07 w=6.1e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net122 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP25 pm nmin net128 VNW p12 l=1.3e-07 w=4.5e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP17 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP27 bm nmset net112 VNW p12 l=1.3e-07 w=2.7e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRHQX4MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS SN net62 VPW n12 l=1.3e-07 w=7.5e-07
MXN23 net62 cn net82 VPW n12 l=1.3e-07 w=7.5e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=7.5e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN25 VSS RN net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP28 net122 c cn VNW p12 l=1.3e-07 w=6.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.03e-06
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP29 pm nmin net128 VNW p12 l=1.3e-07 w=6.8e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP30 m RN net144 VNW p12 l=1.3e-07 w=3.1e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP31 bm nmset net112 VNW p12 l=1.3e-07 w=3.6e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRHQX8MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS SN net62 VPW n12 l=1.3e-07 w=7.5e-07
MXN23 net62 cn net82 VPW n12 l=1.3e-07 w=7.5e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=7.5e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN25 VSS RN net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP28 net122 c cn VNW p12 l=1.3e-07 w=6.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.03e-06
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP29 pm nmin net128 VNW p12 l=1.3e-07 w=6.8e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP30 m RN net144 VNW p12 l=1.3e-07 w=3.1e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP31 bm nmset net112 VNW p12 l=1.3e-07 w=3.6e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRX1MTR Q QN VDD VNW VPW VSS CK D RN SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm c XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MXN2 m NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MXN3 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MXN8 bm cn net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 NSN s net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm cn XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net_NRN NRN VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP6 m pm net_NRN VNW p12 l=1.3e-07 w=3.6e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MXP7 bm c net75 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net_NRN s net75 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSRX2MTR Q QN VDD VNW VPW VSS CK D RN SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm c XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MXN2 m NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MXN3 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MXN4 bm cn net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 NSN s net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm cn XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net_NRN NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 m pm net_NRN VNW p12 l=1.3e-07 w=4.4e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.4e-07
MXP7 bm c net75 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net_NRN s net75 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRX4MTR Q QN VDD VNW VPW VSS CK D RN SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI4_MXNOE pm c XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MXN2 m NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=4.7e-07
MXN3 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MXN4 bm cn net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 NSN s net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN SN VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm cn XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net_NRN NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 m pm net_NRN VNW p12 l=1.3e-07 w=4.4e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.7e-07
MXP7 bm c net75 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net_NRN s net75 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSX1MTR Q QN VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm BSN VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MXN1 bm cn net134 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 BSN s net134 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 BSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net73 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSX2MTR Q QN VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN0 m pm BSN VPW n12 l=1.3e-07 w=2.1e-07
MXN0_2 m pm BSN VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MXN1 bm cn net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN4 BSN s net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.1e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm c net73 VNW p12 l=1.3e-07 w=1.5e-07
MXP6 VDD s net73 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSX4MTR Q QN VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=2e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=2e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 m pm BSN VPW n12 l=1.3e-07 w=3.3e-07
MXN0_2 m pm BSN VPW n12 l=1.3e-07 w=3.3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=5.2e-07
MXN1 bm cn net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN4 BSN s net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN SN VSS VPW n12 l=1.3e-07 w=1.08e-06
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=5.6e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.4e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.2e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm c net73 VNW p12 l=1.3e-07 w=1.5e-07
MXP6 VDD s net73 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFTRX1MTR Q QN VDD VNW VPW VSS CK D RN
MXN4 net129 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net132 D net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm cn net132 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
mXI4_MXNOE bm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g11_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP4 net62 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm c net62 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI4_MXPOEN bm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g11_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFTRX2MTR Q QN VDD VNW VPW VSS CK D RN
MXN6 net129 RN VSS VPW n12 l=1.3e-07 w=2.6e-07
MXN5 net132 D net129 VPW n12 l=1.3e-07 w=2.6e-07
MXN1 pm cn net132 VPW n12 l=1.3e-07 w=2.6e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI4_MXNOE bm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g11_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 net62 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP5 pm c net62 VNW p12 l=1.3e-07 w=2.6e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.7e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI4_MXPOEN bm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g11_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFTRX4MTR Q QN VDD VNW VPW VSS CK D RN
MXN8 net129 RN VSS VPW n12 l=1.3e-07 w=5e-07
MXN7 net132 D net129 VPW n12 l=1.3e-07 w=5e-07
MXN1 pm cn net132 VPW n12 l=1.3e-07 w=5e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=4e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=8e-07
mXI4_MXNOE bm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g11_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g11_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 net62 RN VDD VNW p12 l=1.3e-07 w=2.5e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP6 pm c net62 VNW p12 l=1.3e-07 w=5.1e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.6e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_3 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_4 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI47_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI4_MXPOEN bm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g11_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g11_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFX1MTR Q QN VDD VNW VPW VSS CK D
mXI14_MXNA1 XI14_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNOE pm cn XI14_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI12_MXNOE nm c XI12_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI11_MXNOE nm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI14_MXPA1 XI14_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI14_MXPOEN pm c XI14_p1 VNW p12 l=1.3e-07 w=3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI12_MXPOEN nm cn XI12_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI11_MXPOEN nm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFX2MTR Q QN VDD VNW VPW VSS CK D
mXI14_MXNA1 XI14_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNOE pm cn XI14_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=4e-07
mXI12_MXNOE nm c XI12_n1 VPW n12 l=1.3e-07 w=4e-07
mXI11_MXNOE nm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1 XI14_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI14_MXPOEN pm c XI14_p1 VNW p12 l=1.3e-07 w=3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=4.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI12_MXPOEN nm cn XI12_p1 VNW p12 l=1.3e-07 w=4.9e-07
mXI11_MXPOEN nm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFX4MTR Q QN VDD VNW VPW VSS CK D
mXI14_MXNA1 XI14_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNOE pm cn XI14_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=5.8e-07
mXI12_MXNOE nm c XI12_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI11_MXNOE nm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1 XI14_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI14_MXPOEN pm c XI14_p1 VNW p12 l=1.3e-07 w=3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g14_MXPA1_2 cn CK VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.7e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI12_MXPOEN nm cn XI12_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI11_MXPOEN nm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends



.SUBCKT EDFFHQX1MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 VSS s net104 VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=3.6e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=4e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=3e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 nmsi E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=4.5e-07
MXP0 cn c net053 VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP2 pm nmsi net047 VNW p12 l=1.3e-07 w=4.4e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=7.9e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT EDFFHQX2MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 VSS s net104 VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=5.1e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.2e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.6e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=3.9e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 nmsi E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=4.5e-07
MXP0 cn c net053 VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=8e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 pm nmsi net047 VNW p12 l=1.3e-07 w=6.2e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFHQX4MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=2.3e-07
MXN3 VSS s net104 VPW n12 l=1.3e-07 w=2.3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=5.1e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmsi E net73 VNW p12 l=1.3e-07 w=2.8e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=5e-07
MXP4 cn c net053 VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 pm nmsi net047 VNW p12 l=1.3e-07 w=6.2e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFHQX8MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=2.3e-07
MXN3 VSS s net104 VPW n12 l=1.3e-07 w=2.3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=5.1e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmsi E net73 VNW p12 l=1.3e-07 w=2.8e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=5e-07
MXP4 cn c net053 VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 pm nmsi net047 VNW p12 l=1.3e-07 w=6.2e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFTRX1MTR Q QN VDD VNW VPW VSS CK D E RN
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net122 s net140 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net122 nmen net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net107 E net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net140 D net107 VPW n12 l=1.3e-07 w=1.8e-07
MX_t3 net106 RN VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t19 pm cn net140 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI11_MXNOE bnm c XI11_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI5_MXNOE bnm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bnm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 net77 s net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 VDD nmen net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net76 D net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 VDD RN net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net77 c pm VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI11_MXPA1 XI11_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI11_MXPOEN bnm cn XI11_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI5_MXPOEN bnm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bnm VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT EDFFTRX2MTR Q QN VDD VNW VPW VSS CK D E RN
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net122 s net140 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net122 nmen net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net107 E net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net140 D net107 VPW n12 l=1.3e-07 w=1.8e-07
MX_t3 net106 RN VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t19 pm cn net140 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 m VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI11_MXNOE bnm c XI11_n1 VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE bnm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g1_MXNA1 Q bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 net77 s net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 VDD nmen net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net76 D net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 VDD RN net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net77 c pm VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI11_MXPA1 XI11_p1 m VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI11_MXPOEN bnm cn XI11_p1 VNW p12 l=1.3e-07 w=5.2e-07
mXI5_MXPOEN bnm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g1_MXPA1 Q bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFTRX4MTR Q QN VDD VNW VPW VSS CK D E RN
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net122 s net140 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net122 nmen net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net107 E net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net140 D net107 VPW n12 l=1.3e-07 w=1.8e-07
MX_t3 net106 RN VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t19 pm cn net140 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 m VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI11_MXNOE bnm c XI11_n1 VPW n12 l=1.3e-07 w=6.3e-07
mXI5_MXNOE bnm cn XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g1_MXNA1 Q bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 net77 s net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 VDD nmen net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net76 D net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 VDD RN net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net77 c pm VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI11_MXPA1 XI11_p1 m VDD VNW p12 l=1.3e-07 w=8.2e-07
mXI11_MXPOEN bnm cn XI11_p1 VNW p12 l=1.3e-07 w=8.2e-07
mXI5_MXPOEN bnm c XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g1_MXPA1 Q bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFX1MTR Q QN VDD VNW VPW VSS CK D E
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net120 s net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net120 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net123 E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net129 D net123 VPW n12 l=1.3e-07 w=1.8e-07
MX_t19 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI1_MXNOE nm c XI1_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net38 s net36 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 VDD E net36 VNW p12 l=1.3e-07 w=3.8e-07
MX_t5 VDD nmen net39 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net39 D net38 VNW p12 l=1.3e-07 w=3.8e-07
MXP2 net38 c pm VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI1_MXPOEN nm cn XI1_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT EDFFX2MTR Q QN VDD VNW VPW VSS CK D E
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net120 s net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net120 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net123 E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net129 D net123 VPW n12 l=1.3e-07 w=1.8e-07
MX_t19 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI1_MXNOE nm c XI1_n1 VPW n12 l=1.3e-07 w=4.3e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net38 s net36 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 VDD E net36 VNW p12 l=1.3e-07 w=3.8e-07
MX_t5 VDD nmen net39 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net39 D net38 VNW p12 l=1.3e-07 w=3.8e-07
MXP2 net38 c pm VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI1_MXPOEN nm cn XI1_p1 VNW p12 l=1.3e-07 w=5.2e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFX4MTR Q QN VDD VNW VPW VSS CK D E
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net120 s net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net120 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net123 E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net129 D net123 VPW n12 l=1.3e-07 w=1.8e-07
MX_t19 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI1_MXNOE nm c XI1_n1 VPW n12 l=1.3e-07 w=6.4e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net38 s net36 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 VDD E net36 VNW p12 l=1.3e-07 w=3.8e-07
MX_t5 VDD nmen net39 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net39 D net38 VNW p12 l=1.3e-07 w=3.8e-07
MXP2 net38 c pm VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.7e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI1_MXPOEN nm cn XI1_p1 VNW p12 l=1.3e-07 w=7.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=5e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MDFFHQX1MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=2.1e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 net135 cn VSS VPW n12 l=1.3e-07 w=3.3e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=3.3e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=3.7e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t9 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=2.6e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=3e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=3e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=4.2e-07
MXP0 cn c net50 VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=4e-07
MXP1 pm nmsi net61 VNW p12 l=1.3e-07 w=4e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=7.3e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MDFFHQX2MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=3.1e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=3e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN1 net135 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=4.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=4.4e-07
MXP2 cn c net50 VNW p12 l=1.3e-07 w=4.4e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=7.6e-07
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP5 pm nmsi net61 VNW p12 l=1.3e-07 w=5.9e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=9.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=9.8e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MDFFHQX4MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=5e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN2 net135 cn VSS VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=5.6e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net50 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net61 VNW p12 l=1.3e-07 w=1.01e-06
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MDFFHQX8MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=4.9e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN2 net135 cn VSS VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=5.6e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.3e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net50 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net61 VNW p12 l=1.3e-07 w=1.01e-06
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends

***********************************************************

.SUBCKT SDFFHQNX1MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net71 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net48 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 pm nmsi net60 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFHQNX2MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net71 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net48 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.6e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 pm nmsi net60 VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT SDFFHQNX4MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=2.9e-07
MXN2 net71 cn VSS VPW n12 l=1.3e-07 w=2.9e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.2e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=5e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net48 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP3 pm nmsi net60 VNW p12 l=1.3e-07 w=3.5e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=6.1e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFHQNX8MTR QN VDD VNW VPW VSS CK D SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=3.4e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3e-07
MXN3 net71 cn VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 pm nmsi net71 VPW n12 l=1.3e-07 w=5.4e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNOE bm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g2_MXNA1_2 s bm VSS VPW n12 l=1.3e-07 w=4.8e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=4.2e-07
MX_t10 net48 CK VDD VNW p12 l=1.3e-07 w=4.8e-07
MXP4 net48 c cn VNW p12 l=1.3e-07 w=4.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.3e-07
MX_t8 net60 c VDD VNW p12 l=1.3e-07 w=6.5e-07
MXP5 pm nmsi net60 VNW p12 l=1.3e-07 w=6.5e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.5e-07
mXI7_MXPOEN bm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=6e-07
mX_g2_MXPA1_2 s bm VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFHQX1MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.1e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=3.3e-07
MXN1 net54 cn VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.7e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP0 net065 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.6e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=4e-07
MXP2 pm nmsi net71 VNW p12 l=1.3e-07 w=4e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.3e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
.ends


.SUBCKT SDFFHQX2MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=1.9e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=3.1e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=4.8e-07
MXN2 net54 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP3 net065 c cn VNW p12 l=1.3e-07 w=4.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP4 pm nmsi net71 VNW p12 l=1.3e-07 w=5.9e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
.ends


.SUBCKT SDFFHQX4MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=3.2e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.5e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.4e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=6.9e-07
MXN3 net54 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP5 net065 c cn VNW p12 l=1.3e-07 w=7.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=6.7e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP6 pm nmsi net71 VNW p12 l=1.3e-07 w=8e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT SDFFHQX8MTR Q VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 VSS CK cn VPW n12 l=1.3e-07 w=5.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.5e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.4e-07
MX_t3 pm nmsi net54 VPW n12 l=1.3e-07 w=6.9e-07
MXN3 net54 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.9e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP1 net065 CK VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP5 net065 c cn VNW p12 l=1.3e-07 w=7.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=6.7e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=5e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=8.3e-07
MX_t8 net71 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP6 pm nmsi net71 VNW p12 l=1.3e-07 w=8e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT SDFFHX1MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.3e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net0107 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 net104 cn VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 net079 c cn VNW p12 l=1.3e-07 w=4.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.8e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.8e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 nmsi SI net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP10 pm nmsi net087 VNW p12 l=1.3e-07 w=4.4e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.9e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFHX2MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=3.2e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net0107 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=5.1e-07
MXN7 net104 cn VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP13 net079 c cn VNW p12 l=1.3e-07 w=4.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.9e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 nmsi SI net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP12 pm nmsi net087 VNW p12 l=1.3e-07 w=6.2e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g6_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.1e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT SDFFHX4MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.4e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=2.9e-07
MXN8 net0107 SE VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=7e-07
MXN9 net104 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 net079 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=7e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP14 nmsi SI net76 VNW p12 l=1.3e-07 w=3.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 pm nmsi net087 VNW p12 l=1.3e-07 w=8.7e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g6_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT SDFFHX8MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI62_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.4e-07
MX_t20 nmsi SI net0107 VPW n12 l=1.3e-07 w=2.9e-07
MXN8 net0107 SE VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t3 pm nmsi net104 VPW n12 l=1.3e-07 w=7e-07
MXN9 net104 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI60_MXNOE pm c XI60_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI60_MXNA1 XI60_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI14_MXNOE bm cn XI14_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI14_MXNA1 XI14_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP13 net079 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI62_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=7e-07
MX_t22 net76 nmse VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP14 nmsi SI net76 VNW p12 l=1.3e-07 w=3.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t8 net087 c VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 pm nmsi net087 VNW p12 l=1.3e-07 w=8.7e-07
mXI60_MXPOEN pm cn XI60_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPA1 XI60_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g6_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI14_MXPOEN bm c XI14_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI14_MXPA1 XI14_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT SDFFNHX1MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmsi SI n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 n1 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=4.3e-07
MXN5 net58 cn VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=4e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP2 net87 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP8 p1 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmsi SI p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=6.8e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP10 pm nmsi net93 VNW p12 l=1.3e-07 w=3.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=4.8e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFNHX2MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmsi SI n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 n1 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=6.1e-07
MXN1 net58 cn VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP2 net87 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP8 p1 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmsi SI p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=8.4e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP5 pm nmsi net93 VNW p12 l=1.3e-07 w=4.6e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFNHX4MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.7e-07
MXN5 nmsi SI net058 VPW n12 l=1.3e-07 w=2.7e-07
MXN7 net058 SE VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=4.6e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=5.4e-07
MXN1 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MX_t3_2 pm nmsi net58 VPW n12 l=1.3e-07 w=5.4e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI59_MXNOE_2 nm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP10 net87 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.3e-07
MXP14 p1 nmse VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP9 nmsi SI p1 VNW p12 l=1.3e-07 w=3.3e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g10_MXPA1_2 cn net185 VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP13 pm nmsi net93 VNW p12 l=1.3e-07 w=6.9e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN_2 nm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g1_MXPA1_3 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT SDFFNHX8MTR Q QN VDD VNW VPW VSS CKN D SE SI
mX_g14_MXNA1 net185 CKN VSS VPW n12 l=1.3e-07 w=4.7e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.1e-07
MXN7 nmsi SI n1 VPW n12 l=1.3e-07 w=5.1e-07
MXN6 n1 SE VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g10_MXNA1 cn net185 VSS VPW n12 l=1.3e-07 w=5e-07
MX_t3 pm nmsi net58 VPW n12 l=1.3e-07 w=7.4e-07
MXN1 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 net58 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MX_t3_2 pm nmsi net58 VPW n12 l=1.3e-07 w=7.4e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI59_MXNOE nm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI59_MXNOE_2 nm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE nm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net185 CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MX_t10 net87 CKN VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP14 net87 cn c VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.5e-07
MXP8 p1 nmse VDD VNW p12 l=1.3e-07 w=3.4e-07
MXP15 nmsi SI p1 VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 cn net185 VDD VNW p12 l=1.3e-07 w=7.2e-07
mX_g10_MXPA1_2 cn net185 VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP0 net93 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP13 pm nmsi net93 VNW p12 l=1.3e-07 w=6.9e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.7e-07
mXI59_MXPOEN nm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN_2 nm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI8_MXPOEN nm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFNSRHX1MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net0207 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net0207 VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MX_t30 nmsi SI net172 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 net172 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS SN net163 VPW n12 l=1.3e-07 w=4.3e-07
MXN17 net163 cn net160 VPW n12 l=1.3e-07 w=4.3e-07
MX_t26 pm nmsi net160 VPW n12 l=1.3e-07 w=4.3e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 net0106 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t12 net0106 pm net166 VPW n12 l=1.3e-07 w=4.5e-07
MXN19 VSS RN net166 VPW n12 l=1.3e-07 w=4.5e-07
MXN20 net0106 nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE bm c net0106 VPW n12 l=1.3e-07 w=4e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net181 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net181 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 net0207 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net080 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net080 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn net0207 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP16 nmsi SI net117 VNW p12 l=1.3e-07 w=2.3e-07
MX_t32 net117 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP17 pm nmsi net0125 VNW p12 l=1.3e-07 w=3.3e-07
MX_t24 net0125 c VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI23_MXPA1 XI23_p1 net0106 VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 net0106 pm VDD VNW p12 l=1.3e-07 w=4.8e-07
MXP18 net111 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net0106 RN net111 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net0106 VNW p12 l=1.3e-07 w=4.8e-07
MXP21 bm nmset net126 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 net126 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP24 bm c net132 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net132 nmset net135 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net135 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT SDFFNSRHX2MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net261 CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net261 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=1.8e-07
MX_t30 nmsi SI net168 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 net168 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN26 VSS SN net149 VPW n12 l=1.3e-07 w=6.1e-07
MXN25 net149 cn net153 VPW n12 l=1.3e-07 w=6.1e-07
MX_t26 pm nmsi net153 VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 net129 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN27 net129 pm net145 VPW n12 l=1.3e-07 w=6.3e-07
MXN28 VSS RN net145 VPW n12 l=1.3e-07 w=6.3e-07
MXN20 net129 nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE bm c net129 VPW n12 l=1.3e-07 w=5.5e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net261 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net109 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net109 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn net261 VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=2.3e-07
MXP16 nmsi SI net91 VNW p12 l=1.3e-07 w=2.3e-07
MX_t32 net91 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP25 pm nmsi net83 VNW p12 l=1.3e-07 w=4.6e-07
MX_t24 net83 c VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI23_MXPA1 XI23_p1 net129 VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 net129 pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP18 net103 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net129 RN net103 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net129 VNW p12 l=1.3e-07 w=6.7e-07
MXP28 bm nmset net79 VNW p12 l=1.3e-07 w=2.8e-07
MXP20 net79 RN VDD VNW p12 l=1.3e-07 w=2.8e-07
MXP24 bm c net123 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net123 nmset net119 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net119 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFNSRHX4MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net261 CKN VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net261 VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=2.7e-07
MX_t30 nmsi SI net168 VPW n12 l=1.3e-07 w=2.7e-07
MXN29 net168 SE VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN31 VSS SN net149 VPW n12 l=1.3e-07 w=7.6e-07
MXN30 net149 cn net153 VPW n12 l=1.3e-07 w=7.6e-07
MX_t26 pm nmsi net153 VPW n12 l=1.3e-07 w=7.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 net129 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN27 net129 pm net145 VPW n12 l=1.3e-07 w=8.4e-07
MXN32 VSS RN net145 VPW n12 l=1.3e-07 w=8.4e-07
MXN20 net129 nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI74_MXNOE bm c net129 VPW n12 l=1.3e-07 w=5.5e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net261 CKN VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net109 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP29 net109 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 cn net261 VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=3.2e-07
MXP30 nmsi SI net91 VNW p12 l=1.3e-07 w=3.3e-07
MX_t32 net91 nmse VDD VNW p12 l=1.3e-07 w=3.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP31 pm nmsi net83 VNW p12 l=1.3e-07 w=6.9e-07
MX_t24 net83 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI23_MXPA1 XI23_p1 net129 VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t10_2 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP18 net103 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net129 RN net103 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net129 VNW p12 l=1.3e-07 w=6.7e-07
MXP32 bm nmset net79 VNW p12 l=1.3e-07 w=3.6e-07
MXP20 net79 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP24 bm c net123 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net123 nmset net119 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net119 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFNSRHX8MTR Q QN VDD VNW VPW VSS CKN D RN SE SI SN
mX_g14_MXNA1 net261 CKN VSS VPW n12 l=1.3e-07 w=4.7e-07
MX_t6 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn net261 VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g10_MXNA1_2 cn net261 VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI65_MXNOE nmsi nmse nmin VPW n12 l=1.3e-07 w=5.4e-07
MX_t30 nmsi SI net168 VPW n12 l=1.3e-07 w=5.1e-07
MXN33 net168 SE VSS VPW n12 l=1.3e-07 w=5.1e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN31 VSS SN net149 VPW n12 l=1.3e-07 w=7.6e-07
MXN30 net149 cn net153 VPW n12 l=1.3e-07 w=7.6e-07
MX_t26 pm nmsi net153 VPW n12 l=1.3e-07 w=7.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI23_MXNA1 XI23_n1 net129 VSS VPW n12 l=1.3e-07 w=2.5e-07
MXN27 net129 pm net145 VPW n12 l=1.3e-07 w=8.7e-07
MXN34 VSS RN net145 VPW n12 l=1.3e-07 w=8.7e-07
MXN20 net129 nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI74_MXNOE bm c net129 VPW n12 l=1.3e-07 w=5.5e-07
MXN22 bm cn net184 VPW n12 l=1.3e-07 w=1.8e-07
MXN23 net184 RN net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS s net161 VPW n12 l=1.3e-07 w=1.8e-07
MXN21 bm nmset VSS VPW n12 l=1.3e-07 w=3e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 net261 CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MX_t4 net109 CKN VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP33 net109 cn c VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 cn net261 VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g10_MXPA1_2 cn net261 VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=1.03e-06
mXI65_MXPOEN nmsi SE nmin VNW p12 l=1.3e-07 w=5.8e-07
MXP34 nmsi SI net91 VNW p12 l=1.3e-07 w=5.6e-07
MX_t32 net91 nmse VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=3.3e-07
MX_t11 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP31 pm nmsi net83 VNW p12 l=1.3e-07 w=6.9e-07
MX_t24 net83 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI23_MXPA1 XI23_p1 net129 VDD VNW p12 l=1.3e-07 w=3.1e-07
MX_t10 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t10_2 net129 pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP18 net103 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net129 RN net103 VNW p12 l=1.3e-07 w=2.3e-07
mXI74_MXPOEN bm cn net129 VNW p12 l=1.3e-07 w=6.7e-07
MXP35 bm nmset net79 VNW p12 l=1.3e-07 w=3.5e-07
MXP20 net79 RN VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP24 bm c net123 VNW p12 l=1.3e-07 w=2.3e-07
MXP23 net123 nmset net119 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 VDD s net119 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQNX1MTR QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net108 SE net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 VSS SI net108 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net111 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net129 D net111 VPW n12 l=1.3e-07 w=1.8e-07
MX_t1 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE pm c XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.7e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net69 nmse net65 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net65 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net68 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net69 D net68 VNW p12 l=1.3e-07 w=3.8e-07
MXP5 pm c net69 VNW p12 l=1.3e-07 w=3.8e-07
mXI1_MXPOEN pm cn XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFQNX2MTR QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net108 SE net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 VSS SI net108 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net111 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net129 D net111 VPW n12 l=1.3e-07 w=1.8e-07
MX_t1 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE pm c XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.7e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP6 net69 nmse net65 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net65 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net68 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net69 D net68 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 pm c net69 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN pm cn XI1_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQNX4MTR QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net108 SE net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 VSS SI net108 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net111 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net129 D net111 VPW n12 l=1.3e-07 w=1.8e-07
MX_t1 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE pm c XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.7e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP6 net69 nmse net65 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net65 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net68 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net69 D net68 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 pm c net69 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN pm cn XI1_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQX1MTR Q VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net064 SE net055 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 VSS SI net064 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net059 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net055 D net059 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm cn net055 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE pm c XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net105 m VSS VPW n12 l=1.3e-07 w=2.8e-07
MX_t12 ns c net105 VPW n12 l=1.3e-07 w=2.8e-07
mXI15_MXNOE ns cn XI15_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI15_MXNA1 XI15_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net076 nmse net070 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net070 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net074 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net076 D net074 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 pm c net076 VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN pm cn XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MX_t14 net80 m VDD VNW p12 l=1.3e-07 w=3.4e-07
MXP7 ns cn net80 VNW p12 l=1.3e-07 w=3.4e-07
mXI15_MXPOEN ns c XI15_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI15_MXPA1 XI15_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFQX2MTR Q VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net064 SE net055 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 VSS SI net064 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net059 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net055 D net059 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm cn net055 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE pm c XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net105 m VSS VPW n12 l=1.3e-07 w=3.9e-07
MX_t12 ns c net105 VPW n12 l=1.3e-07 w=3.9e-07
mXI15_MXNOE ns cn XI15_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI15_MXNA1 XI15_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net076 nmse net070 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net070 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net074 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net076 D net074 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 pm c net076 VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN pm cn XI16_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI16_MXPA1 XI16_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=4.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MX_t14 net80 m VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP8 ns cn net80 VNW p12 l=1.3e-07 w=4.9e-07
mXI15_MXPOEN ns c XI15_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI15_MXPA1 XI15_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFQX4MTR Q VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net064 SE net055 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 VSS SI net064 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net059 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net055 D net059 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm cn net055 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE pm c XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net105 m VSS VPW n12 l=1.3e-07 w=4.4e-07
MX_t12 ns c net105 VPW n12 l=1.3e-07 w=4.4e-07
mXI15_MXNOE ns cn XI15_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI15_MXNA1 XI15_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net076 nmse net070 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net070 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net074 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net076 D net074 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 pm c net076 VNW p12 l=1.3e-07 w=3.8e-07
mXI16_MXPOEN pm cn XI16_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI16_MXPA1 XI16_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MX_t14 net80 m VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP9 ns cn net80 VNW p12 l=1.3e-07 w=6.4e-07
mXI15_MXPOEN ns c XI15_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI15_MXPA1 XI15_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRHQX1MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=3.5e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=3.5e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS RN net128 VPW n12 l=1.3e-07 w=4.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=4.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.7e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP8 net065 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=2.7e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP13 pm nmsi p1 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=6.6e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.3e-07
MX_t15 bm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 bm c net109 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=2.3e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFRHQX2MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS RN net128 VPW n12 l=1.3e-07 w=5.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=5.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP14 net065 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.9e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 pm nmsi p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
MX_t10_2 m pm VDD VNW p12 l=1.3e-07 w=5.1e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 bm RN VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP16 bm c net109 VNW p12 l=1.3e-07 w=1.5e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=1.5e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRHQX4MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS RN net128 VPW n12 l=1.3e-07 w=5.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=5.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP14 net065 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.9e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 pm nmsi p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
MX_t10_2 m pm VDD VNW p12 l=1.3e-07 w=5.1e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 bm RN VDD VNW p12 l=1.3e-07 w=3e-07
MXP16 bm c net109 VNW p12 l=1.3e-07 w=1.5e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=1.5e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRHQX8MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mXI69_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 n1 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 pm nmsi n1 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS RN net128 VPW n12 l=1.3e-07 w=5.9e-07
MX_t11 m pm net128 VPW n12 l=1.3e-07 w=5.9e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MX_t18 bm cn net149 VPW n12 l=1.3e-07 w=1.5e-07
MXN7 net149 RN net146 VPW n12 l=1.3e-07 w=1.5e-07
MXN8 VSS s net146 VPW n12 l=1.3e-07 w=1.5e-07
mXI26_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t4 net065 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP14 net065 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
mXI69_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.9e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 p1 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 pm nmsi p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
MX_t10_2 m pm VDD VNW p12 l=1.3e-07 w=5.1e-07
MX_t7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 bm RN VDD VNW p12 l=1.3e-07 w=3e-07
MXP16 bm c net109 VNW p12 l=1.3e-07 w=1.5e-07
MXP9 VDD s net109 VNW p12 l=1.3e-07 w=1.5e-07
mXI26_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRQX1MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net130 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net130 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net138 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MX_t9 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN7 pm c net123 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net118 m net123 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net118 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE net76 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE net76 cn XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 s net76 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net97 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 nmrs SE net97 VNW p12 l=1.3e-07 w=3e-07
MXP1 nmrs nmse net105 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net105 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI74_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN net76 cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN net76 c XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s net76 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFRQX2MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net130 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net130 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net138 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MX_t9 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm c net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 net118 m net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN6 net118 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE net76 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE net76 cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1 s net76 XI1_n1 VPW n12 l=1.3e-07 w=2.7e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net97 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 nmrs SE net97 VNW p12 l=1.3e-07 w=3e-07
MXP1 nmrs nmse net105 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net105 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI74_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm cn net89 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD m net89 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN net76 cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN net76 c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s net76 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRQX4MTR Q VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net130 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net130 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net138 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MX_t9 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI74_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm c net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 net118 m net123 VPW n12 l=1.3e-07 w=1.5e-07
MXN6 net118 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE net76 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE net76 cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1 s net76 XI1_n1 VPW n12 l=1.3e-07 w=4.9e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net97 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 nmrs SE net97 VNW p12 l=1.3e-07 w=3e-07
MXP1 nmrs nmse net105 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net105 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI74_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm cn net89 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD m net89 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI59_MXPOEN net76 cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN net76 c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 s net76 VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRX1MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net104 D net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MXN9 nmrs nmse net104 VPW n12 l=1.3e-07 w=2.4e-07
MXN7 nmrs SE net77 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net77 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
MXN12 pm c net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN13 net83 m net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net83 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNOE bm cn XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 s bm XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net139 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP10 nmrs SE net139 VNW p12 l=1.3e-07 w=3e-07
MXP8 nmrs nmse net115 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net115 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm cn net124 VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD m net124 VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPOEN bm c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFRX2MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net104 D net_clr_ VPW n12 l=1.3e-07 w=2.5e-07
MXN9 nmrs nmse net104 VPW n12 l=1.3e-07 w=2.5e-07
MXN7 nmrs SE net77 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net77 SI net_clr_ VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net_clr_ RN VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.9e-07
MXN12 pm c net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN16 net83 m net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN17 net83 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4.2e-07
mXI0_MXNOE bm cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1 s bm XI1_n1 VPW n12 l=1.3e-07 w=2.7e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net139 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP10 nmrs SE net139 VNW p12 l=1.3e-07 w=3e-07
MXP8 nmrs nmse net115 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net115 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
MXP13 pm cn net124 VNW p12 l=1.3e-07 w=1.5e-07
MXP12 VDD m net124 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.4e-07
mXI0_MXPOEN bm c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFRX4MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net104 D net_clr_ VPW n12 l=1.3e-07 w=4.9e-07
MXN9 nmrs nmse net104 VPW n12 l=1.3e-07 w=4.9e-07
MXN7 nmrs SE net77 VPW n12 l=1.3e-07 w=2.4e-07
MXN16 net77 SI net_clr_ VPW n12 l=1.3e-07 w=2.4e-07
MXN11 net_clr_ RN VSS VPW n12 l=1.3e-07 w=6.5e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=3.7e-07
MXN12 pm c net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN18 net83 m net89 VPW n12 l=1.3e-07 w=1.5e-07
MXN19 net83 RN VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g6_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=6.4e-07
mXI0_MXNOE bm cn XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1 s bm XI1_n1 VPW n12 l=1.3e-07 w=4.4e-07
mXI70_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI70_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net139 D VDD VNW p12 l=1.3e-07 w=6e-07
MXP14 nmrs SE net139 VNW p12 l=1.3e-07 w=6e-07
MXP13 nmrs nmse net115 VNW p12 l=1.3e-07 w=2.9e-07
MXP7 net115 SI VDD VNW p12 l=1.3e-07 w=2.9e-07
MXP3 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=3.9e-07
MXP15 pm cn net124 VNW p12 l=1.3e-07 w=1.5e-07
MXP12 VDD m net124 VNW p12 l=1.3e-07 w=1.5e-07
mX_g6_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.4e-07
mXI0_MXPOEN bm c XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mXI70_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI70_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSHQX1MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net0112 SN VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN3 net169 cn net0112 VPW n12 l=1.3e-07 w=4.5e-07
MX_t11 pm nmsi net169 VPW n12 l=1.3e-07 w=4.5e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP3 net088 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=3e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm nmsi net56 VNW p12 l=1.3e-07 w=3.7e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT SDFFSHQX2MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=3.4e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net0104 SN VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN8 net169 cn net0104 VPW n12 l=1.3e-07 w=6.5e-07
MX_t11 pm nmsi net169 VPW n12 l=1.3e-07 w=6.5e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP8 net088 c cn VNW p12 l=1.3e-07 w=4.9e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=4.2e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=4.2e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=2.3e-07
MXP9 pm nmsi net56 VNW p12 l=1.3e-07 w=5.4e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.01e-06
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSHQX4MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net0104 SN VSS VPW n12 l=1.3e-07 w=7.4e-07
MXN10 net169 cn net0104 VPW n12 l=1.3e-07 w=7.4e-07
MX_t11 pm nmsi net169 VPW n12 l=1.3e-07 w=7.4e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.9e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP10 net088 c cn VNW p12 l=1.3e-07 w=5.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=3.8e-07
MXP11 pm nmsi net56 VNW p12 l=1.3e-07 w=6.9e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSHQX8MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI73_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net0104 SN VSS VPW n12 l=1.3e-07 w=7.5e-07
MXN12 net169 cn net0104 VPW n12 l=1.3e-07 w=7.5e-07
MXN13 pm nmsi net169 VPW n12 l=1.3e-07 w=7.5e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN5 bm cn net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 VSS s net160 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 bm nmset_ VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g3_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.9e-07
MX_t4 net088 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP10 net088 c cn VNW p12 l=1.3e-07 w=5.2e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI73_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 VDD SN pm VNW p12 l=1.3e-07 w=3.8e-07
MXP11 pm nmsi net56 VNW p12 l=1.3e-07 w=6.9e-07
MX_t8 net56 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP7 net72 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net75 nmset_ net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net75 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSQX1MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmrs SE net150 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net150 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net123 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 nmrs nmse net123 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN11 bm cn net141 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 NSN s net141 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 nmrs SE net83 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net83 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 VDD SI net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net113 nmse nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 VDD pm m VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD SN m VNW p12 l=1.3e-07 w=2.3e-07
MXP13 VDD SN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP14 net107 c bm VNW p12 l=1.3e-07 w=2.3e-07
MXP15 net107 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSQX2MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmrs SE net150 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net150 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net123 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 nmrs nmse net123 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN11 bm cn net141 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 NSN s net141 VPW n12 l=1.3e-07 w=1.5e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 nmrs SE net83 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net83 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 VDD SI net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net113 nmse nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 VDD pm m VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD SN m VNW p12 l=1.3e-07 w=2.3e-07
MXP13 VDD SN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP16 net107 c bm VNW p12 l=1.3e-07 w=1.5e-07
MXP15 net107 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSQX4MTR Q VDD VNW VPW VSS CK D SE SI SN
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmrs SE net150 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net150 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net123 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 nmrs nmse net123 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN11 bm cn net141 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 NSN s net141 VPW n12 l=1.3e-07 w=1.5e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 nmrs SE net83 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net83 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 VDD SI net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net113 nmse nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 VDD pm m VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP12 VDD SN m VNW p12 l=1.3e-07 w=2.3e-07
MXP13 VDD SN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP16 net107 c bm VNW p12 l=1.3e-07 w=1.5e-07
MXP15 net107 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRHQX1MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 net142 SN VSS VPW n12 l=1.3e-07 w=4.1e-07
MXN12 net166 cn net142 VPW n12 l=1.3e-07 w=4.1e-07
MX_t25 pm nmsi net166 VPW n12 l=1.3e-07 w=4.1e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=4.3e-07
MXN14 net170 RN VSS VPW n12 l=1.3e-07 w=4.3e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP12 net111 c cn VNW p12 l=1.3e-07 w=4.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmsi net131 VNW p12 l=1.3e-07 w=3.1e-07
MX_t28 net131 c VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 m RN net117 VNW p12 l=1.3e-07 w=2.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.6e-07
MXP21 bm nmset net93 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSRHQX2MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 net142 SN VSS VPW n12 l=1.3e-07 w=5.9e-07
MXN19 net166 cn net142 VPW n12 l=1.3e-07 w=5.9e-07
MXN20 pm nmsi net166 VPW n12 l=1.3e-07 w=5.9e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=6.1e-07
MXN21 net170 RN VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP12 net111 c cn VNW p12 l=1.3e-07 w=4.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7e-07
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmsi net131 VNW p12 l=1.3e-07 w=4.5e-07
MXP22 net131 c VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 m RN net117 VNW p12 l=1.3e-07 w=2.3e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP23 bm nmset net93 VNW p12 l=1.3e-07 w=2.7e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRHQX4MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN20 net142 SN VSS VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net166 cn net142 VPW n12 l=1.3e-07 w=7.5e-07
MX_t25 pm nmsi net166 VPW n12 l=1.3e-07 w=7.5e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=7.2e-07
MXN21 net170 RN VSS VPW n12 l=1.3e-07 w=7.2e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN22 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP22 net111 c cn VNW p12 l=1.3e-07 w=5.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.2e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.9e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP23 pm nmsi net131 VNW p12 l=1.3e-07 w=6.8e-07
MX_t28 net131 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP26 m RN net117 VNW p12 l=1.3e-07 w=3.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP27 bm nmset net93 VNW p12 l=1.3e-07 w=3.6e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRHQX8MTR Q VDD VNW VPW VSS CK D RN SE SI SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI80_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g10_MXNA1_2 c nck VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g13_MXNA1 wlnmin D VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI71_MXNOE nmsi nmse wlnmin VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNOE nmsi SE XI1_n1 VPW n12 l=1.3e-07 w=2.6e-07
mXI1_MXNA1 XI1_n1 SI VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN20 net142 SN VSS VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net166 cn net142 VPW n12 l=1.3e-07 w=7.5e-07
MX_t25 pm nmsi net166 VPW n12 l=1.3e-07 w=7.5e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 m pm net170 VPW n12 l=1.3e-07 w=7.2e-07
MXN21 net170 RN VSS VPW n12 l=1.3e-07 w=7.2e-07
MX_t6 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN16 bm cn net162 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net162 RN net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN18 VSS s net159 VPW n12 l=1.3e-07 w=1.8e-07
MXN22 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP11 net111 CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP22 net111 c cn VNW p12 l=1.3e-07 w=5.2e-07
mXI80_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g13_MXPA1 wlnmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI71_MXPOEN nmsi SE wlnmin VNW p12 l=1.3e-07 w=3.2e-07
mXI1_MXPOEN nmsi nmse XI1_p1 VNW p12 l=1.3e-07 w=2.9e-07
mXI1_MXPA1 XI1_p1 SI VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP23 pm nmsi net131 VNW p12 l=1.3e-07 w=6.8e-07
MX_t28 net131 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP15 net117 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP26 m RN net117 VNW p12 l=1.3e-07 w=3.1e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP27 bm nmset net93 VNW p12 l=1.3e-07 w=3.6e-07
MXP17 net93 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP20 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP19 net105 nmset net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP18 VDD s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRX1MTR Q QN VDD VNW VPW VSS CK D RN SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE pm c XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MX_t15 NSN NRN m VPW n12 l=1.3e-07 w=1.9e-07
mXI60_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MXN5 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MX_t20 bm cn net75 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN s net75 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN pm cn XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 brn NRN VDD VNW p12 l=1.3e-07 w=4.9e-07
MX_t11 m pm brn VNW p12 l=1.3e-07 w=3.6e-07
MX_t12 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t16 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MXP6 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 brn s net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSRX2MTR Q QN VDD VNW VPW VSS CK D RN SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE pm c XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MX_t15 NSN NRN m VPW n12 l=1.3e-07 w=1.9e-07
mXI60_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MXN5 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MX_t20 bm cn net75 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN s net75 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN pm cn XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 brn NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP7 m pm brn VNW p12 l=1.3e-07 w=4.4e-07
MX_t12 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t16 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.4e-07
MXP6 bm c net105 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 brn s net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSRX4MTR Q QN VDD VNW VPW VSS CK D RN SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=2.5e-07
mXI8_MXNOE pm c XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MX_t15 NSN NRN m VPW n12 l=1.3e-07 w=1.9e-07
mXI60_MXNOE bm c m VPW n12 l=1.3e-07 w=4.7e-07
MXN5 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MX_t20 bm cn net91 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN s net91 VPW n12 l=1.3e-07 w=1.8e-07
MX_t14 NSN SN VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=3e-07
mXI8_MXPOEN pm cn XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 brn NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP7 m pm brn VNW p12 l=1.3e-07 w=4.4e-07
MX_t12 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t16 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI60_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.7e-07
MXP6 bm c net101 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 brn s net101 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSX1MTR Q QN VDD VNW VPW VSS CK D SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE pm c XI2_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNA1 XI2_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MX_t11 m pm BSN VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MX_t19 bm cn net138 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 BSN s net138 VPW n12 l=1.3e-07 w=1.8e-07
MX_t33 BSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI33_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN pm cn XI2_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPA1 XI2_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MX_t24 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 bm c net104 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 VDD s net104 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI33_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFSX2MTR Q QN VDD VNW VPW VSS CK D SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE pm c XI2_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNA1 XI2_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
MX_t11 m pm BSN VPW n12 l=1.3e-07 w=2.1e-07
MX_t11_2 m pm BSN VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MX_t19 bm cn net138 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN s net138 VPW n12 l=1.3e-07 w=1.5e-07
MX_t33 BSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN pm cn XI2_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPA1 XI2_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.4e-07
MX_t24 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm c net104 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD s net104 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI34_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFSX4MTR Q QN VDD VNW VPW VSS CK D SE SI SN
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE nmrs SE XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 D VSS VPW n12 l=1.3e-07 w=2e-07
mXI3_MXNOE nmrs nmse XI3_n1 VPW n12 l=1.3e-07 w=2e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=2e-07
mXI2_MXNOE pm c XI2_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNA1 XI2_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.8e-07
MX_t11 m pm BSN VPW n12 l=1.3e-07 w=3.5e-07
MX_t11_2 m pm BSN VPW n12 l=1.3e-07 w=3.5e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=5.2e-07
MX_t19 bm cn net138 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN s net138 VPW n12 l=1.3e-07 w=1.5e-07
MX_t33 BSN SN VSS VPW n12 l=1.3e-07 w=1.08e-06
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI35_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI35_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN nmrs SE XI3_p1 VNW p12 l=1.3e-07 w=2.8e-07
mXI3_MXPA1 XI3_p1 D VDD VNW p12 l=1.3e-07 w=2.8e-07
mXI0_MXPA1 XI0_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPOEN nmrs nmse XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.4e-07
mXI2_MXPOEN pm cn XI2_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPA1 XI2_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=7.8e-07
MX_t10 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
MX_t24 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm c net104 VNW p12 l=1.3e-07 w=1.5e-07
MXP5 VDD s net104 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.9e-07
mXI35_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI35_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFTRX1MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net074 RN VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN5 net181 D net074 VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net181 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net193 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net193 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE bm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net96 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP7 nmrs SE net96 VNW p12 l=1.3e-07 w=3e-07
MXP6 nmrs nmse net114 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net114 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net105 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmrs RN net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI43_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI8_MXPOEN bm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFTRX2MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net074 RN VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN5 net181 D net074 VPW n12 l=1.3e-07 w=2.4e-07
MX_t7 nmrs nmse net181 VPW n12 l=1.3e-07 w=2.4e-07
MX_t3 nmrs SE net193 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net193 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mXI43_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI8_MXNOE bm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI47_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net96 D VDD VNW p12 l=1.3e-07 w=3e-07
MXP7 nmrs SE net96 VNW p12 l=1.3e-07 w=3e-07
MXP6 nmrs nmse net114 VNW p12 l=1.3e-07 w=2.3e-07
MX_t1 net114 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net105 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 nmrs RN net105 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI43_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI8_MXPOEN bm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFTRX4MTR Q QN VDD VNW VPW VSS CK D RN SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net074 RN VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN8 net181 D net074 VPW n12 l=1.3e-07 w=4.2e-07
MX_t7 nmrs nmse net181 VPW n12 l=1.3e-07 w=4.2e-07
MX_t3 nmrs SE net193 VPW n12 l=1.3e-07 w=2.3e-07
MXN7 net193 SI VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI43_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI69_MXNOE pm cn nmrs VPW n12 l=1.3e-07 w=3.4e-07
mXI7_MXNOE pm c XI7_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 XI7_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=4e-07
mXI59_MXNOE bm c m VPW n12 l=1.3e-07 w=8e-07
mXI8_MXNOE bm cn XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI49_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI49_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 net96 D VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP11 nmrs SE net96 VNW p12 l=1.3e-07 w=5.4e-07
MXP10 nmrs nmse net114 VNW p12 l=1.3e-07 w=2.7e-07
MX_t1 net114 SI VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP8 net105 SE VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP13 nmrs RN net105 VNW p12 l=1.3e-07 w=2.7e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI43_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI69_MXPOEN pm c nmrs VNW p12 l=1.3e-07 w=4.1e-07
mXI7_MXPOEN pm cn XI7_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 XI7_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_3 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_4 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mXI59_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI59_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI8_MXPOEN bm c XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=4.3e-07
mXI49_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI49_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SDFFX1MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net137 SE net116 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net116 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net137 D net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 pm cn net137 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNOE pm c XI17_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 XI17_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI57_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI15_MXNOE sn c XI15_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI16_MXNOE sn cn XI16_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI16_MXNA1 XI16_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI58_MXNA1 Q sn VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 s sn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net77 nmse net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net73 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net76 SE VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net77 D net76 VNW p12 l=1.3e-07 w=3.8e-07
MXP4 pm c net77 VNW p12 l=1.3e-07 w=3.8e-07
mXI17_MXPOEN pm cn XI17_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPA1 XI17_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI57_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI15_MXPOEN sn cn XI15_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI16_MXPOEN sn c XI16_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI16_MXPA1 XI16_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s sn VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPA1 Q sn VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SDFFX2MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net137 SE net116 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net116 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net137 D net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 pm cn net137 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNOE pm c XI17_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 XI17_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI57_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI15_MXNOE sn c XI15_n1 VPW n12 l=1.3e-07 w=3.5e-07
mXI16_MXNOE sn cn XI16_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI16_MXNA1 XI16_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s sn VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI61_MXNA1 Q sn VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP5 net77 nmse net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net73 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net76 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net77 D net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm c net77 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPOEN pm cn XI17_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI17_MXPA1 XI17_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI57_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI15_MXPOEN sn cn XI15_p1 VNW p12 l=1.3e-07 w=4.9e-07
mXI16_MXPOEN sn c XI16_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI16_MXPA1 XI16_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s sn VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI61_MXPA1 Q sn VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT SDFFX4MTR Q QN VDD VNW VPW VSS CK D SE SI
mX_g8_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net137 SE net116 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net116 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net137 D net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 pm cn net137 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNOE pm c XI17_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 XI17_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI57_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=5.8e-07
mXI15_MXNOE sn c XI15_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI16_MXNOE sn cn XI16_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI16_MXNA1 XI16_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s sn VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI62_MXNA1 Q sn VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI62_MXNA1_2 Q sn VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g8_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP5 net77 nmse net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net73 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net76 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net77 D net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 pm c net77 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPOEN pm cn XI17_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI17_MXPA1 XI17_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=4.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI57_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI15_MXPOEN sn cn XI15_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI16_MXPOEN sn c XI16_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI16_MXPA1 XI16_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s sn VDD VNW p12 l=1.3e-07 w=4.2e-07
mXI62_MXPA1 Q sn VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI62_MXPA1_2 Q sn VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT SEDFFHQX1MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=2.3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=3.6e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.4e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=3e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP4 net079 c cn VNW p12 l=1.3e-07 w=4.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP5 pm nmsi net78 VNW p12 l=1.3e-07 w=4.4e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.4e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SEDFFHQX2MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=5.1e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=5.6e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=3.9e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP6 net079 c cn VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 pm nmsi net78 VNW p12 l=1.3e-07 w=6.2e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFHQX4MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=5.1e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=7e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.8e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 net079 c cn VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.8e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 pm nmsi net78 VNW p12 l=1.3e-07 w=6.2e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFHQX8MTR Q VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNA1 XI16_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI16_MXNOE nmsi SE XI16_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI65_MXNOE nmsi nmse2 nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g8_MXNA1 nmse2 se2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 se2 E XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA2 nmen2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNA1 nmen2 E VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 en2 nmen2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI8_MXNOE nmsi nmen2 XI8_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI8_MXNA1 XI8_n1 s VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t6 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 net0121 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 pm nmsi net0121 VPW n12 l=1.3e-07 w=5.1e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI93_MXNOE bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNOE bm cn XI13_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI13_MXNA1 XI13_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPA1 XI16_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI16_MXPOEN nmsi nmse XI16_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
mXI65_MXPOEN nmsi se2 nmin VNW p12 l=1.3e-07 w=7e-07
mX_g8_MXPA1 nmse2 se2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 se2 E VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 se2 nmse VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI7_MXPA2 XI7_p1 SE VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI7_MXPA1 nmen2 E XI7_p1 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 en2 nmen2 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI8_MXPOEN nmsi en2 XI8_p1 VNW p12 l=1.3e-07 w=2.8e-07
mXI8_MXPA1 XI8_p1 s VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t10 net079 CK VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 net079 c cn VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.8e-07
MXP0 net78 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 pm nmsi net78 VNW p12 l=1.3e-07 w=6.2e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI93_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPOEN bm c XI13_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI13_MXPA1 XI13_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFTRX1MTR Q QN VDD VNW VPW VSS CK D E RN SE SI
MX_t9 nmrs RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmrs SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI44_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmsi SI VSS VPW n12 l=1.3e-07 w=1.7e-07
mXI38_MXNOE nmin_pass2 bse nmsi VPW n12 l=1.3e-07 w=1.8e-07
mXI39_MXNOE nmin_pass2 nmse nmin_pass1 VPW n12 l=1.3e-07 w=1.8e-07
mXI45_MXNA1 bse nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNOE nmin_pass1 be nmin VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE nmin_pass1 nmen s VPW n12 l=1.3e-07 w=1.8e-07
mX_g12_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 be nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net169 nmrs VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t5 net169 nmin_pass2 VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t4 pm cn net169 VPW n12 l=1.3e-07 w=2e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g18_MXNA1 nm m VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI59_MXNOE bnm c nm VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNOE bnm cn XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI46_MXNA1 QN bnm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP4 nmrs RN net108 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net108 SE VDD VNW p12 l=1.3e-07 w=3e-07
mXI44_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmsi SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI38_MXPOEN nmin_pass2 nmse nmsi VNW p12 l=1.3e-07 w=2.3e-07
mXI39_MXPOEN nmin_pass2 bse nmin_pass1 VNW p12 l=1.3e-07 w=2.3e-07
mXI45_MXPA1 bse nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPOEN nmin_pass1 nmen nmin VNW p12 l=1.3e-07 w=2.3e-07
mXI40_MXPOEN nmin_pass1 be s VNW p12 l=1.3e-07 w=2.3e-07
mX_g12_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 be nmen VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
MX_t1 net102 nmrs VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net111 nmin_pass2 net102 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 pm c net111 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g18_MXPA1 nm m VDD VNW p12 l=1.3e-07 w=4.1e-07
mXI59_MXPOEN bnm cn nm VNW p12 l=1.3e-07 w=4.1e-07
mXI1_MXPOEN bnm c XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI46_MXPA1 QN bnm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SEDFFTRX2MTR Q QN VDD VNW VPW VSS CK D E RN SE SI
MX_t9 nmrs RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmrs SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI44_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmsi SI VSS VPW n12 l=1.3e-07 w=1.7e-07
mXI38_MXNOE nmin_pass2 bse nmsi VPW n12 l=1.3e-07 w=1.8e-07
mXI39_MXNOE nmin_pass2 nmse nmin_pass1 VPW n12 l=1.3e-07 w=1.8e-07
mXI45_MXNA1 bse nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNOE nmin_pass1 be nmin VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE nmin_pass1 nmen s VPW n12 l=1.3e-07 w=1.8e-07
mX_g12_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 be nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN5 net169 nmrs VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t5 net169 nmin_pass2 VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t4 pm cn net169 VPW n12 l=1.3e-07 w=2e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g18_MXNA1 nm m VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE bnm c nm VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNOE bnm cn XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI47_MXNA1 QN bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmrs RN net108 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net108 SE VDD VNW p12 l=1.3e-07 w=3e-07
mXI44_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmsi SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI38_MXPOEN nmin_pass2 nmse nmsi VNW p12 l=1.3e-07 w=2.3e-07
mXI39_MXPOEN nmin_pass2 bse nmin_pass1 VNW p12 l=1.3e-07 w=2.3e-07
mXI45_MXPA1 bse nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPOEN nmin_pass1 nmen nmin VNW p12 l=1.3e-07 w=2.3e-07
mXI40_MXPOEN nmin_pass1 be s VNW p12 l=1.3e-07 w=2.3e-07
mX_g12_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 be nmen VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.2e-07
MX_t1 net102 nmrs VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net111 nmin_pass2 net102 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 pm c net111 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g18_MXPA1 nm m VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI59_MXPOEN bnm cn nm VNW p12 l=1.3e-07 w=5.9e-07
mXI1_MXPOEN bnm c XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI47_MXPA1 QN bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFTRX4MTR Q QN VDD VNW VPW VSS CK D E RN SE SI
MX_t9 nmrs RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmrs SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI44_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmsi SI VSS VPW n12 l=1.3e-07 w=1.7e-07
mXI38_MXNOE nmin_pass2 bse nmsi VPW n12 l=1.3e-07 w=1.8e-07
mXI39_MXNOE nmin_pass2 nmse nmin_pass1 VPW n12 l=1.3e-07 w=1.8e-07
mXI45_MXNA1 bse nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNOE nmin_pass1 be nmin VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE nmin_pass1 nmen s VPW n12 l=1.3e-07 w=1.8e-07
mX_g12_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 be nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN5 net169 nmrs VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t5 net169 nmin_pass2 VSS VPW n12 l=1.3e-07 w=2.3e-07
MX_t4 pm cn net169 VPW n12 l=1.3e-07 w=2e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g18_MXNA1 nm m VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI59_MXNOE bnm c nm VPW n12 l=1.3e-07 w=7.4e-07
mXI1_MXNOE bnm cn XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI48_MXNA1 QN bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI48_MXNA1_2 QN bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmrs RN net108 VNW p12 l=1.3e-07 w=3e-07
MX_t7 net108 SE VDD VNW p12 l=1.3e-07 w=3e-07
mXI44_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 nmsi SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI38_MXPOEN nmin_pass2 nmse nmsi VNW p12 l=1.3e-07 w=2.3e-07
mXI39_MXPOEN nmin_pass2 bse nmin_pass1 VNW p12 l=1.3e-07 w=2.3e-07
mXI45_MXPA1 bse nmse VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPOEN nmin_pass1 nmen nmin VNW p12 l=1.3e-07 w=2.3e-07
mXI40_MXPOEN nmin_pass1 be s VNW p12 l=1.3e-07 w=2.3e-07
mX_g12_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 be nmen VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t1 net102 nmrs VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net111 nmin_pass2 net102 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 pm c net111 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.9e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g18_MXPA1 nm m VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI59_MXPOEN bnm cn nm VNW p12 l=1.3e-07 w=8e-07
mXI1_MXPOEN bnm c XI1_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI48_MXPA1 QN bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI48_MXPA1_2 QN bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFX1MTR Q QN VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net180 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net187 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net190 SE net187 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net190 D net181 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net181 E net180 VPW n12 l=1.3e-07 w=1.8e-07
MX_t16 net196 nmen net180 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net196 s net190 VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 pm cn net190 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI3_MXNOE nm c XI3_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI4_MXNOE nm cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI41_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t6 net85 SE VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t8 net97 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net96 nmse net97 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net96 D net91 VNW p12 l=1.3e-07 w=4.7e-07
MX_t5 net91 nmen net85 VNW p12 l=1.3e-07 w=4.7e-07
MXP9 net88 E net85 VNW p12 l=1.3e-07 w=4.7e-07
MXP10 net88 s net96 VNW p12 l=1.3e-07 w=4.7e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm c net96 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI40_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI3_MXPOEN nm cn XI3_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI4_MXPOEN nm c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.4e-07
mXI41_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SEDFFX2MTR Q QN VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net100 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net92 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net88 SE net92 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net88 D net76 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net76 E net100 VPW n12 l=1.3e-07 w=1.8e-07
MX_t16 net84 nmen net100 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net84 s net88 VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 pm cn net88 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI3_MXNOE nm c XI3_n1 VPW n12 l=1.3e-07 w=4.4e-07
mXI4_MXNOE nm cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI42_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t6 net127 SE VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t8 net111 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net113 nmse net111 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net113 D net131 VNW p12 l=1.3e-07 w=4.7e-07
MX_t5 net131 nmen net127 VNW p12 l=1.3e-07 w=4.7e-07
MXP9 net105 E net127 VNW p12 l=1.3e-07 w=4.7e-07
MXP10 net105 s net113 VNW p12 l=1.3e-07 w=4.7e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm c net113 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI40_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI3_MXPOEN nm cn XI3_p1 VNW p12 l=1.3e-07 w=5.4e-07
mXI4_MXPOEN nm c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI42_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SEDFFX4MTR Q QN VDD VNW VPW VSS CK D E SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net100 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net92 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net88 SE net92 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net88 D net76 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net76 E net100 VPW n12 l=1.3e-07 w=1.8e-07
MX_t16 net84 nmen net100 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net84 s net88 VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 pm cn net88 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI40_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI3_MXNOE nm c XI3_n1 VPW n12 l=1.3e-07 w=6.4e-07
mXI4_MXNOE nm cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI43_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI43_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 net127 SE VDD VNW p12 l=1.3e-07 w=2.4e-07
MXP14_2 net127 SE VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t8 net111 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 net113 nmse net111 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net113 D net131 VNW p12 l=1.3e-07 w=4.7e-07
MX_t5 net131 nmen net127 VNW p12 l=1.3e-07 w=4.7e-07
MXP12 net105 E net127 VNW p12 l=1.3e-07 w=4.6e-07
MXP13 net105 s net113 VNW p12 l=1.3e-07 w=4.6e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 pm c net113 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI40_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI3_MXPOEN nm cn XI3_p1 VNW p12 l=1.3e-07 w=7.3e-07
mXI4_MXPOEN nm c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI43_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI43_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SMDFFHQX1MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=1.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=2.1e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN4 VSS cn net107 VPW n12 l=1.3e-07 w=3.3e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=3.3e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=3.7e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=2.6e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=2.6e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=3e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=3e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=4.2e-07
MXP0 cn c net085 VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=4e-07
MXP3 pm nmsi net060 VNW p12 l=1.3e-07 w=4e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=7.3e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT SMDFFHQX2MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=1.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=3.1e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=3e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN5 VSS cn net107 VPW n12 l=1.3e-07 w=4.8e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=4.8e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=4.4e-07
MXP4 cn c net085 VNW p12 l=1.3e-07 w=4.4e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP5 pm nmsi net060 VNW p12 l=1.3e-07 w=5.9e-07
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=9.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=9.8e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SMDFFHQX4MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=2.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=5e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN6 VSS cn net107 VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=5.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=3.4e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net085 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net060 VNW p12 l=1.3e-07 w=1.01e-06
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT SMDFFHQX8MTR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
mX_g9_MXNA1 nmse SE VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 XI24_n1 SI VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI24_MXNOE nmsi SE XI24_n1 VPW n12 l=1.3e-07 w=2.8e-07
MX_t8 nmsi nn1 d1n VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 d1n D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g8_MXNA1 nn1 n1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 n1 S0 net119 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net119 nmse VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 n2 SE VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 n2 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 nn2 n2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi n2 d0n VPW n12 l=1.3e-07 w=5e-07
mX_g16_MXNA1 d0n D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN6 VSS cn net107 VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net107 VPW n12 l=1.3e-07 w=5.6e-07
mXI23_MXNOE pm c XI23_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA1 XI23_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI22_MXNOE bm cn XI22_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 XI22_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXPA1 nmse SE VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI24_MXPA1 XI24_p1 SI VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI24_MXPOEN nmsi nmse XI24_p1 VNW p12 l=1.3e-07 w=3.4e-07
mX_g13_MXPA1 d1n D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t9 d1n n1 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g8_MXPA1 nn1 n1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t38 VDD S0 n1 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD nmse n1 VNW p12 l=1.3e-07 w=2.3e-07
MX_t43 VDD SE net85 VNW p12 l=1.3e-07 w=3.6e-07
MXP1 net85 S0 n2 VNW p12 l=1.3e-07 w=3.6e-07
mX_g6_MXPA1 nn2 n2 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 d0n nn2 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 d0n D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net085 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net085 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net060 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net060 VNW p12 l=1.3e-07 w=1.01e-06
mXI23_MXPOEN pm cn XI23_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI23_MXPA1 XI23_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI22_MXPOEN bm c XI22_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 XI22_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


