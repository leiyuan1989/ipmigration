* 
* No part of this file can be released without the consent of SMIC.
*
* Note: SMIC recommends that users set VNTOL=1E-9 at .option for more smooth convergence.
*************************************************************************************************************
* 0.18um Mixed Signal 1P6M with MIM Salicide 1.8V/3.3V RF SPICE Model (for HSPICE only)  *
*************************************************************************************************************
*
* Release version    : 1.5
*
* Release date       : 01/20/2007
*
* Simulation tool    : Synopsys Star-HSPICE version 2005.9
*
*
*  Inductor   :
*
*        *------------------------------------------* 
*        | Inductor subckt |   diff_ind_rf    |
*        *------------------------------------------*
**********************************
* 0.18um differential Inductor *
**********************************
* 1=port1(M6), 2=port2(M5)
* R means inner redius; N means turns
* Spacing is fixed at 1.5um and width is fixed at 8um
.subckt diff_ind_rf 1 2 R=radius N=turns
* inductor scalable model parameters
.param
+L00  = 'max(((-0.00043*R*1E+6+0.0326)*N*N*N+(0.00798*R*1E+6-0.4421)*N*N+(-0.0296*R*1E+6+1.95)*N+(0.0437*R*1E+6-2.5533))*1E-9, 1E-12)'
+R00  = 'max((-0.0005414*R*1E+6+0.022909)*N*N*N+(0.0091377*R*1E+6-0.359131)*N*N+(-0.0398784*R*1E+6+2.084685)*N+(0.0643148*R*1E+6-2.873445), 1E-6)'
+L01  = '1.33E-010'
+R01  = '125'
+L10  = 'max(((-0.00043*R*1E+6+0.0326)*N*N*N+(0.00798*R*1E+6-0.4421)*N*N+(-0.0296*R*1E+6+1.95)*N+(0.0437*R*1E+6-2.5533))*1E-9, 1E-12)'
+R10  = 'max((-0.0005414*R*1E+6+0.022909)*N*N*N+(0.0091377*R*1E+6-0.359131)*N*N+(-0.0398784*R*1E+6+2.084685)*N+(0.0643148*R*1E+6-2.873445), 1E-6)'
+L11  = '1.33E-010'
+R11  = '125'
+COXM   = 'max((0.67851*L00*L00*L00*1E+9*1E+9*1E+9-8.27182*L00*L00*1E+9*1E+9+34.35047*L00*1E+9+30.06634)*1E-15, 1E-18)'
+RSM    = 'max((42.31593*L00*L00*L00*1E+9*1E+9*1E+9-411.80075*L00*L00*1E+9*1E+9+1389.18524*L00*1E+9+1419.43733), 1E-6)'
+CSM    = 'max((0.1322*L00*L00*L00*1E+9*1E+9*1E+9-1.7049*L00*L00*1E+9*1E+9+9.96*L00*1E+9-1.3483)*1E-15, 1E-18)'
+CPASS  = 'max(((-0.0068648*R*1E+6+0.732611)*N*N*N+(0.1468104*R*1E+6-10.650026)*N*N+(-0.697329*R*1E+6+51.120355)*N+(1.1635258*R*1E+6-82.029203))*1E-15, 1E-18)'
+CCI    = 'max(((0.012491*R*1E+6-0.569096)*N*N*N+(-0.20918*R*1E+6+6.17064)*N*N+(0.913908*R*1E+6+9.895997)*N+(-0.14843*R*1E+6-95.477512))*1E-15, 1E-18)'
+CCO    = 'max(((0.012491*R*1E+6-0.569096)*N*N*N+(-0.20918*R*1E+6+6.17064)*N*N+(0.913908*R*1E+6+9.895997)*N+(-0.14843*R*1E+6-95.477512))*1E-15, 1E-18)'
+RCI    = 'max((49.11941*L00*L00*L00*1E+9*1E+9*1E+9-503.65103*L00*L00*1E+9*1E+9+1625.77739*L00*1E+9+1312.52424), 1E-6)'
+RCO    = 'max((49.11941*L00*L00*L00*1E+9*1E+9*1E+9-503.65103*L00*L00*1E+9*1E+9+1625.77739*L00*1E+9+1312.52424), 1E-6)'
+COXI   = 'max(((-0.020551*R*1E+6+1.147253)*N*N+(0.194817*R*1E+6-1.934667)*N+(-0.108661*R*1E+6-12.53573))*1E-15, 1E-18)'
+RSI    = 'max((13.34945*L00*L00*L00*1E+9*1E+9*1E+9-135.42118*L00*L00*1E+9*1E+9+436.81570*L00*1E+9+319.07449), 1E-6)'
+CSI    = 'max(((0.00202687*R*1E+6-0.009606)*N*N*N+(-0.040912*R*1E+6-0.125553)*N*N+(0.209166*R*1E+6+7.262962)*N+(-0.105972*R*1E+6-22.808747))*1E-15, 1E-18)'
+COXO   = 'max(((-0.020551*R*1E+6+1.147253)*N*N+(0.194817*R*1E+6-1.934667)*N+(-0.108661*R*1E+6-12.53573))*1E-15, 1E-18)'
+RSO    = 'max((13.34945*L00*L00*L00*1E+9*1E+9*1E+9-135.42118*L00*L00*1E+9*1E+9+436.81570*L00*1E+9+319.07449), 1E-6)'
+CSO    = 'max(((0.00202687*R*1E+6-0.009606)*N*N*N+(-0.040912*R*1E+6-0.125553)*N*N+(0.209166*R*1E+6+7.262962)*N+(-0.105972*R*1E+6-22.808747))*1E-15, 1E-18)'
* equivalent circuit
L00_rf  1 N1 L00 
R00_rf  N1 NM R00  
L01_rf  N1 N11 L01 
R01_rf  N11 NM R01  
L10_rf  NM N2 L10  
R10_rf  N2 2 R10  
L11_rf  N2 N21 L11 
R11_rf  N21 2 R11   
COXM_rf  NM NSM COXM  
RSM_rf  NSM 0 RSM  
CSM_rf  NSM 0 CSM 
CPASS_rf  1 2 CPASS 
CCI_rf  1 NM CCI 
CCO_rf  NM 2 CCO  
RCI_rf  NSI NSM RCI  
RCO_rf  NSM NSO RCO  
COXI_rf 1 NSI COXI  
RSI_rf  NSI 0 RSI  
CSI_rf  NSI 0 CSI  
COXO_rf 2 NSO COXO  
RSO_rf  NSO 0 RSO  
CSO_rf  NSO 0 CSO
K01 L10_rf L01_rf 0.205
K11 L00_rf L11_rf 0.205
.ends diff_ind_rf
