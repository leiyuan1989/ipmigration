* ---------------------------------------------------------------------------- 
* 
*     library Calibre-based CDL file 
* 
*     Date: Feb 19, 2010 11:19:35 PM IST 
* 
*     CellBuilder version 3.2.3 -- built on Dec 04, 2009 
*     Copyright (c) 2002-2009 ARM, Inc. 
*     The confidential and proprietary information contained in this file 
*     may only be used by a person authorised under and to the extent 
*     permitted by a subsisting licensing agreement from ARM Limited. 
*      
*     (C) COPYRIGHT 2004-2010 ARM Limited. 
*     ALL RIGHTS RESERVED 
*      
*     This entire notice must be reproduced on all copies of this file 
*     and copies of this file may only be made by a person if such person 
*     is permitted to do so under the terms of a subsisting license 
*     agreement from ARM Limited. 
* 
* ----------------------------------------------------------------------------



.SUBCKT A2SDFFQN_X0P5M_A9TR QN VDD VNW VPW VSS A B CK SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 22 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 22 VPW nch L=4e-08 W=1.2e-07 
M3 23 3 VSS VPW nch L=4e-08 W=2.45e-07 
M4 6 B 23 VPW nch L=4e-08 W=2.45e-07 
M5 4 A 6 VPW nch L=4e-08 W=2.45e-07 
M6 7 13 4 VPW nch L=4e-08 W=1.2e-07 
M7 24 12 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 8 24 VPW nch L=4e-08 W=1.2e-07 
M9 8 7 VSS VPW nch L=4e-08 W=1.2e-07 
M10 9 12 8 VPW nch L=4e-08 W=1.2e-07 
M11 25 13 9 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 10 25 VPW nch L=4e-08 W=1.2e-07 
M13 VSS 9 10 VPW nch L=4e-08 W=1.2e-07 
M14 QN 9 VSS VPW nch L=4e-08 W=1.55e-07 
M15 VSS 13 12 VPW nch L=4e-08 W=1.2e-07 
M16 13 CK VSS VPW nch L=4e-08 W=1.2e-07 
M17 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M18 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M19 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M20 5 SE VDD VNW pch L=4e-08 W=2.55e-07 
M21 4 B 5 VNW pch L=4e-08 W=2.55e-07 
M22 4 A 5 VNW pch L=4e-08 W=2.55e-07 
M23 7 12 4 VNW pch L=4e-08 W=1.2e-07 
M24 20 13 7 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M26 8 7 VDD VNW pch L=4e-08 W=1.8e-07 
M27 9 13 8 VNW pch L=4e-08 W=1.2e-07 
M28 21 12 9 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 10 21 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 9 10 VNW pch L=4e-08 W=1.2e-07 
M31 QN 9 VDD VNW pch L=4e-08 W=2e-07 
M32 VDD 13 12 VNW pch L=4e-08 W=2.5e-07 
M33 13 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT A2SDFFQN_X1M_A9TR QN VDD VNW VPW VSS A B CK SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 22 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 22 VPW nch L=4e-08 W=1.2e-07 
M3 23 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 6 B 23 VPW nch L=4e-08 W=3.1e-07 
M5 4 A 6 VPW nch L=4e-08 W=3.1e-07 
M6 7 13 4 VPW nch L=4e-08 W=1.6e-07 
M7 24 12 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 8 24 VPW nch L=4e-08 W=1.2e-07 
M9 8 7 VSS VPW nch L=4e-08 W=1.6e-07 
M10 9 12 8 VPW nch L=4e-08 W=1.6e-07 
M11 25 13 9 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 10 25 VPW nch L=4e-08 W=1.2e-07 
M13 VSS 9 10 VPW nch L=4e-08 W=1.2e-07 
M14 QN 9 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 13 12 VPW nch L=4e-08 W=1.2e-07 
M16 13 CK VSS VPW nch L=4e-08 W=1.2e-07 
M17 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M18 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M19 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M20 5 SE VDD VNW pch L=4e-08 W=3.1e-07 
M21 4 B 5 VNW pch L=4e-08 W=3.1e-07 
M22 4 A 5 VNW pch L=4e-08 W=3.1e-07 
M23 7 12 4 VNW pch L=4e-08 W=1.6e-07 
M24 20 13 7 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M26 8 7 VDD VNW pch L=4e-08 W=2.3e-07 
M27 9 13 8 VNW pch L=4e-08 W=1.6e-07 
M28 21 12 9 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 10 21 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 9 10 VNW pch L=4e-08 W=1.2e-07 
M31 QN 9 VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD 13 12 VNW pch L=4e-08 W=2.5e-07 
M33 13 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT A2SDFFQN_X2M_A9TR QN VDD VNW VPW VSS A B CK SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 22 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 22 VPW nch L=4e-08 W=1.2e-07 
M3 23 3 VSS VPW nch L=4e-08 W=3.5e-07 
M4 6 B 23 VPW nch L=4e-08 W=3.5e-07 
M5 4 A 6 VPW nch L=4e-08 W=3.5e-07 
M6 7 13 4 VPW nch L=4e-08 W=2.5e-07 
M7 24 12 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 8 24 VPW nch L=4e-08 W=1.2e-07 
M9 8 7 VSS VPW nch L=4e-08 W=2.5e-07 
M10 9 12 8 VPW nch L=4e-08 W=2.5e-07 
M11 25 13 9 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 10 25 VPW nch L=4e-08 W=1.2e-07 
M13 VSS 9 10 VPW nch L=4e-08 W=1.2e-07 
M14 QN 9 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 9 QN VPW nch L=4e-08 W=3.1e-07 
M16 VSS 13 12 VPW nch L=4e-08 W=1.3e-07 
M17 13 CK VSS VPW nch L=4e-08 W=1.3e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M21 5 SE VDD VNW pch L=4e-08 W=3.4e-07 
M22 4 B 5 VNW pch L=4e-08 W=3.4e-07 
M23 4 A 5 VNW pch L=4e-08 W=3.4e-07 
M24 7 12 4 VNW pch L=4e-08 W=2.5e-07 
M25 20 13 7 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M27 8 7 VDD VNW pch L=4e-08 W=3.2e-07 
M28 9 13 8 VNW pch L=4e-08 W=2.5e-07 
M29 21 12 9 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 10 21 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 9 10 VNW pch L=4e-08 W=1.2e-07 
M32 QN 9 VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD 9 QN VNW pch L=4e-08 W=3.8e-07 
M34 VDD 13 12 VNW pch L=4e-08 W=2.7e-07 
M35 13 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT A2SDFFQN_X3M_A9TR QN VDD VNW VPW VSS A B CK SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 22 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 22 VPW nch L=4e-08 W=1.2e-07 
M3 23 3 VSS VPW nch L=4e-08 W=3.5e-07 
M4 6 B 23 VPW nch L=4e-08 W=3.5e-07 
M5 4 A 6 VPW nch L=4e-08 W=3.5e-07 
M6 7 13 4 VPW nch L=4e-08 W=3.1e-07 
M7 24 12 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 8 24 VPW nch L=4e-08 W=1.2e-07 
M9 8 7 VSS VPW nch L=4e-08 W=3.1e-07 
M10 9 12 8 VPW nch L=4e-08 W=2.75e-07 
M11 25 13 9 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 10 25 VPW nch L=4e-08 W=1.2e-07 
M13 VSS 9 10 VPW nch L=4e-08 W=1.2e-07 
M14 QN 9 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 9 QN VPW nch L=4e-08 W=3.1e-07 
M16 QN 9 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 13 12 VPW nch L=4e-08 W=1.4e-07 
M18 13 CK VSS VPW nch L=4e-08 W=1.4e-07 
M19 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M20 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M21 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M22 5 SE VDD VNW pch L=4e-08 W=3.4e-07 
M23 4 B 5 VNW pch L=4e-08 W=3.4e-07 
M24 4 A 5 VNW pch L=4e-08 W=3.4e-07 
M25 7 12 4 VNW pch L=4e-08 W=3.1e-07 
M26 20 13 7 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M28 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M29 9 13 8 VNW pch L=4e-08 W=3.1e-07 
M30 21 12 9 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 10 21 VNW pch L=4e-08 W=1.2e-07 
M32 VDD 9 10 VNW pch L=4e-08 W=1.2e-07 
M33 QN 9 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 9 QN VNW pch L=4e-08 W=3.8e-07 
M35 QN 9 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 13 12 VNW pch L=4e-08 W=2.9e-07 
M37 13 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT A2SDFFQ_X0P5M_A9TR Q VDD VNW VPW VSS A B CK SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 22 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 22 VPW nch L=4e-08 W=1.2e-07 
M3 23 3 VSS VPW nch L=4e-08 W=2.5e-07 
M4 6 B 23 VPW nch L=4e-08 W=2.5e-07 
M5 4 A 6 VPW nch L=4e-08 W=2.5e-07 
M6 7 13 4 VPW nch L=4e-08 W=1.2e-07 
M7 24 12 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 8 24 VPW nch L=4e-08 W=1.2e-07 
M9 8 7 VSS VPW nch L=4e-08 W=1.2e-07 
M10 9 12 8 VPW nch L=4e-08 W=1.2e-07 
M11 25 13 9 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 10 25 VPW nch L=4e-08 W=1.2e-07 
M13 VSS 9 10 VPW nch L=4e-08 W=1.2e-07 
M14 Q 10 VSS VPW nch L=4e-08 W=1.55e-07 
M15 VSS 13 12 VPW nch L=4e-08 W=1.2e-07 
M16 13 CK VSS VPW nch L=4e-08 W=1.2e-07 
M17 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M18 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M19 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M20 5 SE VDD VNW pch L=4e-08 W=2.5e-07 
M21 4 B 5 VNW pch L=4e-08 W=2.5e-07 
M22 4 A 5 VNW pch L=4e-08 W=2.5e-07 
M23 7 12 4 VNW pch L=4e-08 W=1.2e-07 
M24 20 13 7 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M26 8 7 VDD VNW pch L=4e-08 W=1.55e-07 
M27 9 13 8 VNW pch L=4e-08 W=1.2e-07 
M28 21 12 9 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 10 21 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 9 10 VNW pch L=4e-08 W=1.55e-07 
M31 Q 10 VDD VNW pch L=4e-08 W=2e-07 
M32 VDD 13 12 VNW pch L=4e-08 W=2.5e-07 
M33 13 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT A2SDFFQ_X1M_A9TR Q VDD VNW VPW VSS A B CK SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 22 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 22 VPW nch L=4e-08 W=1.2e-07 
M3 23 3 VSS VPW nch L=4e-08 W=3.2e-07 
M4 6 B 23 VPW nch L=4e-08 W=3.2e-07 
M5 4 A 6 VPW nch L=4e-08 W=3.2e-07 
M6 7 13 4 VPW nch L=4e-08 W=1.6e-07 
M7 24 12 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 8 24 VPW nch L=4e-08 W=1.2e-07 
M9 8 7 VSS VPW nch L=4e-08 W=1.6e-07 
M10 9 12 8 VPW nch L=4e-08 W=1.6e-07 
M11 25 13 9 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 10 25 VPW nch L=4e-08 W=1.2e-07 
M13 VSS 9 10 VPW nch L=4e-08 W=1.75e-07 
M14 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 13 12 VPW nch L=4e-08 W=1.2e-07 
M16 13 CK VSS VPW nch L=4e-08 W=1.2e-07 
M17 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M18 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M19 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M20 5 SE VDD VNW pch L=4e-08 W=3e-07 
M21 4 B 5 VNW pch L=4e-08 W=3e-07 
M22 4 A 5 VNW pch L=4e-08 W=3e-07 
M23 7 12 4 VNW pch L=4e-08 W=1.6e-07 
M24 20 13 7 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M26 8 7 VDD VNW pch L=4e-08 W=2.05e-07 
M27 9 13 8 VNW pch L=4e-08 W=1.6e-07 
M28 21 12 9 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 10 21 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 9 10 VNW pch L=4e-08 W=2.45e-07 
M31 Q 10 VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD 13 12 VNW pch L=4e-08 W=2.5e-07 
M33 13 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT A2SDFFQ_X2M_A9TR Q VDD VNW VPW VSS A B CK SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 22 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 22 VPW nch L=4e-08 W=1.2e-07 
M3 23 3 VSS VPW nch L=4e-08 W=3.6e-07 
M4 6 B 23 VPW nch L=4e-08 W=3.6e-07 
M5 4 A 6 VPW nch L=4e-08 W=3.6e-07 
M6 7 13 4 VPW nch L=4e-08 W=2.5e-07 
M7 24 12 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 8 24 VPW nch L=4e-08 W=1.2e-07 
M9 8 7 VSS VPW nch L=4e-08 W=2.5e-07 
M10 9 12 8 VPW nch L=4e-08 W=2.5e-07 
M11 25 13 9 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 10 25 VPW nch L=4e-08 W=1.2e-07 
M13 VSS 9 10 VPW nch L=4e-08 W=2.5e-07 
M14 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 10 Q VPW nch L=4e-08 W=3.1e-07 
M16 VSS 13 12 VPW nch L=4e-08 W=1.3e-07 
M17 13 CK VSS VPW nch L=4e-08 W=1.3e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M21 5 SE VDD VNW pch L=4e-08 W=3.3e-07 
M22 4 B 5 VNW pch L=4e-08 W=3.3e-07 
M23 4 A 5 VNW pch L=4e-08 W=3.3e-07 
M24 7 12 4 VNW pch L=4e-08 W=2.5e-07 
M25 20 13 7 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M27 8 7 VDD VNW pch L=4e-08 W=3.1e-07 
M28 9 13 8 VNW pch L=4e-08 W=2.5e-07 
M29 21 12 9 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 10 21 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 9 10 VNW pch L=4e-08 W=3.8e-07 
M32 Q 10 VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD 10 Q VNW pch L=4e-08 W=3.8e-07 
M34 VDD 13 12 VNW pch L=4e-08 W=2.7e-07 
M35 13 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT A2SDFFQ_X3M_A9TR Q VDD VNW VPW VSS A B CK SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 22 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 22 VPW nch L=4e-08 W=1.2e-07 
M3 23 3 VSS VPW nch L=4e-08 W=3.6e-07 
M4 6 B 23 VPW nch L=4e-08 W=3.6e-07 
M5 4 A 6 VPW nch L=4e-08 W=3.6e-07 
M6 7 13 4 VPW nch L=4e-08 W=3.1e-07 
M7 24 12 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 8 24 VPW nch L=4e-08 W=1.2e-07 
M9 8 7 VSS VPW nch L=4e-08 W=3.5e-07 
M10 9 12 8 VPW nch L=4e-08 W=3.1e-07 
M11 25 13 9 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 10 25 VPW nch L=4e-08 W=1.2e-07 
M13 VSS 9 10 VPW nch L=4e-08 W=2.5e-07 
M14 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 10 Q VPW nch L=4e-08 W=3.1e-07 
M16 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 13 12 VPW nch L=4e-08 W=1.4e-07 
M18 13 CK VSS VPW nch L=4e-08 W=1.4e-07 
M19 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M20 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M21 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M22 5 SE VDD VNW pch L=4e-08 W=3.3e-07 
M23 4 B 5 VNW pch L=4e-08 W=3.3e-07 
M24 4 A 5 VNW pch L=4e-08 W=3.3e-07 
M25 7 12 4 VNW pch L=4e-08 W=3.1e-07 
M26 20 13 7 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M28 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M29 9 13 8 VNW pch L=4e-08 W=3.1e-07 
M30 21 12 9 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 10 21 VNW pch L=4e-08 W=1.2e-07 
M32 VDD 9 10 VNW pch L=4e-08 W=3.8e-07 
M33 Q 10 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 10 Q VNW pch L=4e-08 W=3.8e-07 
M35 Q 10 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 13 12 VNW pch L=4e-08 W=2.9e-07 
M37 13 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT A2SDFFQ_X4M_A9TR Q VDD VNW VPW VSS A B CK SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 22 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 22 VPW nch L=4e-08 W=1.2e-07 
M3 23 3 VSS VPW nch L=4e-08 W=3.6e-07 
M4 6 B 23 VPW nch L=4e-08 W=3.6e-07 
M5 4 A 6 VPW nch L=4e-08 W=3.6e-07 
M6 7 13 4 VPW nch L=4e-08 W=3.1e-07 
M7 24 12 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 8 24 VPW nch L=4e-08 W=1.2e-07 
M9 8 7 VSS VPW nch L=4e-08 W=3.5e-07 
M10 9 12 8 VPW nch L=4e-08 W=3.1e-07 
M11 25 13 9 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 10 25 VPW nch L=4e-08 W=1.2e-07 
M13 10 9 VSS VPW nch L=4e-08 W=2.5e-07 
M14 VSS 9 10 VPW nch L=4e-08 W=2.5e-07 
M15 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 10 Q VPW nch L=4e-08 W=3.1e-07 
M17 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M18 VSS 10 Q VPW nch L=4e-08 W=3.1e-07 
M19 VSS 13 12 VPW nch L=4e-08 W=1.4e-07 
M20 13 CK VSS VPW nch L=4e-08 W=1.4e-07 
M21 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M22 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M23 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M24 5 SE VDD VNW pch L=4e-08 W=3.3e-07 
M25 4 B 5 VNW pch L=4e-08 W=3.3e-07 
M26 4 A 5 VNW pch L=4e-08 W=3.3e-07 
M27 7 12 4 VNW pch L=4e-08 W=3.1e-07 
M28 20 13 7 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M30 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M31 9 13 8 VNW pch L=4e-08 W=3.1e-07 
M32 21 12 9 VNW pch L=4e-08 W=1.2e-07 
M33 VDD 10 21 VNW pch L=4e-08 W=1.2e-07 
M34 10 9 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 9 10 VNW pch L=4e-08 W=3.8e-07 
M36 Q 10 VDD VNW pch L=4e-08 W=3.8e-07 
M37 VDD 10 Q VNW pch L=4e-08 W=3.8e-07 
M38 Q 10 VDD VNW pch L=4e-08 W=3.8e-07 
M39 VDD 10 Q VNW pch L=4e-08 W=3.8e-07 
M40 VDD 13 12 VNW pch L=4e-08 W=2.9e-07 
M41 13 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT ADDFCIN_X1M_A9TR CO SUM VDD VNW VPW VSS A B CIN
M0 VSS 4 1 VPW nch L=4e-08 W=3.15e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.15e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.15e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.15e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.15e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.15e-07 
M6 7 B VSS VPW nch L=4e-08 W=1.55e-07 
M7 9 5 8 VPW nch L=4e-08 W=1.55e-07 
M8 7 6 9 VPW nch L=4e-08 W=1.55e-07 
M9 11 6 8 VPW nch L=4e-08 W=1.55e-07 
M10 10 5 11 VPW nch L=4e-08 W=1.55e-07 
M11 VSS 10 8 VPW nch L=4e-08 W=1.55e-07 
M12 10 CIN VSS VPW nch L=4e-08 W=1.55e-07 
M13 VSS 11 SUM VPW nch L=4e-08 W=2.95e-07 
M14 CO 9 VSS VPW nch L=4e-08 W=2.95e-07 
M15 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M16 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M17 5 B 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 7 5 VNW pch L=4e-08 W=3.8e-07 
M19 6 7 1 VNW pch L=4e-08 W=3.8e-07 
M20 4 B 6 VNW pch L=4e-08 W=3.8e-07 
M21 7 B VDD VNW pch L=4e-08 W=2.6e-07 
M22 9 5 7 VNW pch L=4e-08 W=2.6e-07 
M23 8 6 9 VNW pch L=4e-08 W=2.6e-07 
M24 11 6 10 VNW pch L=4e-08 W=2.6e-07 
M25 8 5 11 VNW pch L=4e-08 W=2.6e-07 
M26 VDD 10 8 VNW pch L=4e-08 W=2.6e-07 
M27 10 CIN VDD VNW pch L=4e-08 W=2.6e-07 
M28 VDD 11 SUM VNW pch L=4e-08 W=3.8e-07 
M29 CO 9 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT ADDFCIN_X1P4M_A9TR CO SUM VDD VNW VPW VSS A B CIN
M0 VSS 4 1 VPW nch L=4e-08 W=3.15e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.15e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.15e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.15e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.15e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.15e-07 
M6 7 B VSS VPW nch L=4e-08 W=2.3e-07 
M7 9 5 8 VPW nch L=4e-08 W=2.3e-07 
M8 7 6 9 VPW nch L=4e-08 W=2.3e-07 
M9 11 6 8 VPW nch L=4e-08 W=2.3e-07 
M10 10 5 11 VPW nch L=4e-08 W=2.3e-07 
M11 VSS 10 8 VPW nch L=4e-08 W=2.3e-07 
M12 10 CIN VSS VPW nch L=4e-08 W=2.3e-07 
M13 SUM 11 VSS VPW nch L=4e-08 W=2.2e-07 
M14 VSS 11 SUM VPW nch L=4e-08 W=2.2e-07 
M15 CO 9 VSS VPW nch L=4e-08 W=2.2e-07 
M16 VSS 9 CO VPW nch L=4e-08 W=2.2e-07 
M17 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M19 5 B 1 VNW pch L=4e-08 W=3.8e-07 
M20 4 7 5 VNW pch L=4e-08 W=3.8e-07 
M21 6 7 1 VNW pch L=4e-08 W=3.8e-07 
M22 4 B 6 VNW pch L=4e-08 W=3.8e-07 
M23 7 B VDD VNW pch L=4e-08 W=3.8e-07 
M24 9 5 7 VNW pch L=4e-08 W=3.8e-07 
M25 8 6 9 VNW pch L=4e-08 W=3.8e-07 
M26 11 6 10 VNW pch L=4e-08 W=3.8e-07 
M27 8 5 11 VNW pch L=4e-08 W=3.8e-07 
M28 VDD 10 8 VNW pch L=4e-08 W=3.8e-07 
M29 10 CIN VDD VNW pch L=4e-08 W=3.8e-07 
M30 SUM 11 VDD VNW pch L=4e-08 W=2.85e-07 
M31 VDD 11 SUM VNW pch L=4e-08 W=2.85e-07 
M32 CO 9 VDD VNW pch L=4e-08 W=2.85e-07 
M33 VDD 9 CO VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT ADDFCIN_X2M_A9TR CO SUM VDD VNW VPW VSS A B CIN
M0 VSS 4 1 VPW nch L=4e-08 W=3.15e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.15e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.15e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.15e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.15e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.15e-07 
M6 7 B VSS VPW nch L=4e-08 W=2.3e-07 
M7 9 5 8 VPW nch L=4e-08 W=2.3e-07 
M8 7 6 9 VPW nch L=4e-08 W=2.3e-07 
M9 11 6 8 VPW nch L=4e-08 W=2.3e-07 
M10 10 5 11 VPW nch L=4e-08 W=2.3e-07 
M11 VSS 10 8 VPW nch L=4e-08 W=2.3e-07 
M12 10 CIN VSS VPW nch L=4e-08 W=2.3e-07 
M13 SUM 11 VSS VPW nch L=4e-08 W=2.95e-07 
M14 VSS 11 SUM VPW nch L=4e-08 W=2.95e-07 
M15 CO 9 VSS VPW nch L=4e-08 W=2.95e-07 
M16 VSS 9 CO VPW nch L=4e-08 W=2.95e-07 
M17 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M19 5 B 1 VNW pch L=4e-08 W=3.8e-07 
M20 4 7 5 VNW pch L=4e-08 W=3.8e-07 
M21 6 7 1 VNW pch L=4e-08 W=3.8e-07 
M22 4 B 6 VNW pch L=4e-08 W=3.8e-07 
M23 7 B VDD VNW pch L=4e-08 W=3.8e-07 
M24 9 5 7 VNW pch L=4e-08 W=3.8e-07 
M25 8 6 9 VNW pch L=4e-08 W=3.8e-07 
M26 11 6 10 VNW pch L=4e-08 W=3.8e-07 
M27 8 5 11 VNW pch L=4e-08 W=3.8e-07 
M28 VDD 10 8 VNW pch L=4e-08 W=3.8e-07 
M29 10 CIN VDD VNW pch L=4e-08 W=3.8e-07 
M30 SUM 11 VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD 11 SUM VNW pch L=4e-08 W=3.8e-07 
M32 CO 9 VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD 9 CO VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT ADDFH_X1M_A9TR CO SUM VDD VNW VPW VSS A B CI
M0 VSS 4 1 VPW nch L=4e-08 W=3.15e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.15e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.15e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.15e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.15e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.15e-07 
M6 7 B VSS VPW nch L=4e-08 W=1.55e-07 
M7 9 5 8 VPW nch L=4e-08 W=1.55e-07 
M8 7 6 9 VPW nch L=4e-08 W=1.55e-07 
M9 11 6 8 VPW nch L=4e-08 W=1.55e-07 
M10 10 5 11 VPW nch L=4e-08 W=1.55e-07 
M11 VSS 8 10 VPW nch L=4e-08 W=1.55e-07 
M12 8 CI VSS VPW nch L=4e-08 W=1.55e-07 
M13 VSS 11 SUM VPW nch L=4e-08 W=2.95e-07 
M14 CO 9 VSS VPW nch L=4e-08 W=2.95e-07 
M15 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M16 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M17 5 B 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 7 5 VNW pch L=4e-08 W=3.8e-07 
M19 6 7 1 VNW pch L=4e-08 W=3.8e-07 
M20 4 B 6 VNW pch L=4e-08 W=3.8e-07 
M21 7 B VDD VNW pch L=4e-08 W=2.6e-07 
M22 9 5 7 VNW pch L=4e-08 W=2.6e-07 
M23 8 6 9 VNW pch L=4e-08 W=2.6e-07 
M24 11 6 10 VNW pch L=4e-08 W=2.6e-07 
M25 8 5 11 VNW pch L=4e-08 W=2.6e-07 
M26 VDD 8 10 VNW pch L=4e-08 W=2.6e-07 
M27 8 CI VDD VNW pch L=4e-08 W=2.6e-07 
M28 VDD 11 SUM VNW pch L=4e-08 W=3.8e-07 
M29 CO 9 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT ADDFH_X1P4M_A9TR CO SUM VDD VNW VPW VSS A B CI
M0 VSS 4 1 VPW nch L=4e-08 W=3.15e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.15e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.15e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.15e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.15e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.15e-07 
M6 7 B VSS VPW nch L=4e-08 W=2.3e-07 
M7 9 5 8 VPW nch L=4e-08 W=2.3e-07 
M8 7 6 9 VPW nch L=4e-08 W=2.3e-07 
M9 11 6 8 VPW nch L=4e-08 W=2.3e-07 
M10 10 5 11 VPW nch L=4e-08 W=2.3e-07 
M11 VSS 8 10 VPW nch L=4e-08 W=2.3e-07 
M12 8 CI VSS VPW nch L=4e-08 W=2.3e-07 
M13 SUM 11 VSS VPW nch L=4e-08 W=2.2e-07 
M14 VSS 11 SUM VPW nch L=4e-08 W=2.2e-07 
M15 CO 9 VSS VPW nch L=4e-08 W=2.2e-07 
M16 VSS 9 CO VPW nch L=4e-08 W=2.2e-07 
M17 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M19 5 B 1 VNW pch L=4e-08 W=3.8e-07 
M20 4 7 5 VNW pch L=4e-08 W=3.8e-07 
M21 6 7 1 VNW pch L=4e-08 W=3.8e-07 
M22 4 B 6 VNW pch L=4e-08 W=3.8e-07 
M23 7 B VDD VNW pch L=4e-08 W=3.8e-07 
M24 9 5 7 VNW pch L=4e-08 W=3.8e-07 
M25 8 6 9 VNW pch L=4e-08 W=3.8e-07 
M26 11 6 10 VNW pch L=4e-08 W=3.8e-07 
M27 8 5 11 VNW pch L=4e-08 W=3.8e-07 
M28 VDD 8 10 VNW pch L=4e-08 W=3.8e-07 
M29 8 CI VDD VNW pch L=4e-08 W=3.8e-07 
M30 SUM 11 VDD VNW pch L=4e-08 W=2.85e-07 
M31 VDD 11 SUM VNW pch L=4e-08 W=2.85e-07 
M32 CO 9 VDD VNW pch L=4e-08 W=2.85e-07 
M33 VDD 9 CO VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT ADDFH_X2M_A9TR CO SUM VDD VNW VPW VSS A B CI
M0 VSS 4 1 VPW nch L=4e-08 W=3.15e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.15e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.15e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.15e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.15e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.15e-07 
M6 7 B VSS VPW nch L=4e-08 W=2.3e-07 
M7 9 5 8 VPW nch L=4e-08 W=2.3e-07 
M8 7 6 9 VPW nch L=4e-08 W=2.3e-07 
M9 11 6 8 VPW nch L=4e-08 W=2.3e-07 
M10 10 5 11 VPW nch L=4e-08 W=2.3e-07 
M11 VSS 8 10 VPW nch L=4e-08 W=2.3e-07 
M12 8 CI VSS VPW nch L=4e-08 W=2.3e-07 
M13 SUM 11 VSS VPW nch L=4e-08 W=2.95e-07 
M14 VSS 11 SUM VPW nch L=4e-08 W=2.95e-07 
M15 CO 9 VSS VPW nch L=4e-08 W=2.95e-07 
M16 VSS 9 CO VPW nch L=4e-08 W=2.95e-07 
M17 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M19 5 B 1 VNW pch L=4e-08 W=3.8e-07 
M20 4 7 5 VNW pch L=4e-08 W=3.8e-07 
M21 6 7 1 VNW pch L=4e-08 W=3.8e-07 
M22 4 B 6 VNW pch L=4e-08 W=3.8e-07 
M23 7 B VDD VNW pch L=4e-08 W=3.8e-07 
M24 9 5 7 VNW pch L=4e-08 W=3.8e-07 
M25 8 6 9 VNW pch L=4e-08 W=3.8e-07 
M26 11 6 10 VNW pch L=4e-08 W=3.8e-07 
M27 8 5 11 VNW pch L=4e-08 W=3.8e-07 
M28 VDD 8 10 VNW pch L=4e-08 W=3.8e-07 
M29 8 CI VDD VNW pch L=4e-08 W=3.8e-07 
M30 SUM 11 VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD 11 SUM VNW pch L=4e-08 W=3.8e-07 
M32 CO 9 VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD 9 CO VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT ADDF_X1M_A9TR CO S VDD VNW VPW VSS A B CI
M0 VSS 6 CO VPW nch L=4e-08 W=3.1e-07 
M1 4 A VSS VPW nch L=4e-08 W=2.2e-07 
M2 VSS B 4 VPW nch L=4e-08 W=2.2e-07 
M3 17 B VSS VPW nch L=4e-08 W=2.2e-07 
M4 6 A 17 VPW nch L=4e-08 W=2.2e-07 
M5 4 CI 6 VPW nch L=4e-08 W=2.2e-07 
M6 7 CI VSS VPW nch L=4e-08 W=3.5e-07 
M7 VSS A 7 VPW nch L=4e-08 W=3.5e-07 
M8 7 B VSS VPW nch L=4e-08 W=3.5e-07 
M9 9 6 7 VPW nch L=4e-08 W=3.5e-07 
M10 18 CI 9 VPW nch L=4e-08 W=2e-07 
M11 19 A 18 VPW nch L=4e-08 W=2e-07 
M12 VSS B 19 VPW nch L=4e-08 W=2e-07 
M13 S 9 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VDD 6 CO VNW pch L=4e-08 W=4e-07 
M15 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M16 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M17 14 B VDD VNW pch L=4e-08 W=3.8e-07 
M18 6 A 14 VNW pch L=4e-08 W=3.8e-07 
M19 5 CI 6 VNW pch L=4e-08 W=3.8e-07 
M20 8 CI VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD A 8 VNW pch L=4e-08 W=3.8e-07 
M22 8 B VDD VNW pch L=4e-08 W=3.8e-07 
M23 9 6 8 VNW pch L=4e-08 W=3.8e-07 
M24 15 CI 9 VNW pch L=4e-08 W=3.8e-07 
M25 16 A 15 VNW pch L=4e-08 W=3.8e-07 
M26 VDD B 16 VNW pch L=4e-08 W=3.8e-07 
M27 S 9 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT ADDF_X1P4M_A9TR CO S VDD VNW VPW VSS A B CI
M0 CO 6 VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS 6 CO VPW nch L=4e-08 W=2.2e-07 
M2 4 A VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS B 4 VPW nch L=4e-08 W=2.2e-07 
M4 17 B VSS VPW nch L=4e-08 W=2.2e-07 
M5 6 A 17 VPW nch L=4e-08 W=2.2e-07 
M6 4 CI 6 VPW nch L=4e-08 W=2.2e-07 
M7 7 CI VSS VPW nch L=4e-08 W=3.5e-07 
M8 VSS A 7 VPW nch L=4e-08 W=3.5e-07 
M9 7 B VSS VPW nch L=4e-08 W=3.5e-07 
M10 9 6 7 VPW nch L=4e-08 W=3.5e-07 
M11 18 CI 9 VPW nch L=4e-08 W=2e-07 
M12 19 A 18 VPW nch L=4e-08 W=2e-07 
M13 VSS B 19 VPW nch L=4e-08 W=2e-07 
M14 S 9 VSS VPW nch L=4e-08 W=2.2e-07 
M15 VSS 9 S VPW nch L=4e-08 W=2.2e-07 
M16 CO 6 VDD VNW pch L=4e-08 W=2.85e-07 
M17 VDD 6 CO VNW pch L=4e-08 W=2.85e-07 
M18 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M19 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M20 14 B VDD VNW pch L=4e-08 W=3.8e-07 
M21 6 A 14 VNW pch L=4e-08 W=3.8e-07 
M22 5 CI 6 VNW pch L=4e-08 W=3.8e-07 
M23 8 CI VDD VNW pch L=4e-08 W=3.8e-07 
M24 VDD A 8 VNW pch L=4e-08 W=3.8e-07 
M25 8 B VDD VNW pch L=4e-08 W=3.8e-07 
M26 9 6 8 VNW pch L=4e-08 W=3.8e-07 
M27 15 CI 9 VNW pch L=4e-08 W=3.8e-07 
M28 16 A 15 VNW pch L=4e-08 W=3.8e-07 
M29 VDD B 16 VNW pch L=4e-08 W=3.8e-07 
M30 S 9 VDD VNW pch L=4e-08 W=2.85e-07 
M31 VDD 9 S VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT ADDF_X2M_A9TR CO S VDD VNW VPW VSS A B CI
M0 CO 6 VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS 6 CO VPW nch L=4e-08 W=3.1e-07 
M2 4 A VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS B 4 VPW nch L=4e-08 W=2.2e-07 
M4 17 B VSS VPW nch L=4e-08 W=2.2e-07 
M5 6 A 17 VPW nch L=4e-08 W=2.2e-07 
M6 4 CI 6 VPW nch L=4e-08 W=2.2e-07 
M7 7 CI VSS VPW nch L=4e-08 W=3.5e-07 
M8 VSS A 7 VPW nch L=4e-08 W=3.5e-07 
M9 7 B VSS VPW nch L=4e-08 W=3.5e-07 
M10 9 6 7 VPW nch L=4e-08 W=3.5e-07 
M11 18 CI 9 VPW nch L=4e-08 W=2e-07 
M12 19 A 18 VPW nch L=4e-08 W=2e-07 
M13 VSS B 19 VPW nch L=4e-08 W=2e-07 
M14 S 9 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 9 S VPW nch L=4e-08 W=3.1e-07 
M16 CO 6 VDD VNW pch L=4e-08 W=4e-07 
M17 VDD 6 CO VNW pch L=4e-08 W=4e-07 
M18 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M19 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M20 14 B VDD VNW pch L=4e-08 W=3.8e-07 
M21 6 A 14 VNW pch L=4e-08 W=3.8e-07 
M22 5 CI 6 VNW pch L=4e-08 W=3.8e-07 
M23 8 CI VDD VNW pch L=4e-08 W=3.8e-07 
M24 VDD A 8 VNW pch L=4e-08 W=3.8e-07 
M25 8 B VDD VNW pch L=4e-08 W=3.8e-07 
M26 9 6 8 VNW pch L=4e-08 W=3.8e-07 
M27 15 CI 9 VNW pch L=4e-08 W=3.8e-07 
M28 16 A 15 VNW pch L=4e-08 W=3.8e-07 
M29 VDD B 16 VNW pch L=4e-08 W=3.8e-07 
M30 S 9 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 9 S VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT ADDH_X1M_A9TR CO S VDD VNW VPW VSS A B
M0 VSS 4 CO VPW nch L=4e-08 W=3.1e-07 
M1 11 B VSS VPW nch L=4e-08 W=3.2e-07 
M2 4 A 11 VPW nch L=4e-08 W=3.2e-07 
M3 VSS B 5 VPW nch L=4e-08 W=2.35e-07 
M4 5 A VSS VPW nch L=4e-08 W=2.35e-07 
M5 6 4 5 VPW nch L=4e-08 W=2.35e-07 
M6 S 6 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VDD 4 CO VNW pch L=4e-08 W=4e-07 
M8 4 B VDD VNW pch L=4e-08 W=2.8e-07 
M9 VDD A 4 VNW pch L=4e-08 W=2.8e-07 
M10 10 B VDD VNW pch L=4e-08 W=2.8e-07 
M11 6 A 10 VNW pch L=4e-08 W=2.8e-07 
M12 VDD 4 6 VNW pch L=4e-08 W=1.3e-07 
M13 S 6 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT ADDH_X1P4M_A9TR CO S VDD VNW VPW VSS A B
M0 CO 4 VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS 4 CO VPW nch L=4e-08 W=2.2e-07 
M2 11 B VSS VPW nch L=4e-08 W=4e-07 
M3 4 A 11 VPW nch L=4e-08 W=4e-07 
M4 VSS B 5 VPW nch L=4e-08 W=3.35e-07 
M5 5 A VSS VPW nch L=4e-08 W=3.35e-07 
M6 6 4 5 VPW nch L=4e-08 W=3.35e-07 
M7 S 6 VSS VPW nch L=4e-08 W=2.2e-07 
M8 VSS 6 S VPW nch L=4e-08 W=2.2e-07 
M9 CO 4 VDD VNW pch L=4e-08 W=2.85e-07 
M10 VDD 4 CO VNW pch L=4e-08 W=2.85e-07 
M11 4 B VDD VNW pch L=4e-08 W=3.45e-07 
M12 VDD A 4 VNW pch L=4e-08 W=3.45e-07 
M13 10 B VDD VNW pch L=4e-08 W=3.45e-07 
M14 6 A 10 VNW pch L=4e-08 W=3.45e-07 
M15 VDD 4 6 VNW pch L=4e-08 W=1.85e-07 
M16 S 6 VDD VNW pch L=4e-08 W=2.85e-07 
M17 VDD 6 S VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT ADDH_X2M_A9TR CO S VDD VNW VPW VSS A B
M0 CO 4 VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS 4 CO VPW nch L=4e-08 W=3.1e-07 
M2 11 B VSS VPW nch L=4e-08 W=4e-07 
M3 4 A 11 VPW nch L=4e-08 W=4e-07 
M4 VSS B 5 VPW nch L=4e-08 W=4e-07 
M5 5 A VSS VPW nch L=4e-08 W=4e-07 
M6 6 4 5 VPW nch L=4e-08 W=4e-07 
M7 S 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 6 S VPW nch L=4e-08 W=3.1e-07 
M9 CO 4 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD 4 CO VNW pch L=4e-08 W=4e-07 
M11 4 B VDD VNW pch L=4e-08 W=3.45e-07 
M12 VDD A 4 VNW pch L=4e-08 W=3.45e-07 
M13 10 B VDD VNW pch L=4e-08 W=3.8e-07 
M14 6 A 10 VNW pch L=4e-08 W=3.8e-07 
M15 VDD 4 6 VNW pch L=4e-08 W=2.2e-07 
M16 S 6 VDD VNW pch L=4e-08 W=4e-07 
M17 VDD 6 S VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X0P5B_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS B 7 VPW nch L=4e-08 W=1.2e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M3 1 A VDD VNW pch L=4e-08 W=1.4e-07 
M4 VDD B 1 VNW pch L=4e-08 W=1.4e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT AND2_X0P5M_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=1.4e-07 
M1 VSS B 7 VPW nch L=4e-08 W=1.4e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=1.55e-07 
M3 1 A VDD VNW pch L=4e-08 W=1.2e-07 
M4 VDD B 1 VNW pch L=4e-08 W=1.2e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AND2_X0P7B_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=1.25e-07 
M1 VSS B 7 VPW nch L=4e-08 W=1.25e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M3 1 A VDD VNW pch L=4e-08 W=1.45e-07 
M4 VDD B 1 VNW pch L=4e-08 W=1.45e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AND2_X0P7M_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=1.4e-07 
M1 VSS B 7 VPW nch L=4e-08 W=1.4e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M3 1 A VDD VNW pch L=4e-08 W=1.2e-07 
M4 VDD B 1 VNW pch L=4e-08 W=1.2e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AND2_X11B_A9TR Y VDD VNW VPW VSS A B
M0 7 B VSS VPW nch L=4e-08 W=3.45e-07 
M1 3 A 7 VPW nch L=4e-08 W=3.45e-07 
M2 8 A 3 VPW nch L=4e-08 W=3.45e-07 
M3 VSS B 8 VPW nch L=4e-08 W=3.45e-07 
M4 9 B VSS VPW nch L=4e-08 W=3.45e-07 
M5 3 A 9 VPW nch L=4e-08 W=3.45e-07 
M6 10 A 3 VPW nch L=4e-08 W=3.45e-07 
M7 VSS B 10 VPW nch L=4e-08 W=3.45e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=3.55e-07 
M9 VSS 3 Y VPW nch L=4e-08 W=3.55e-07 
M10 Y 3 VSS VPW nch L=4e-08 W=3.55e-07 
M11 VSS 3 Y VPW nch L=4e-08 W=3.55e-07 
M12 Y 3 VSS VPW nch L=4e-08 W=3.55e-07 
M13 VSS 3 Y VPW nch L=4e-08 W=3.55e-07 
M14 Y 3 VSS VPW nch L=4e-08 W=3.55e-07 
M15 3 B VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A 3 VNW pch L=4e-08 W=4e-07 
M17 3 A VDD VNW pch L=4e-08 W=4e-07 
M18 VDD B 3 VNW pch L=4e-08 W=4e-07 
M19 3 B VDD VNW pch L=4e-08 W=4e-07 
M20 VDD A 3 VNW pch L=4e-08 W=4e-07 
M21 3 A VDD VNW pch L=4e-08 W=4e-07 
M22 VDD B 3 VNW pch L=4e-08 W=4e-07 
M23 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M25 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M27 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M29 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M31 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M33 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X11M_A9TR Y VDD VNW VPW VSS A B
M0 8 A 1 VPW nch L=4e-08 W=3.5e-07 
M1 VSS B 8 VPW nch L=4e-08 W=3.5e-07 
M2 9 B VSS VPW nch L=4e-08 W=3.5e-07 
M3 1 A 9 VPW nch L=4e-08 W=3.5e-07 
M4 10 A 1 VPW nch L=4e-08 W=3.5e-07 
M5 VSS B 10 VPW nch L=4e-08 W=3.5e-07 
M6 11 B VSS VPW nch L=4e-08 W=3.5e-07 
M7 1 A 11 VPW nch L=4e-08 W=3.5e-07 
M8 12 A 1 VPW nch L=4e-08 W=3.5e-07 
M9 VSS B 12 VPW nch L=4e-08 W=3.5e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M16 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M18 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M20 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M21 1 B VDD VNW pch L=4e-08 W=3.75e-07 
M22 VDD A 1 VNW pch L=4e-08 W=3.75e-07 
M23 1 A VDD VNW pch L=4e-08 W=3.75e-07 
M24 VDD B 1 VNW pch L=4e-08 W=3.75e-07 
M25 1 B VDD VNW pch L=4e-08 W=3.75e-07 
M26 VDD A 1 VNW pch L=4e-08 W=3.75e-07 
M27 1 A VDD VNW pch L=4e-08 W=3.75e-07 
M28 VDD B 1 VNW pch L=4e-08 W=3.75e-07 
M29 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M31 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M33 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M35 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M37 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M39 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X1B_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=1.5e-07 
M1 VSS B 7 VPW nch L=4e-08 W=1.5e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M3 1 A VDD VNW pch L=4e-08 W=1.75e-07 
M4 VDD B 1 VNW pch L=4e-08 W=1.75e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X1M_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=1.75e-07 
M1 VSS B 7 VPW nch L=4e-08 W=1.75e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M3 1 A VDD VNW pch L=4e-08 W=1.5e-07 
M4 VDD B 1 VNW pch L=4e-08 W=1.5e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X1P4B_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=1.9e-07 
M1 VSS B 7 VPW nch L=4e-08 W=1.9e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M4 1 A VDD VNW pch L=4e-08 W=2.2e-07 
M5 VDD B 1 VNW pch L=4e-08 W=2.2e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AND2_X1P4M_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=2.35e-07 
M1 VSS B 7 VPW nch L=4e-08 W=2.35e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=2.2e-07 
M4 1 A VDD VNW pch L=4e-08 W=2e-07 
M5 VDD B 1 VNW pch L=4e-08 W=2e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AND2_X2B_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=2.5e-07 
M1 VSS B 7 VPW nch L=4e-08 W=2.5e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M4 1 A VDD VNW pch L=4e-08 W=2.9e-07 
M5 VDD B 1 VNW pch L=4e-08 W=2.9e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X2M_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=3.1e-07 
M1 VSS B 7 VPW nch L=4e-08 W=3.1e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M4 1 A VDD VNW pch L=4e-08 W=2.7e-07 
M5 VDD B 1 VNW pch L=4e-08 W=2.7e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X3B_A9TR Y VDD VNW VPW VSS A B
M0 7 B VSS VPW nch L=4e-08 W=2.05e-07 
M1 3 A 7 VPW nch L=4e-08 W=2.05e-07 
M2 8 A 3 VPW nch L=4e-08 W=2.05e-07 
M3 VSS B 8 VPW nch L=4e-08 W=2.05e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.4e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.4e-07 
M6 3 B VDD VNW pch L=4e-08 W=2.35e-07 
M7 VDD A 3 VNW pch L=4e-08 W=2.35e-07 
M8 3 A VDD VNW pch L=4e-08 W=2.35e-07 
M9 VDD B 3 VNW pch L=4e-08 W=2.35e-07 
M10 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M12 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X3M_A9TR Y VDD VNW VPW VSS A B
M0 7 B VSS VPW nch L=4e-08 W=2.45e-07 
M1 3 A 7 VPW nch L=4e-08 W=2.45e-07 
M2 8 A 3 VPW nch L=4e-08 W=2.45e-07 
M3 VSS B 8 VPW nch L=4e-08 W=2.45e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M7 3 B VDD VNW pch L=4e-08 W=2.1e-07 
M8 VDD A 3 VNW pch L=4e-08 W=2.1e-07 
M9 3 A VDD VNW pch L=4e-08 W=2.1e-07 
M10 VDD B 3 VNW pch L=4e-08 W=2.1e-07 
M11 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M13 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X4B_A9TR Y VDD VNW VPW VSS A B
M0 7 B VSS VPW nch L=4e-08 W=2.55e-07 
M1 3 A 7 VPW nch L=4e-08 W=2.55e-07 
M2 8 A 3 VPW nch L=4e-08 W=2.55e-07 
M3 VSS B 8 VPW nch L=4e-08 W=2.55e-07 
M4 VSS 3 Y VPW nch L=4e-08 W=3e-07 
M5 Y 3 VSS VPW nch L=4e-08 W=3e-07 
M6 VSS 3 Y VPW nch L=4e-08 W=3e-07 
M7 3 B VDD VNW pch L=4e-08 W=2.95e-07 
M8 VDD A 3 VNW pch L=4e-08 W=2.95e-07 
M9 3 A VDD VNW pch L=4e-08 W=2.95e-07 
M10 VDD B 3 VNW pch L=4e-08 W=2.95e-07 
M11 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M13 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X4M_A9TR Y VDD VNW VPW VSS A B
M0 7 B VSS VPW nch L=4e-08 W=3.15e-07 
M1 3 A 7 VPW nch L=4e-08 W=3.15e-07 
M2 8 A 3 VPW nch L=4e-08 W=3.15e-07 
M3 VSS B 8 VPW nch L=4e-08 W=3.15e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M8 3 B VDD VNW pch L=4e-08 W=2.7e-07 
M9 VDD A 3 VNW pch L=4e-08 W=2.7e-07 
M10 3 A VDD VNW pch L=4e-08 W=2.7e-07 
M11 VDD B 3 VNW pch L=4e-08 W=2.7e-07 
M12 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M13 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X6B_A9TR Y VDD VNW VPW VSS A B
M0 8 B VSS VPW nch L=4e-08 W=3.9e-07 
M1 2 A 8 VPW nch L=4e-08 W=3.9e-07 
M2 9 A 2 VPW nch L=4e-08 W=3.9e-07 
M3 VSS B 9 VPW nch L=4e-08 W=3.9e-07 
M4 Y 2 VSS VPW nch L=4e-08 W=3.35e-07 
M5 VSS 2 Y VPW nch L=4e-08 W=3.35e-07 
M6 Y 2 VSS VPW nch L=4e-08 W=3.35e-07 
M7 VSS 2 Y VPW nch L=4e-08 W=3.35e-07 
M8 2 A VDD VNW pch L=4e-08 W=3e-07 
M9 VDD B 2 VNW pch L=4e-08 W=3e-07 
M10 2 B VDD VNW pch L=4e-08 W=3e-07 
M11 VDD A 2 VNW pch L=4e-08 W=3e-07 
M12 2 A VDD VNW pch L=4e-08 W=3e-07 
M13 VDD B 2 VNW pch L=4e-08 W=3e-07 
M14 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M16 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M17 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M18 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 2 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X6M_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=3.2e-07 
M1 VSS B 7 VPW nch L=4e-08 W=3.2e-07 
M2 8 B VSS VPW nch L=4e-08 W=3.2e-07 
M3 1 A 8 VPW nch L=4e-08 W=3.2e-07 
M4 9 A 1 VPW nch L=4e-08 W=3.2e-07 
M5 VSS B 9 VPW nch L=4e-08 W=3.2e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M12 1 A VDD VNW pch L=4e-08 W=2.75e-07 
M13 VDD B 1 VNW pch L=4e-08 W=2.75e-07 
M14 1 B VDD VNW pch L=4e-08 W=2.75e-07 
M15 VDD A 1 VNW pch L=4e-08 W=2.75e-07 
M16 1 A VDD VNW pch L=4e-08 W=2.75e-07 
M17 VDD B 1 VNW pch L=4e-08 W=2.75e-07 
M18 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M20 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X8B_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=3.3e-07 
M1 VSS B 7 VPW nch L=4e-08 W=3.3e-07 
M2 8 B VSS VPW nch L=4e-08 W=3.3e-07 
M3 1 A 8 VPW nch L=4e-08 W=3.3e-07 
M4 9 A 1 VPW nch L=4e-08 W=3.3e-07 
M5 VSS B 9 VPW nch L=4e-08 W=3.3e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=3.6e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=3.6e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=3.6e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=3.6e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=3.6e-07 
M11 1 A VDD VNW pch L=4e-08 W=3.8e-07 
M12 VDD B 1 VNW pch L=4e-08 W=3.8e-07 
M13 1 B VDD VNW pch L=4e-08 W=3.8e-07 
M14 VDD A 1 VNW pch L=4e-08 W=3.8e-07 
M15 1 A VDD VNW pch L=4e-08 W=3.8e-07 
M16 VDD B 1 VNW pch L=4e-08 W=3.8e-07 
M17 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M19 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M21 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M23 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND2_X8M_A9TR Y VDD VNW VPW VSS A B
M0 7 A 1 VPW nch L=4e-08 W=4e-07 
M1 VSS B 7 VPW nch L=4e-08 W=4e-07 
M2 8 B VSS VPW nch L=4e-08 W=4e-07 
M3 1 A 8 VPW nch L=4e-08 W=4e-07 
M4 9 A 1 VPW nch L=4e-08 W=4e-07 
M5 VSS B 9 VPW nch L=4e-08 W=4e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M14 1 A VDD VNW pch L=4e-08 W=3.45e-07 
M15 VDD B 1 VNW pch L=4e-08 W=3.45e-07 
M16 1 B VDD VNW pch L=4e-08 W=3.45e-07 
M17 VDD A 1 VNW pch L=4e-08 W=3.45e-07 
M18 1 A VDD VNW pch L=4e-08 W=3.45e-07 
M19 VDD B 1 VNW pch L=4e-08 W=3.45e-07 
M20 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M24 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M26 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND3_X0P5M_A9TR Y VDD VNW VPW VSS A B C
M0 8 A 1 VPW nch L=4e-08 W=1.8e-07 
M1 9 B 8 VPW nch L=4e-08 W=1.8e-07 
M2 VSS C 9 VPW nch L=4e-08 W=1.8e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=1.55e-07 
M4 VDD A 1 VNW pch L=4e-08 W=1.2e-07 
M5 1 B VDD VNW pch L=4e-08 W=1.2e-07 
M6 VDD C 1 VNW pch L=4e-08 W=1.2e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AND3_X0P7M_A9TR Y VDD VNW VPW VSS A B C
M0 8 A 1 VPW nch L=4e-08 W=2.25e-07 
M1 9 B 8 VPW nch L=4e-08 W=2.25e-07 
M2 VSS C 9 VPW nch L=4e-08 W=2.25e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M4 VDD A 1 VNW pch L=4e-08 W=1.5e-07 
M5 1 B VDD VNW pch L=4e-08 W=1.5e-07 
M6 VDD C 1 VNW pch L=4e-08 W=1.5e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AND3_X11M_A9TR Y VDD VNW VPW VSS A B C
M0 9 A 1 VPW nch L=4e-08 W=4e-07 
M1 3 B 9 VPW nch L=4e-08 W=4e-07 
M2 10 B 3 VPW nch L=4e-08 W=4e-07 
M3 1 A 10 VPW nch L=4e-08 W=4e-07 
M4 11 A 1 VPW nch L=4e-08 W=4e-07 
M5 3 B 11 VPW nch L=4e-08 W=4e-07 
M6 12 B 3 VPW nch L=4e-08 W=4e-07 
M7 1 A 12 VPW nch L=4e-08 W=4e-07 
M8 13 A 1 VPW nch L=4e-08 W=4e-07 
M9 3 B 13 VPW nch L=4e-08 W=4e-07 
M10 14 B 3 VPW nch L=4e-08 W=4e-07 
M11 1 A 14 VPW nch L=4e-08 W=4e-07 
M12 15 A 1 VPW nch L=4e-08 W=4e-07 
M13 3 B 15 VPW nch L=4e-08 W=4e-07 
M14 VSS C 3 VPW nch L=4e-08 W=4e-07 
M15 3 C VSS VPW nch L=4e-08 W=4e-07 
M16 VSS C 3 VPW nch L=4e-08 W=4e-07 
M17 3 C VSS VPW nch L=4e-08 W=4e-07 
M18 VSS C 3 VPW nch L=4e-08 W=4e-07 
M19 3 C VSS VPW nch L=4e-08 W=4e-07 
M20 VSS C 3 VPW nch L=4e-08 W=4e-07 
M21 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M22 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M23 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M24 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M25 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M26 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M27 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M28 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M29 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M30 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M31 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M32 VDD A 1 VNW pch L=4e-08 W=2.7e-07 
M33 1 B VDD VNW pch L=4e-08 W=2.7e-07 
M34 VDD B 1 VNW pch L=4e-08 W=2.7e-07 
M35 1 A VDD VNW pch L=4e-08 W=2.7e-07 
M36 VDD A 1 VNW pch L=4e-08 W=2.7e-07 
M37 1 B VDD VNW pch L=4e-08 W=2.7e-07 
M38 VDD B 1 VNW pch L=4e-08 W=2.7e-07 
M39 1 A VDD VNW pch L=4e-08 W=2.7e-07 
M40 VDD A 1 VNW pch L=4e-08 W=2.7e-07 
M41 1 B VDD VNW pch L=4e-08 W=2.7e-07 
M42 VDD B 1 VNW pch L=4e-08 W=2.7e-07 
M43 1 A VDD VNW pch L=4e-08 W=2.7e-07 
M44 VDD A 1 VNW pch L=4e-08 W=2.7e-07 
M45 1 B VDD VNW pch L=4e-08 W=2.7e-07 
M46 VDD C 1 VNW pch L=4e-08 W=2.7e-07 
M47 1 C VDD VNW pch L=4e-08 W=2.7e-07 
M48 VDD C 1 VNW pch L=4e-08 W=2.7e-07 
M49 1 C VDD VNW pch L=4e-08 W=2.7e-07 
M50 VDD C 1 VNW pch L=4e-08 W=2.7e-07 
M51 1 C VDD VNW pch L=4e-08 W=2.7e-07 
M52 VDD C 1 VNW pch L=4e-08 W=2.7e-07 
M53 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M54 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M55 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M56 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M57 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M58 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M59 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M60 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M61 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M62 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M63 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND3_X1M_A9TR Y VDD VNW VPW VSS A B C
M0 8 A 1 VPW nch L=4e-08 W=2.8e-07 
M1 9 B 8 VPW nch L=4e-08 W=2.8e-07 
M2 VSS C 9 VPW nch L=4e-08 W=2.8e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VDD A 1 VNW pch L=4e-08 W=1.85e-07 
M5 1 B VDD VNW pch L=4e-08 W=1.85e-07 
M6 VDD C 1 VNW pch L=4e-08 W=1.85e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND3_X1P4M_A9TR Y VDD VNW VPW VSS A B C
M0 8 A 1 VPW nch L=4e-08 W=3.75e-07 
M1 9 B 8 VPW nch L=4e-08 W=3.75e-07 
M2 VSS C 9 VPW nch L=4e-08 W=3.75e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=2.2e-07 
M5 VDD A 1 VNW pch L=4e-08 W=2.5e-07 
M6 1 B VDD VNW pch L=4e-08 W=2.5e-07 
M7 VDD C 1 VNW pch L=4e-08 W=2.5e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AND3_X2M_A9TR Y VDD VNW VPW VSS A B C
M0 8 C VSS VPW nch L=4e-08 W=2.65e-07 
M1 9 B 8 VPW nch L=4e-08 W=2.65e-07 
M2 3 A 9 VPW nch L=4e-08 W=2.65e-07 
M3 10 A 3 VPW nch L=4e-08 W=2.65e-07 
M4 11 B 10 VPW nch L=4e-08 W=2.65e-07 
M5 VSS C 11 VPW nch L=4e-08 W=2.65e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M8 3 C VDD VNW pch L=4e-08 W=1.75e-07 
M9 VDD B 3 VNW pch L=4e-08 W=1.75e-07 
M10 3 A VDD VNW pch L=4e-08 W=1.75e-07 
M11 VDD A 3 VNW pch L=4e-08 W=1.75e-07 
M12 3 B VDD VNW pch L=4e-08 W=1.75e-07 
M13 VDD C 3 VNW pch L=4e-08 W=1.75e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND3_X3M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=3.7e-07 
M1 1 C VSS VPW nch L=4e-08 W=3.7e-07 
M2 9 B 1 VPW nch L=4e-08 W=3.7e-07 
M3 4 A 9 VPW nch L=4e-08 W=3.7e-07 
M4 10 A 4 VPW nch L=4e-08 W=3.7e-07 
M5 1 B 10 VPW nch L=4e-08 W=3.7e-07 
M6 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M8 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M9 4 C VDD VNW pch L=4e-08 W=2.45e-07 
M10 VDD C 4 VNW pch L=4e-08 W=2.45e-07 
M11 4 B VDD VNW pch L=4e-08 W=2.45e-07 
M12 VDD A 4 VNW pch L=4e-08 W=2.45e-07 
M13 4 A VDD VNW pch L=4e-08 W=2.45e-07 
M14 VDD B 4 VNW pch L=4e-08 W=2.45e-07 
M15 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M17 Y 4 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND3_X4M_A9TR Y VDD VNW VPW VSS A B C
M0 9 A 1 VPW nch L=4e-08 W=3.3e-07 
M1 3 B 9 VPW nch L=4e-08 W=3.3e-07 
M2 10 B 3 VPW nch L=4e-08 W=3.3e-07 
M3 1 A 10 VPW nch L=4e-08 W=3.3e-07 
M4 11 A 1 VPW nch L=4e-08 W=3.3e-07 
M5 3 B 11 VPW nch L=4e-08 W=3.3e-07 
M6 VSS C 3 VPW nch L=4e-08 W=3.3e-07 
M7 3 C VSS VPW nch L=4e-08 W=3.3e-07 
M8 VSS C 3 VPW nch L=4e-08 W=3.3e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M13 VDD A 1 VNW pch L=4e-08 W=2.2e-07 
M14 1 B VDD VNW pch L=4e-08 W=2.2e-07 
M15 VDD B 1 VNW pch L=4e-08 W=2.2e-07 
M16 1 A VDD VNW pch L=4e-08 W=2.2e-07 
M17 VDD A 1 VNW pch L=4e-08 W=2.2e-07 
M18 1 B VDD VNW pch L=4e-08 W=2.2e-07 
M19 VDD C 1 VNW pch L=4e-08 W=2.2e-07 
M20 1 C VDD VNW pch L=4e-08 W=2.2e-07 
M21 VDD C 1 VNW pch L=4e-08 W=2.2e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M24 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND3_X6M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=3.7e-07 
M1 1 C VSS VPW nch L=4e-08 W=3.7e-07 
M2 VSS C 1 VPW nch L=4e-08 W=3.7e-07 
M3 1 C VSS VPW nch L=4e-08 W=3.7e-07 
M4 9 B 1 VPW nch L=4e-08 W=3.7e-07 
M5 4 A 9 VPW nch L=4e-08 W=3.7e-07 
M6 10 A 4 VPW nch L=4e-08 W=3.7e-07 
M7 1 B 10 VPW nch L=4e-08 W=3.7e-07 
M8 11 B 1 VPW nch L=4e-08 W=3.7e-07 
M9 4 A 11 VPW nch L=4e-08 W=3.7e-07 
M10 12 A 4 VPW nch L=4e-08 W=3.7e-07 
M11 1 B 12 VPW nch L=4e-08 W=3.7e-07 
M12 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M16 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M18 4 C VDD VNW pch L=4e-08 W=2.45e-07 
M19 VDD C 4 VNW pch L=4e-08 W=2.45e-07 
M20 4 C VDD VNW pch L=4e-08 W=2.45e-07 
M21 VDD C 4 VNW pch L=4e-08 W=2.45e-07 
M22 4 B VDD VNW pch L=4e-08 W=2.45e-07 
M23 VDD A 4 VNW pch L=4e-08 W=2.45e-07 
M24 4 A VDD VNW pch L=4e-08 W=2.45e-07 
M25 VDD B 4 VNW pch L=4e-08 W=2.45e-07 
M26 4 B VDD VNW pch L=4e-08 W=2.45e-07 
M27 VDD A 4 VNW pch L=4e-08 W=2.45e-07 
M28 4 A VDD VNW pch L=4e-08 W=2.45e-07 
M29 VDD B 4 VNW pch L=4e-08 W=2.45e-07 
M30 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M32 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M33 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M34 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND3_X8M_A9TR Y VDD VNW VPW VSS A B C
M0 9 A 1 VPW nch L=4e-08 W=4e-07 
M1 3 B 9 VPW nch L=4e-08 W=4e-07 
M2 10 B 3 VPW nch L=4e-08 W=4e-07 
M3 1 A 10 VPW nch L=4e-08 W=4e-07 
M4 11 A 1 VPW nch L=4e-08 W=4e-07 
M5 3 B 11 VPW nch L=4e-08 W=4e-07 
M6 12 B 3 VPW nch L=4e-08 W=4e-07 
M7 1 A 12 VPW nch L=4e-08 W=4e-07 
M8 13 A 1 VPW nch L=4e-08 W=4e-07 
M9 3 B 13 VPW nch L=4e-08 W=4e-07 
M10 VSS C 3 VPW nch L=4e-08 W=4e-07 
M11 3 C VSS VPW nch L=4e-08 W=4e-07 
M12 VSS C 3 VPW nch L=4e-08 W=4e-07 
M13 3 C VSS VPW nch L=4e-08 W=4e-07 
M14 VSS C 3 VPW nch L=4e-08 W=4e-07 
M15 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M17 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M18 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M19 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M20 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M21 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M22 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M23 VDD A 1 VNW pch L=4e-08 W=2.65e-07 
M24 1 B VDD VNW pch L=4e-08 W=2.65e-07 
M25 VDD B 1 VNW pch L=4e-08 W=2.65e-07 
M26 1 A VDD VNW pch L=4e-08 W=2.65e-07 
M27 VDD A 1 VNW pch L=4e-08 W=2.65e-07 
M28 1 B VDD VNW pch L=4e-08 W=2.65e-07 
M29 VDD B 1 VNW pch L=4e-08 W=2.65e-07 
M30 1 A VDD VNW pch L=4e-08 W=2.65e-07 
M31 VDD A 1 VNW pch L=4e-08 W=2.65e-07 
M32 1 B VDD VNW pch L=4e-08 W=2.65e-07 
M33 VDD C 1 VNW pch L=4e-08 W=2.65e-07 
M34 1 C VDD VNW pch L=4e-08 W=2.65e-07 
M35 VDD C 1 VNW pch L=4e-08 W=2.65e-07 
M36 1 C VDD VNW pch L=4e-08 W=2.65e-07 
M37 VDD C 1 VNW pch L=4e-08 W=2.65e-07 
M38 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M40 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M41 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M42 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M43 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M44 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M45 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND4_X0P5M_A9TR Y VDD VNW VPW VSS A B C D
M0 9 A 1 VPW nch L=4e-08 W=2.55e-07 
M1 10 B 9 VPW nch L=4e-08 W=2.55e-07 
M2 11 C 10 VPW nch L=4e-08 W=2.55e-07 
M3 VSS D 11 VPW nch L=4e-08 W=2.55e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.55e-07 
M5 1 A VDD VNW pch L=4e-08 W=1.45e-07 
M6 VDD B 1 VNW pch L=4e-08 W=1.45e-07 
M7 1 C VDD VNW pch L=4e-08 W=1.45e-07 
M8 VDD D 1 VNW pch L=4e-08 W=1.45e-07 
M9 Y 1 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AND4_X0P7M_A9TR Y VDD VNW VPW VSS A B C D
M0 9 A 1 VPW nch L=4e-08 W=3.15e-07 
M1 10 B 9 VPW nch L=4e-08 W=3.15e-07 
M2 11 C 10 VPW nch L=4e-08 W=3.15e-07 
M3 VSS D 11 VPW nch L=4e-08 W=3.15e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M5 1 A VDD VNW pch L=4e-08 W=1.8e-07 
M6 VDD B 1 VNW pch L=4e-08 W=1.8e-07 
M7 1 C VDD VNW pch L=4e-08 W=1.8e-07 
M8 VDD D 1 VNW pch L=4e-08 W=1.8e-07 
M9 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AND4_X1M_A9TR Y VDD VNW VPW VSS A B C D
M0 9 A 1 VPW nch L=4e-08 W=3.8e-07 
M1 10 B 9 VPW nch L=4e-08 W=3.8e-07 
M2 11 C 10 VPW nch L=4e-08 W=3.8e-07 
M3 VSS D 11 VPW nch L=4e-08 W=3.8e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M5 1 A VDD VNW pch L=4e-08 W=2.2e-07 
M6 VDD B 1 VNW pch L=4e-08 W=2.2e-07 
M7 1 C VDD VNW pch L=4e-08 W=2.2e-07 
M8 VDD D 1 VNW pch L=4e-08 W=2.2e-07 
M9 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND4_X1P4M_A9TR Y VDD VNW VPW VSS A B C D
M0 10 C 1 VPW nch L=4e-08 W=3.2e-07 
M1 VSS D 10 VPW nch L=4e-08 W=3.2e-07 
M2 11 D VSS VPW nch L=4e-08 W=3.2e-07 
M3 1 C 11 VPW nch L=4e-08 W=3.2e-07 
M4 12 B 1 VPW nch L=4e-08 W=3.2e-07 
M5 3 A 12 VPW nch L=4e-08 W=3.2e-07 
M6 13 A 3 VPW nch L=4e-08 W=3.2e-07 
M7 1 B 13 VPW nch L=4e-08 W=3.2e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=2.2e-07 
M9 VSS 3 Y VPW nch L=4e-08 W=2.2e-07 
M10 3 C VDD VNW pch L=4e-08 W=1.85e-07 
M11 VDD D 3 VNW pch L=4e-08 W=1.85e-07 
M12 3 D VDD VNW pch L=4e-08 W=1.85e-07 
M13 VDD C 3 VNW pch L=4e-08 W=1.85e-07 
M14 3 B VDD VNW pch L=4e-08 W=1.85e-07 
M15 VDD A 3 VNW pch L=4e-08 W=1.85e-07 
M16 3 A VDD VNW pch L=4e-08 W=1.85e-07 
M17 VDD B 3 VNW pch L=4e-08 W=1.85e-07 
M18 Y 3 VDD VNW pch L=4e-08 W=2.85e-07 
M19 VDD 3 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AND4_X2M_A9TR Y VDD VNW VPW VSS A B C D
M0 10 C 1 VPW nch L=4e-08 W=4e-07 
M1 VSS D 10 VPW nch L=4e-08 W=4e-07 
M2 11 D VSS VPW nch L=4e-08 W=4e-07 
M3 1 C 11 VPW nch L=4e-08 W=4e-07 
M4 12 B 1 VPW nch L=4e-08 W=4e-07 
M5 3 A 12 VPW nch L=4e-08 W=4e-07 
M6 13 A 3 VPW nch L=4e-08 W=4e-07 
M7 1 B 13 VPW nch L=4e-08 W=4e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M10 3 C VDD VNW pch L=4e-08 W=2.25e-07 
M11 VDD D 3 VNW pch L=4e-08 W=2.25e-07 
M12 3 D VDD VNW pch L=4e-08 W=2.25e-07 
M13 VDD C 3 VNW pch L=4e-08 W=2.25e-07 
M14 3 B VDD VNW pch L=4e-08 W=2.25e-07 
M15 VDD A 3 VNW pch L=4e-08 W=2.25e-07 
M16 3 A VDD VNW pch L=4e-08 W=2.25e-07 
M17 VDD B 3 VNW pch L=4e-08 W=2.25e-07 
M18 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND4_X3M_A9TR Y VDD VNW VPW VSS A B C D
M0 3 A 1 VPW nch L=4e-08 W=3.8e-07 
M1 1 A 3 VPW nch L=4e-08 W=3.8e-07 
M2 12 A 1 VPW nch L=4e-08 W=3.8e-07 
M3 4 B 12 VPW nch L=4e-08 W=3.8e-07 
M4 3 B 4 VPW nch L=4e-08 W=3.8e-07 
M5 4 B 3 VPW nch L=4e-08 W=3.8e-07 
M6 5 C 4 VPW nch L=4e-08 W=3.8e-07 
M7 4 C 5 VPW nch L=4e-08 W=3.8e-07 
M8 13 C 4 VPW nch L=4e-08 W=3.8e-07 
M9 VSS D 13 VPW nch L=4e-08 W=3.8e-07 
M10 5 D VSS VPW nch L=4e-08 W=3.8e-07 
M11 VSS D 5 VPW nch L=4e-08 W=3.8e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M15 1 A VDD VNW pch L=4e-08 W=2.15e-07 
M16 VDD A 1 VNW pch L=4e-08 W=2.15e-07 
M17 1 A VDD VNW pch L=4e-08 W=2.15e-07 
M18 VDD B 1 VNW pch L=4e-08 W=2.15e-07 
M19 1 B VDD VNW pch L=4e-08 W=2.15e-07 
M20 VDD B 1 VNW pch L=4e-08 W=2.15e-07 
M21 1 C VDD VNW pch L=4e-08 W=2.15e-07 
M22 VDD C 1 VNW pch L=4e-08 W=2.15e-07 
M23 1 C VDD VNW pch L=4e-08 W=2.15e-07 
M24 VDD D 1 VNW pch L=4e-08 W=2.15e-07 
M25 1 D VDD VNW pch L=4e-08 W=2.15e-07 
M26 VDD D 1 VNW pch L=4e-08 W=2.15e-07 
M27 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M29 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND4_X4M_A9TR Y VDD VNW VPW VSS A B C D
M0 10 C 1 VPW nch L=4e-08 W=3.7e-07 
M1 VSS D 10 VPW nch L=4e-08 W=3.7e-07 
M2 11 D VSS VPW nch L=4e-08 W=3.7e-07 
M3 1 C 11 VPW nch L=4e-08 W=3.7e-07 
M4 12 C 1 VPW nch L=4e-08 W=3.7e-07 
M5 VSS D 12 VPW nch L=4e-08 W=3.7e-07 
M6 13 D VSS VPW nch L=4e-08 W=3.7e-07 
M7 1 C 13 VPW nch L=4e-08 W=3.7e-07 
M8 14 B 1 VPW nch L=4e-08 W=3.7e-07 
M9 3 A 14 VPW nch L=4e-08 W=3.7e-07 
M10 15 A 3 VPW nch L=4e-08 W=3.7e-07 
M11 1 B 15 VPW nch L=4e-08 W=3.7e-07 
M12 16 B 1 VPW nch L=4e-08 W=3.7e-07 
M13 3 A 16 VPW nch L=4e-08 W=3.7e-07 
M14 17 A 3 VPW nch L=4e-08 W=3.7e-07 
M15 1 B 17 VPW nch L=4e-08 W=3.7e-07 
M16 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M18 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M20 3 C VDD VNW pch L=4e-08 W=2.1e-07 
M21 VDD D 3 VNW pch L=4e-08 W=2.1e-07 
M22 3 D VDD VNW pch L=4e-08 W=2.1e-07 
M23 VDD C 3 VNW pch L=4e-08 W=2.1e-07 
M24 3 C VDD VNW pch L=4e-08 W=2.1e-07 
M25 VDD D 3 VNW pch L=4e-08 W=2.1e-07 
M26 3 D VDD VNW pch L=4e-08 W=2.1e-07 
M27 VDD C 3 VNW pch L=4e-08 W=2.1e-07 
M28 3 B VDD VNW pch L=4e-08 W=2.1e-07 
M29 VDD A 3 VNW pch L=4e-08 W=2.1e-07 
M30 3 A VDD VNW pch L=4e-08 W=2.1e-07 
M31 VDD B 3 VNW pch L=4e-08 W=2.1e-07 
M32 3 B VDD VNW pch L=4e-08 W=2.1e-07 
M33 VDD A 3 VNW pch L=4e-08 W=2.1e-07 
M34 3 A VDD VNW pch L=4e-08 W=2.1e-07 
M35 VDD B 3 VNW pch L=4e-08 W=2.1e-07 
M36 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M38 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND4_X6M_A9TR Y VDD VNW VPW VSS A B C D
M0 10 C 1 VPW nch L=4e-08 W=3.75e-07 
M1 VSS D 10 VPW nch L=4e-08 W=3.75e-07 
M2 11 D VSS VPW nch L=4e-08 W=3.75e-07 
M3 1 C 11 VPW nch L=4e-08 W=3.75e-07 
M4 12 C 1 VPW nch L=4e-08 W=3.75e-07 
M5 VSS D 12 VPW nch L=4e-08 W=3.75e-07 
M6 13 D VSS VPW nch L=4e-08 W=3.75e-07 
M7 1 C 13 VPW nch L=4e-08 W=3.75e-07 
M8 14 C 1 VPW nch L=4e-08 W=3.75e-07 
M9 VSS D 14 VPW nch L=4e-08 W=3.75e-07 
M10 15 D VSS VPW nch L=4e-08 W=3.75e-07 
M11 1 C 15 VPW nch L=4e-08 W=3.75e-07 
M12 16 B 1 VPW nch L=4e-08 W=3.75e-07 
M13 3 A 16 VPW nch L=4e-08 W=3.75e-07 
M14 17 A 3 VPW nch L=4e-08 W=3.75e-07 
M15 1 B 17 VPW nch L=4e-08 W=3.75e-07 
M16 18 B 1 VPW nch L=4e-08 W=3.75e-07 
M17 3 A 18 VPW nch L=4e-08 W=3.75e-07 
M18 19 A 3 VPW nch L=4e-08 W=3.75e-07 
M19 1 B 19 VPW nch L=4e-08 W=3.75e-07 
M20 20 B 1 VPW nch L=4e-08 W=3.75e-07 
M21 3 A 20 VPW nch L=4e-08 W=3.75e-07 
M22 21 A 3 VPW nch L=4e-08 W=3.75e-07 
M23 1 B 21 VPW nch L=4e-08 W=3.75e-07 
M24 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M25 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M26 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M27 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M28 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M29 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M30 3 C VDD VNW pch L=4e-08 W=2.15e-07 
M31 VDD D 3 VNW pch L=4e-08 W=2.15e-07 
M32 3 D VDD VNW pch L=4e-08 W=2.15e-07 
M33 VDD C 3 VNW pch L=4e-08 W=2.15e-07 
M34 3 C VDD VNW pch L=4e-08 W=2.15e-07 
M35 VDD D 3 VNW pch L=4e-08 W=2.15e-07 
M36 3 D VDD VNW pch L=4e-08 W=2.15e-07 
M37 VDD C 3 VNW pch L=4e-08 W=2.15e-07 
M38 3 C VDD VNW pch L=4e-08 W=2.15e-07 
M39 VDD D 3 VNW pch L=4e-08 W=2.15e-07 
M40 3 D VDD VNW pch L=4e-08 W=2.15e-07 
M41 VDD C 3 VNW pch L=4e-08 W=2.15e-07 
M42 3 B VDD VNW pch L=4e-08 W=2.15e-07 
M43 VDD A 3 VNW pch L=4e-08 W=2.15e-07 
M44 3 A VDD VNW pch L=4e-08 W=2.15e-07 
M45 VDD B 3 VNW pch L=4e-08 W=2.15e-07 
M46 3 B VDD VNW pch L=4e-08 W=2.15e-07 
M47 VDD A 3 VNW pch L=4e-08 W=2.15e-07 
M48 3 A VDD VNW pch L=4e-08 W=2.15e-07 
M49 VDD B 3 VNW pch L=4e-08 W=2.15e-07 
M50 3 B VDD VNW pch L=4e-08 W=2.15e-07 
M51 VDD A 3 VNW pch L=4e-08 W=2.15e-07 
M52 3 A VDD VNW pch L=4e-08 W=2.15e-07 
M53 VDD B 3 VNW pch L=4e-08 W=2.15e-07 
M54 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M55 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M56 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M57 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M58 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M59 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AND4_X8M_A9TR Y VDD VNW VPW VSS A B C D
M0 10 C 1 VPW nch L=4e-08 W=3.75e-07 
M1 VSS D 10 VPW nch L=4e-08 W=3.75e-07 
M2 11 D VSS VPW nch L=4e-08 W=3.75e-07 
M3 1 C 11 VPW nch L=4e-08 W=3.75e-07 
M4 12 C 1 VPW nch L=4e-08 W=3.75e-07 
M5 VSS D 12 VPW nch L=4e-08 W=3.75e-07 
M6 13 D VSS VPW nch L=4e-08 W=3.75e-07 
M7 1 C 13 VPW nch L=4e-08 W=3.75e-07 
M8 14 C 1 VPW nch L=4e-08 W=3.75e-07 
M9 VSS D 14 VPW nch L=4e-08 W=3.75e-07 
M10 15 D VSS VPW nch L=4e-08 W=3.75e-07 
M11 1 C 15 VPW nch L=4e-08 W=3.75e-07 
M12 16 C 1 VPW nch L=4e-08 W=3.75e-07 
M13 VSS D 16 VPW nch L=4e-08 W=3.75e-07 
M14 17 D VSS VPW nch L=4e-08 W=3.75e-07 
M15 1 C 17 VPW nch L=4e-08 W=3.75e-07 
M16 18 B 1 VPW nch L=4e-08 W=3.75e-07 
M17 3 A 18 VPW nch L=4e-08 W=3.75e-07 
M18 19 A 3 VPW nch L=4e-08 W=3.75e-07 
M19 1 B 19 VPW nch L=4e-08 W=3.75e-07 
M20 20 B 1 VPW nch L=4e-08 W=3.75e-07 
M21 3 A 20 VPW nch L=4e-08 W=3.75e-07 
M22 21 A 3 VPW nch L=4e-08 W=3.75e-07 
M23 1 B 21 VPW nch L=4e-08 W=3.75e-07 
M24 22 B 1 VPW nch L=4e-08 W=3.75e-07 
M25 3 A 22 VPW nch L=4e-08 W=3.75e-07 
M26 23 A 3 VPW nch L=4e-08 W=3.75e-07 
M27 1 B 23 VPW nch L=4e-08 W=3.75e-07 
M28 24 B 1 VPW nch L=4e-08 W=3.75e-07 
M29 3 A 24 VPW nch L=4e-08 W=3.75e-07 
M30 25 A 3 VPW nch L=4e-08 W=3.75e-07 
M31 1 B 25 VPW nch L=4e-08 W=3.75e-07 
M32 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M33 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M34 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M35 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M36 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M37 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M38 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M39 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M40 3 C VDD VNW pch L=4e-08 W=2.15e-07 
M41 VDD D 3 VNW pch L=4e-08 W=2.15e-07 
M42 3 D VDD VNW pch L=4e-08 W=2.15e-07 
M43 VDD C 3 VNW pch L=4e-08 W=2.15e-07 
M44 3 C VDD VNW pch L=4e-08 W=2.15e-07 
M45 VDD D 3 VNW pch L=4e-08 W=2.15e-07 
M46 3 D VDD VNW pch L=4e-08 W=2.15e-07 
M47 VDD C 3 VNW pch L=4e-08 W=2.15e-07 
M48 3 C VDD VNW pch L=4e-08 W=2.15e-07 
M49 VDD D 3 VNW pch L=4e-08 W=2.15e-07 
M50 3 D VDD VNW pch L=4e-08 W=2.15e-07 
M51 VDD C 3 VNW pch L=4e-08 W=2.15e-07 
M52 3 C VDD VNW pch L=4e-08 W=2.15e-07 
M53 VDD D 3 VNW pch L=4e-08 W=2.15e-07 
M54 3 D VDD VNW pch L=4e-08 W=2.15e-07 
M55 VDD C 3 VNW pch L=4e-08 W=2.15e-07 
M56 3 B VDD VNW pch L=4e-08 W=2.15e-07 
M57 VDD A 3 VNW pch L=4e-08 W=2.15e-07 
M58 3 A VDD VNW pch L=4e-08 W=2.15e-07 
M59 VDD B 3 VNW pch L=4e-08 W=2.15e-07 
M60 3 B VDD VNW pch L=4e-08 W=2.15e-07 
M61 VDD A 3 VNW pch L=4e-08 W=2.15e-07 
M62 3 A VDD VNW pch L=4e-08 W=2.15e-07 
M63 VDD B 3 VNW pch L=4e-08 W=2.15e-07 
M64 3 B VDD VNW pch L=4e-08 W=2.15e-07 
M65 VDD A 3 VNW pch L=4e-08 W=2.15e-07 
M66 3 A VDD VNW pch L=4e-08 W=2.15e-07 
M67 VDD B 3 VNW pch L=4e-08 W=2.15e-07 
M68 3 B VDD VNW pch L=4e-08 W=2.15e-07 
M69 VDD A 3 VNW pch L=4e-08 W=2.15e-07 
M70 3 A VDD VNW pch L=4e-08 W=2.15e-07 
M71 VDD B 3 VNW pch L=4e-08 W=2.15e-07 
M72 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M73 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M74 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M75 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M76 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M77 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M78 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M79 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO1B2_X0P5M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 8 B0 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS B1 8 VPW nch L=4e-08 W=1.2e-07 
M2 9 A0N VSS VPW nch L=4e-08 W=1.75e-07 
M3 Y 1 9 VPW nch L=4e-08 W=1.75e-07 
M4 1 B0 VDD VNW pch L=4e-08 W=1.35e-07 
M5 VDD B1 1 VNW pch L=4e-08 W=1.35e-07 
M6 Y A0N VDD VNW pch L=4e-08 W=1.95e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=1.95e-07 
.ENDS


.SUBCKT AO1B2_X0P7M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 8 B0 1 VPW nch L=4e-08 W=1.25e-07 
M1 VSS B1 8 VPW nch L=4e-08 W=1.25e-07 
M2 9 A0N VSS VPW nch L=4e-08 W=2.5e-07 
M3 Y 1 9 VPW nch L=4e-08 W=2.5e-07 
M4 1 B0 VDD VNW pch L=4e-08 W=1.35e-07 
M5 VDD B1 1 VNW pch L=4e-08 W=1.35e-07 
M6 Y A0N VDD VNW pch L=4e-08 W=2.75e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT AO1B2_X1M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 8 B0 1 VPW nch L=4e-08 W=1.6e-07 
M1 VSS B1 8 VPW nch L=4e-08 W=1.6e-07 
M2 9 A0N VSS VPW nch L=4e-08 W=3.55e-07 
M3 Y 1 9 VPW nch L=4e-08 W=3.55e-07 
M4 1 B0 VDD VNW pch L=4e-08 W=1.75e-07 
M5 VDD B1 1 VNW pch L=4e-08 W=1.75e-07 
M6 Y A0N VDD VNW pch L=4e-08 W=3.9e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT AO1B2_X1P4M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 8 B0 1 VPW nch L=4e-08 W=2.15e-07 
M1 VSS B1 8 VPW nch L=4e-08 W=2.15e-07 
M2 9 A0N VSS VPW nch L=4e-08 W=2.5e-07 
M3 Y 1 9 VPW nch L=4e-08 W=2.5e-07 
M4 10 1 Y VPW nch L=4e-08 W=2.5e-07 
M5 VSS A0N 10 VPW nch L=4e-08 W=2.5e-07 
M6 1 B0 VDD VNW pch L=4e-08 W=2.35e-07 
M7 VDD B1 1 VNW pch L=4e-08 W=2.35e-07 
M8 Y A0N VDD VNW pch L=4e-08 W=2.75e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=2.75e-07 
M10 Y 1 VDD VNW pch L=4e-08 W=2.75e-07 
M11 VDD A0N Y VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT AO1B2_X2M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 8 B0 1 VPW nch L=4e-08 W=2.85e-07 
M1 VSS B1 8 VPW nch L=4e-08 W=2.85e-07 
M2 9 A0N VSS VPW nch L=4e-08 W=3.55e-07 
M3 Y 1 9 VPW nch L=4e-08 W=3.55e-07 
M4 10 1 Y VPW nch L=4e-08 W=3.55e-07 
M5 VSS A0N 10 VPW nch L=4e-08 W=3.55e-07 
M6 1 B0 VDD VNW pch L=4e-08 W=3.15e-07 
M7 VDD B1 1 VNW pch L=4e-08 W=3.15e-07 
M8 Y A0N VDD VNW pch L=4e-08 W=3.9e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=3.9e-07 
M10 Y 1 VDD VNW pch L=4e-08 W=3.9e-07 
M11 VDD A0N Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT AO1B2_X3M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 8 B1 VSS VPW nch L=4e-08 W=2.25e-07 
M1 3 B0 8 VPW nch L=4e-08 W=2.25e-07 
M2 9 B0 3 VPW nch L=4e-08 W=2.25e-07 
M3 VSS B1 9 VPW nch L=4e-08 W=2.25e-07 
M4 10 A0N VSS VPW nch L=4e-08 W=3.55e-07 
M5 Y 3 10 VPW nch L=4e-08 W=3.55e-07 
M6 11 3 Y VPW nch L=4e-08 W=3.55e-07 
M7 VSS A0N 11 VPW nch L=4e-08 W=3.55e-07 
M8 12 A0N VSS VPW nch L=4e-08 W=3.55e-07 
M9 Y 3 12 VPW nch L=4e-08 W=3.55e-07 
M10 3 B1 VDD VNW pch L=4e-08 W=2.45e-07 
M11 VDD B0 3 VNW pch L=4e-08 W=2.45e-07 
M12 3 B0 VDD VNW pch L=4e-08 W=2.45e-07 
M13 VDD B1 3 VNW pch L=4e-08 W=2.45e-07 
M14 Y A0N VDD VNW pch L=4e-08 W=3.9e-07 
M15 VDD 3 Y VNW pch L=4e-08 W=3.9e-07 
M16 Y 3 VDD VNW pch L=4e-08 W=3.9e-07 
M17 VDD A0N Y VNW pch L=4e-08 W=3.9e-07 
M18 Y A0N VDD VNW pch L=4e-08 W=3.9e-07 
M19 VDD 3 Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT AO1B2_X4M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 8 B1 VSS VPW nch L=4e-08 W=2.9e-07 
M1 3 B0 8 VPW nch L=4e-08 W=2.9e-07 
M2 9 B0 3 VPW nch L=4e-08 W=2.9e-07 
M3 VSS B1 9 VPW nch L=4e-08 W=2.9e-07 
M4 10 A0N VSS VPW nch L=4e-08 W=3.55e-07 
M5 Y 3 10 VPW nch L=4e-08 W=3.55e-07 
M6 11 3 Y VPW nch L=4e-08 W=3.55e-07 
M7 VSS A0N 11 VPW nch L=4e-08 W=3.55e-07 
M8 12 A0N VSS VPW nch L=4e-08 W=3.55e-07 
M9 Y 3 12 VPW nch L=4e-08 W=3.55e-07 
M10 13 3 Y VPW nch L=4e-08 W=3.55e-07 
M11 VSS A0N 13 VPW nch L=4e-08 W=3.55e-07 
M12 3 B1 VDD VNW pch L=4e-08 W=3.2e-07 
M13 VDD B0 3 VNW pch L=4e-08 W=3.2e-07 
M14 3 B0 VDD VNW pch L=4e-08 W=3.2e-07 
M15 VDD B1 3 VNW pch L=4e-08 W=3.2e-07 
M16 Y A0N VDD VNW pch L=4e-08 W=3.9e-07 
M17 VDD 3 Y VNW pch L=4e-08 W=3.9e-07 
M18 Y 3 VDD VNW pch L=4e-08 W=3.9e-07 
M19 VDD A0N Y VNW pch L=4e-08 W=3.9e-07 
M20 Y A0N VDD VNW pch L=4e-08 W=3.9e-07 
M21 VDD 3 Y VNW pch L=4e-08 W=3.9e-07 
M22 Y 3 VDD VNW pch L=4e-08 W=3.9e-07 
M23 VDD A0N Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT AO1B2_X6M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 8 B0 1 VPW nch L=4e-08 W=2.95e-07 
M1 VSS B1 8 VPW nch L=4e-08 W=2.95e-07 
M2 9 B1 VSS VPW nch L=4e-08 W=2.95e-07 
M3 1 B0 9 VPW nch L=4e-08 W=2.95e-07 
M4 10 B0 1 VPW nch L=4e-08 W=2.95e-07 
M5 VSS B1 10 VPW nch L=4e-08 W=2.95e-07 
M6 11 A0N VSS VPW nch L=4e-08 W=3.55e-07 
M7 Y 1 11 VPW nch L=4e-08 W=3.55e-07 
M8 12 1 Y VPW nch L=4e-08 W=3.55e-07 
M9 VSS A0N 12 VPW nch L=4e-08 W=3.55e-07 
M10 13 A0N VSS VPW nch L=4e-08 W=3.55e-07 
M11 Y 1 13 VPW nch L=4e-08 W=3.55e-07 
M12 14 1 Y VPW nch L=4e-08 W=3.55e-07 
M13 VSS A0N 14 VPW nch L=4e-08 W=3.55e-07 
M14 15 A0N VSS VPW nch L=4e-08 W=3.55e-07 
M15 Y 1 15 VPW nch L=4e-08 W=3.55e-07 
M16 16 1 Y VPW nch L=4e-08 W=3.55e-07 
M17 VSS A0N 16 VPW nch L=4e-08 W=3.55e-07 
M18 1 B0 VDD VNW pch L=4e-08 W=3.25e-07 
M19 VDD B1 1 VNW pch L=4e-08 W=3.25e-07 
M20 1 B1 VDD VNW pch L=4e-08 W=3.25e-07 
M21 VDD B0 1 VNW pch L=4e-08 W=3.25e-07 
M22 1 B0 VDD VNW pch L=4e-08 W=3.25e-07 
M23 VDD B1 1 VNW pch L=4e-08 W=3.25e-07 
M24 Y A0N VDD VNW pch L=4e-08 W=3.4e-07 
M25 VDD 1 Y VNW pch L=4e-08 W=3.4e-07 
M26 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD A0N Y VNW pch L=4e-08 W=4e-07 
M28 Y A0N VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M30 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD A0N Y VNW pch L=4e-08 W=4e-07 
M32 Y A0N VDD VNW pch L=4e-08 W=4e-07 
M33 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M34 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD A0N Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO21A1AI2_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A0 1 VPW nch L=4e-08 W=1.8e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=1.8e-07 
M2 1 B0 VSS VPW nch L=4e-08 W=1.4e-07 
M3 Y C0 1 VPW nch L=4e-08 W=1.7e-07 
M4 VDD A0 2 VNW pch L=4e-08 W=2.3e-07 
M5 2 A1 VDD VNW pch L=4e-08 W=2.3e-07 
M6 Y B0 2 VNW pch L=4e-08 W=2.3e-07 
M7 VDD C0 Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT AO21A1AI2_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A0 1 VPW nch L=4e-08 W=2.2e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=2.2e-07 
M2 1 B0 VSS VPW nch L=4e-08 W=1.7e-07 
M3 Y C0 1 VPW nch L=4e-08 W=2.2e-07 
M4 VDD A0 2 VNW pch L=4e-08 W=2.85e-07 
M5 2 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M6 Y B0 2 VNW pch L=4e-08 W=2.85e-07 
M7 VDD C0 Y VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT AO21A1AI2_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A0 1 VPW nch L=4e-08 W=3.1e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=3.1e-07 
M2 1 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y C0 1 VPW nch L=4e-08 W=3.1e-07 
M4 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M5 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M6 Y B0 2 VNW pch L=4e-08 W=4e-07 
M7 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT AO21A1AI2_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A0 1 VPW nch L=4e-08 W=2.2e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=2.2e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=2.2e-07 
M3 1 A0 11 VPW nch L=4e-08 W=2.2e-07 
M4 VSS B0 1 VPW nch L=4e-08 W=1.7e-07 
M5 1 B0 VSS VPW nch L=4e-08 W=1.7e-07 
M6 Y C0 1 VPW nch L=4e-08 W=2.2e-07 
M7 1 C0 Y VPW nch L=4e-08 W=2.2e-07 
M8 VDD A0 2 VNW pch L=4e-08 W=2.85e-07 
M9 2 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M10 VDD A1 2 VNW pch L=4e-08 W=2.85e-07 
M11 2 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M12 Y B0 2 VNW pch L=4e-08 W=2.85e-07 
M13 2 B0 Y VNW pch L=4e-08 W=2.85e-07 
M14 Y C0 VDD VNW pch L=4e-08 W=1.5e-07 
M15 VDD C0 Y VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT AO21A1AI2_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A0 1 VPW nch L=4e-08 W=3.1e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=3.1e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M3 1 A0 11 VPW nch L=4e-08 W=3.1e-07 
M4 VSS B0 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M6 Y C0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 C0 Y VPW nch L=4e-08 W=3.1e-07 
M8 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M9 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M11 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M12 Y B0 2 VNW pch L=4e-08 W=4e-07 
M13 2 B0 Y VNW pch L=4e-08 W=4e-07 
M14 VDD C0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO21A1AI2_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A0 1 VPW nch L=4e-08 W=3.1e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=3.1e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M3 1 A0 11 VPW nch L=4e-08 W=3.1e-07 
M4 12 A0 1 VPW nch L=4e-08 W=3.1e-07 
M5 VSS A1 12 VPW nch L=4e-08 W=3.1e-07 
M6 1 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M7 VSS B0 1 VPW nch L=4e-08 W=2.4e-07 
M8 1 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M9 Y C0 1 VPW nch L=4e-08 W=3.1e-07 
M10 1 C0 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y C0 1 VPW nch L=4e-08 W=3.1e-07 
M12 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M13 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M15 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M17 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M18 Y B0 2 VNW pch L=4e-08 W=4e-07 
M19 2 B0 Y VNW pch L=4e-08 W=4e-07 
M20 Y B0 2 VNW pch L=4e-08 W=4e-07 
M21 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
M22 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
M23 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT AO21A1AI2_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A0 1 VPW nch L=4e-08 W=3.1e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=3.1e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M3 1 A0 11 VPW nch L=4e-08 W=3.1e-07 
M4 12 A0 1 VPW nch L=4e-08 W=3.1e-07 
M5 VSS A1 12 VPW nch L=4e-08 W=3.1e-07 
M6 13 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M7 1 A0 13 VPW nch L=4e-08 W=3.1e-07 
M8 VSS B0 1 VPW nch L=4e-08 W=2.4e-07 
M9 1 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M10 VSS B0 1 VPW nch L=4e-08 W=2.4e-07 
M11 1 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M12 Y C0 1 VPW nch L=4e-08 W=3.1e-07 
M13 1 C0 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y C0 1 VPW nch L=4e-08 W=3.1e-07 
M15 1 C0 Y VPW nch L=4e-08 W=3.1e-07 
M16 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M17 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M19 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M21 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M23 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M24 Y B0 2 VNW pch L=4e-08 W=4e-07 
M25 2 B0 Y VNW pch L=4e-08 W=4e-07 
M26 Y B0 2 VNW pch L=4e-08 W=4e-07 
M27 2 B0 Y VNW pch L=4e-08 W=4e-07 
M28 VDD C0 Y VNW pch L=4e-08 W=2.8e-07 
M29 Y C0 VDD VNW pch L=4e-08 W=2.8e-07 
M30 VDD C0 Y VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT AO21A1AI2_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 11 A0 1 VPW nch L=4e-08 W=3.1e-07 
M1 VSS A1 11 VPW nch L=4e-08 W=3.1e-07 
M2 12 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M3 1 A0 12 VPW nch L=4e-08 W=3.1e-07 
M4 13 A0 1 VPW nch L=4e-08 W=3.1e-07 
M5 VSS A1 13 VPW nch L=4e-08 W=3.1e-07 
M6 14 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M7 1 A0 14 VPW nch L=4e-08 W=3.1e-07 
M8 15 A0 1 VPW nch L=4e-08 W=3.1e-07 
M9 VSS A1 15 VPW nch L=4e-08 W=3.1e-07 
M10 16 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M11 1 A0 16 VPW nch L=4e-08 W=3.1e-07 
M12 VSS B0 1 VPW nch L=4e-08 W=2.4e-07 
M13 1 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M14 VSS B0 1 VPW nch L=4e-08 W=2.4e-07 
M15 1 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M16 VSS B0 1 VPW nch L=4e-08 W=2.4e-07 
M17 1 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M18 Y C0 1 VPW nch L=4e-08 W=3.1e-07 
M19 1 C0 Y VPW nch L=4e-08 W=3.1e-07 
M20 Y C0 1 VPW nch L=4e-08 W=3.1e-07 
M21 1 C0 Y VPW nch L=4e-08 W=3.1e-07 
M22 Y C0 1 VPW nch L=4e-08 W=3.1e-07 
M23 1 C0 Y VPW nch L=4e-08 W=3.1e-07 
M24 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M25 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M27 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M29 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M31 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M33 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M35 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M36 Y B0 2 VNW pch L=4e-08 W=4e-07 
M37 2 B0 Y VNW pch L=4e-08 W=4e-07 
M38 Y B0 2 VNW pch L=4e-08 W=4e-07 
M39 2 B0 Y VNW pch L=4e-08 W=4e-07 
M40 Y B0 2 VNW pch L=4e-08 W=4e-07 
M41 2 B0 Y VNW pch L=4e-08 W=4e-07 
M42 Y C0 VDD VNW pch L=4e-08 W=3.15e-07 
M43 VDD C0 Y VNW pch L=4e-08 W=3.15e-07 
M44 Y C0 VDD VNW pch L=4e-08 W=3.15e-07 
M45 VDD C0 Y VNW pch L=4e-08 W=3.15e-07 
.ENDS


.SUBCKT AO21B_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 8 A0 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=1.2e-07 
M2 9 1 VSS VPW nch L=4e-08 W=1.75e-07 
M3 Y B0N 9 VPW nch L=4e-08 W=1.75e-07 
M4 1 A0 VDD VNW pch L=4e-08 W=1.35e-07 
M5 VDD A1 1 VNW pch L=4e-08 W=1.35e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=1.95e-07 
M7 VDD B0N Y VNW pch L=4e-08 W=1.95e-07 
.ENDS


.SUBCKT AO21B_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 8 A0 1 VPW nch L=4e-08 W=1.25e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=1.25e-07 
M2 9 1 VSS VPW nch L=4e-08 W=2.5e-07 
M3 Y B0N 9 VPW nch L=4e-08 W=2.5e-07 
M4 1 A0 VDD VNW pch L=4e-08 W=1.35e-07 
M5 VDD A1 1 VNW pch L=4e-08 W=1.35e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=2.75e-07 
M7 VDD B0N Y VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT AO21B_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 8 A0 1 VPW nch L=4e-08 W=1.6e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=1.6e-07 
M2 9 1 VSS VPW nch L=4e-08 W=3.55e-07 
M3 Y B0N 9 VPW nch L=4e-08 W=3.55e-07 
M4 1 A0 VDD VNW pch L=4e-08 W=1.75e-07 
M5 VDD A1 1 VNW pch L=4e-08 W=1.75e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=3.9e-07 
M7 VDD B0N Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT AO21B_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 8 A0 1 VPW nch L=4e-08 W=2.15e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=2.15e-07 
M2 9 1 VSS VPW nch L=4e-08 W=2.5e-07 
M3 Y B0N 9 VPW nch L=4e-08 W=2.5e-07 
M4 10 B0N Y VPW nch L=4e-08 W=2.5e-07 
M5 VSS 1 10 VPW nch L=4e-08 W=2.5e-07 
M6 1 A0 VDD VNW pch L=4e-08 W=2.35e-07 
M7 VDD A1 1 VNW pch L=4e-08 W=2.35e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=2.75e-07 
M9 VDD B0N Y VNW pch L=4e-08 W=2.75e-07 
M10 Y B0N VDD VNW pch L=4e-08 W=2.75e-07 
M11 VDD 1 Y VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT AO21B_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 8 A0 1 VPW nch L=4e-08 W=2.85e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=2.85e-07 
M2 9 1 VSS VPW nch L=4e-08 W=3.55e-07 
M3 Y B0N 9 VPW nch L=4e-08 W=3.55e-07 
M4 10 B0N Y VPW nch L=4e-08 W=3.55e-07 
M5 VSS 1 10 VPW nch L=4e-08 W=3.55e-07 
M6 1 A0 VDD VNW pch L=4e-08 W=3.15e-07 
M7 VDD A1 1 VNW pch L=4e-08 W=3.15e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=3.9e-07 
M9 VDD B0N Y VNW pch L=4e-08 W=3.9e-07 
M10 Y B0N VDD VNW pch L=4e-08 W=3.9e-07 
M11 VDD 1 Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT AO21B_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 8 A1 VSS VPW nch L=4e-08 W=2.25e-07 
M1 3 A0 8 VPW nch L=4e-08 W=2.25e-07 
M2 9 A0 3 VPW nch L=4e-08 W=2.25e-07 
M3 VSS A1 9 VPW nch L=4e-08 W=2.25e-07 
M4 10 3 VSS VPW nch L=4e-08 W=3.55e-07 
M5 Y B0N 10 VPW nch L=4e-08 W=3.55e-07 
M6 11 B0N Y VPW nch L=4e-08 W=3.55e-07 
M7 VSS 3 11 VPW nch L=4e-08 W=3.55e-07 
M8 12 3 VSS VPW nch L=4e-08 W=3.55e-07 
M9 Y B0N 12 VPW nch L=4e-08 W=3.55e-07 
M10 3 A1 VDD VNW pch L=4e-08 W=2.45e-07 
M11 VDD A0 3 VNW pch L=4e-08 W=2.45e-07 
M12 3 A0 VDD VNW pch L=4e-08 W=2.45e-07 
M13 VDD A1 3 VNW pch L=4e-08 W=2.45e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=3.9e-07 
M15 VDD B0N Y VNW pch L=4e-08 W=3.9e-07 
M16 Y B0N VDD VNW pch L=4e-08 W=3.9e-07 
M17 VDD 3 Y VNW pch L=4e-08 W=3.9e-07 
M18 Y 3 VDD VNW pch L=4e-08 W=3.9e-07 
M19 VDD B0N Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT AO21B_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 8 A1 VSS VPW nch L=4e-08 W=2.9e-07 
M1 3 A0 8 VPW nch L=4e-08 W=2.9e-07 
M2 9 A0 3 VPW nch L=4e-08 W=2.9e-07 
M3 VSS A1 9 VPW nch L=4e-08 W=2.9e-07 
M4 10 3 VSS VPW nch L=4e-08 W=3.55e-07 
M5 Y B0N 10 VPW nch L=4e-08 W=3.55e-07 
M6 11 B0N Y VPW nch L=4e-08 W=3.55e-07 
M7 VSS 3 11 VPW nch L=4e-08 W=3.55e-07 
M8 12 3 VSS VPW nch L=4e-08 W=3.55e-07 
M9 Y B0N 12 VPW nch L=4e-08 W=3.55e-07 
M10 13 B0N Y VPW nch L=4e-08 W=3.55e-07 
M11 VSS 3 13 VPW nch L=4e-08 W=3.55e-07 
M12 3 A1 VDD VNW pch L=4e-08 W=3.2e-07 
M13 VDD A0 3 VNW pch L=4e-08 W=3.2e-07 
M14 3 A0 VDD VNW pch L=4e-08 W=3.2e-07 
M15 VDD A1 3 VNW pch L=4e-08 W=3.2e-07 
M16 Y 3 VDD VNW pch L=4e-08 W=3.9e-07 
M17 VDD B0N Y VNW pch L=4e-08 W=3.9e-07 
M18 Y B0N VDD VNW pch L=4e-08 W=3.9e-07 
M19 VDD 3 Y VNW pch L=4e-08 W=3.9e-07 
M20 Y 3 VDD VNW pch L=4e-08 W=3.9e-07 
M21 VDD B0N Y VNW pch L=4e-08 W=3.9e-07 
M22 Y B0N VDD VNW pch L=4e-08 W=3.9e-07 
M23 VDD 3 Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT AO21B_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 8 A0 1 VPW nch L=4e-08 W=2.95e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=2.95e-07 
M2 9 A1 VSS VPW nch L=4e-08 W=2.95e-07 
M3 1 A0 9 VPW nch L=4e-08 W=2.95e-07 
M4 10 A0 1 VPW nch L=4e-08 W=2.95e-07 
M5 VSS A1 10 VPW nch L=4e-08 W=2.95e-07 
M6 11 1 VSS VPW nch L=4e-08 W=3.55e-07 
M7 Y B0N 11 VPW nch L=4e-08 W=3.55e-07 
M8 12 B0N Y VPW nch L=4e-08 W=3.55e-07 
M9 VSS 1 12 VPW nch L=4e-08 W=3.55e-07 
M10 13 1 VSS VPW nch L=4e-08 W=3.55e-07 
M11 Y B0N 13 VPW nch L=4e-08 W=3.55e-07 
M12 14 B0N Y VPW nch L=4e-08 W=3.55e-07 
M13 VSS 1 14 VPW nch L=4e-08 W=3.55e-07 
M14 15 1 VSS VPW nch L=4e-08 W=3.55e-07 
M15 Y B0N 15 VPW nch L=4e-08 W=3.55e-07 
M16 16 B0N Y VPW nch L=4e-08 W=3.55e-07 
M17 VSS 1 16 VPW nch L=4e-08 W=3.55e-07 
M18 1 A0 VDD VNW pch L=4e-08 W=3.25e-07 
M19 VDD A1 1 VNW pch L=4e-08 W=3.25e-07 
M20 1 A1 VDD VNW pch L=4e-08 W=3.25e-07 
M21 VDD A0 1 VNW pch L=4e-08 W=3.25e-07 
M22 1 A0 VDD VNW pch L=4e-08 W=3.25e-07 
M23 VDD A1 1 VNW pch L=4e-08 W=3.25e-07 
M24 Y 1 VDD VNW pch L=4e-08 W=3.9e-07 
M25 VDD B0N Y VNW pch L=4e-08 W=3.9e-07 
M26 Y B0N VDD VNW pch L=4e-08 W=3.9e-07 
M27 VDD 1 Y VNW pch L=4e-08 W=3.9e-07 
M28 Y 1 VDD VNW pch L=4e-08 W=3.9e-07 
M29 VDD B0N Y VNW pch L=4e-08 W=3.9e-07 
M30 Y B0N VDD VNW pch L=4e-08 W=3.9e-07 
M31 VDD 1 Y VNW pch L=4e-08 W=3.9e-07 
M32 Y 1 VDD VNW pch L=4e-08 W=3.9e-07 
M33 VDD B0N Y VNW pch L=4e-08 W=3.9e-07 
M34 Y B0N VDD VNW pch L=4e-08 W=3.9e-07 
M35 VDD 1 Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT AO21_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 9 A1 VSS VPW nch L=4e-08 W=1.8e-07 
M1 4 A0 9 VPW nch L=4e-08 W=1.8e-07 
M2 VSS B0 4 VPW nch L=4e-08 W=1.2e-07 
M3 Y 4 VSS VPW nch L=4e-08 W=1.55e-07 
M4 VDD A1 2 VNW pch L=4e-08 W=3e-07 
M5 2 A0 VDD VNW pch L=4e-08 W=3e-07 
M6 4 B0 2 VNW pch L=4e-08 W=3e-07 
M7 Y 4 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AO21_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 9 A1 VSS VPW nch L=4e-08 W=1.8e-07 
M1 4 A0 9 VPW nch L=4e-08 W=1.8e-07 
M2 VSS B0 4 VPW nch L=4e-08 W=1.2e-07 
M3 Y 4 VSS VPW nch L=4e-08 W=2.2e-07 
M4 VDD A1 2 VNW pch L=4e-08 W=3e-07 
M5 2 A0 VDD VNW pch L=4e-08 W=3e-07 
M6 4 B0 2 VNW pch L=4e-08 W=3e-07 
M7 Y 4 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AO21_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 9 A1 VSS VPW nch L=4e-08 W=2.05e-07 
M1 4 A0 9 VPW nch L=4e-08 W=2.05e-07 
M2 VSS B0 4 VPW nch L=4e-08 W=1.35e-07 
M3 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VDD A1 2 VNW pch L=4e-08 W=3.4e-07 
M5 2 A0 VDD VNW pch L=4e-08 W=3.4e-07 
M6 4 B0 2 VNW pch L=4e-08 W=3.4e-07 
M7 Y 4 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO21_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 10 A1 VSS VPW nch L=4e-08 W=3e-07 
M1 4 A0 10 VPW nch L=4e-08 W=3e-07 
M2 VSS B0 4 VPW nch L=4e-08 W=2e-07 
M3 Y 4 VSS VPW nch L=4e-08 W=2.2e-07 
M4 VSS 4 Y VPW nch L=4e-08 W=2.2e-07 
M5 VDD A0 1 VNW pch L=4e-08 W=2.5e-07 
M6 1 A1 VDD VNW pch L=4e-08 W=2.5e-07 
M7 VDD A1 1 VNW pch L=4e-08 W=2.5e-07 
M8 1 A0 VDD VNW pch L=4e-08 W=2.5e-07 
M9 4 B0 1 VNW pch L=4e-08 W=2.5e-07 
M10 1 B0 4 VNW pch L=4e-08 W=2.5e-07 
M11 Y 4 VDD VNW pch L=4e-08 W=2.85e-07 
M12 VDD 4 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AO21_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 9 A1 VSS VPW nch L=4e-08 W=1.95e-07 
M1 4 A0 9 VPW nch L=4e-08 W=1.95e-07 
M2 10 A0 4 VPW nch L=4e-08 W=1.95e-07 
M3 VSS A1 10 VPW nch L=4e-08 W=1.95e-07 
M4 4 B0 VSS VPW nch L=4e-08 W=1.3e-07 
M5 VSS B0 4 VPW nch L=4e-08 W=1.3e-07 
M6 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M8 VDD A1 2 VNW pch L=4e-08 W=3.2e-07 
M9 2 A0 VDD VNW pch L=4e-08 W=3.2e-07 
M10 VDD A0 2 VNW pch L=4e-08 W=3.2e-07 
M11 2 A1 VDD VNW pch L=4e-08 W=3.2e-07 
M12 4 B0 2 VNW pch L=4e-08 W=3.2e-07 
M13 2 B0 4 VNW pch L=4e-08 W=3.2e-07 
M14 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO21_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 9 A0 1 VPW nch L=4e-08 W=1.95e-07 
M1 VSS A1 9 VPW nch L=4e-08 W=1.95e-07 
M2 10 A1 VSS VPW nch L=4e-08 W=1.95e-07 
M3 1 A0 10 VPW nch L=4e-08 W=1.95e-07 
M4 11 A0 1 VPW nch L=4e-08 W=1.95e-07 
M5 VSS A1 11 VPW nch L=4e-08 W=1.95e-07 
M6 1 B0 VSS VPW nch L=4e-08 W=1.95e-07 
M7 VSS B0 1 VPW nch L=4e-08 W=1.95e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VDD A0 2 VNW pch L=4e-08 W=3.25e-07 
M12 2 A1 VDD VNW pch L=4e-08 W=3.25e-07 
M13 VDD A1 2 VNW pch L=4e-08 W=3.25e-07 
M14 2 A0 VDD VNW pch L=4e-08 W=3.25e-07 
M15 VDD A0 2 VNW pch L=4e-08 W=3.25e-07 
M16 2 A1 VDD VNW pch L=4e-08 W=3.25e-07 
M17 1 B0 2 VNW pch L=4e-08 W=3.25e-07 
M18 2 B0 1 VNW pch L=4e-08 W=3.25e-07 
M19 1 B0 2 VNW pch L=4e-08 W=3.25e-07 
M20 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO21_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 9 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M1 4 A0 9 VPW nch L=4e-08 W=2.4e-07 
M2 10 A0 4 VPW nch L=4e-08 W=2.4e-07 
M3 VSS A1 10 VPW nch L=4e-08 W=2.4e-07 
M4 11 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M5 4 A0 11 VPW nch L=4e-08 W=2.4e-07 
M6 VSS B0 4 VPW nch L=4e-08 W=2.4e-07 
M7 4 B0 VSS VPW nch L=4e-08 W=2.4e-07 
M8 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M10 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M12 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M13 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M15 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M17 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M18 4 B0 2 VNW pch L=4e-08 W=4e-07 
M19 2 B0 4 VNW pch L=4e-08 W=4e-07 
M20 4 B0 2 VNW pch L=4e-08 W=4e-07 
M21 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M23 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO21_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 9 A1 VSS VPW nch L=4e-08 W=2.25e-07 
M1 4 A0 9 VPW nch L=4e-08 W=2.25e-07 
M2 10 A0 4 VPW nch L=4e-08 W=2.25e-07 
M3 VSS A1 10 VPW nch L=4e-08 W=2.25e-07 
M4 11 A1 VSS VPW nch L=4e-08 W=2.25e-07 
M5 4 A0 11 VPW nch L=4e-08 W=2.25e-07 
M6 12 A0 4 VPW nch L=4e-08 W=2.25e-07 
M7 VSS A1 12 VPW nch L=4e-08 W=2.25e-07 
M8 13 A1 VSS VPW nch L=4e-08 W=2.25e-07 
M9 4 A0 13 VPW nch L=4e-08 W=2.25e-07 
M10 VSS B0 4 VPW nch L=4e-08 W=2.5e-07 
M11 4 B0 VSS VPW nch L=4e-08 W=2.5e-07 
M12 VSS B0 4 VPW nch L=4e-08 W=2.5e-07 
M13 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M15 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M17 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M18 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M19 VDD A1 2 VNW pch L=4e-08 W=3.75e-07 
M20 2 A0 VDD VNW pch L=4e-08 W=3.75e-07 
M21 VDD A0 2 VNW pch L=4e-08 W=3.75e-07 
M22 2 A1 VDD VNW pch L=4e-08 W=3.75e-07 
M23 VDD A1 2 VNW pch L=4e-08 W=3.75e-07 
M24 2 A0 VDD VNW pch L=4e-08 W=3.75e-07 
M25 VDD A0 2 VNW pch L=4e-08 W=3.75e-07 
M26 2 A1 VDD VNW pch L=4e-08 W=3.75e-07 
M27 VDD A1 2 VNW pch L=4e-08 W=3.75e-07 
M28 2 A0 VDD VNW pch L=4e-08 W=3.75e-07 
M29 4 B0 2 VNW pch L=4e-08 W=3.75e-07 
M30 2 B0 4 VNW pch L=4e-08 W=3.75e-07 
M31 4 B0 2 VNW pch L=4e-08 W=3.75e-07 
M32 2 B0 4 VNW pch L=4e-08 W=3.75e-07 
M33 4 B0 2 VNW pch L=4e-08 W=3.75e-07 
M34 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M36 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M38 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO22_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 10 A1 VSS VPW nch L=4e-08 W=1.35e-07 
M1 4 A0 10 VPW nch L=4e-08 W=1.35e-07 
M2 11 B0 4 VPW nch L=4e-08 W=1.35e-07 
M3 VSS B1 11 VPW nch L=4e-08 W=1.35e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=1.55e-07 
M5 VDD A1 2 VNW pch L=4e-08 W=2.25e-07 
M6 2 A0 VDD VNW pch L=4e-08 W=2.25e-07 
M7 4 B0 2 VNW pch L=4e-08 W=2.25e-07 
M8 2 B1 4 VNW pch L=4e-08 W=2.25e-07 
M9 Y 4 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AO22_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 10 A1 VSS VPW nch L=4e-08 W=1.7e-07 
M1 4 A0 10 VPW nch L=4e-08 W=1.7e-07 
M2 11 B0 4 VPW nch L=4e-08 W=1.7e-07 
M3 VSS B1 11 VPW nch L=4e-08 W=1.7e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=2.2e-07 
M5 VDD A1 2 VNW pch L=4e-08 W=2.8e-07 
M6 2 A0 VDD VNW pch L=4e-08 W=2.8e-07 
M7 4 B0 2 VNW pch L=4e-08 W=2.8e-07 
M8 2 B1 4 VNW pch L=4e-08 W=2.8e-07 
M9 Y 4 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AO22_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 10 A1 VSS VPW nch L=4e-08 W=2.15e-07 
M1 4 A0 10 VPW nch L=4e-08 W=2.15e-07 
M2 11 B0 4 VPW nch L=4e-08 W=2.15e-07 
M3 VSS B1 11 VPW nch L=4e-08 W=2.15e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M5 VDD A1 2 VNW pch L=4e-08 W=3.5e-07 
M6 2 A0 VDD VNW pch L=4e-08 W=3.5e-07 
M7 4 B0 2 VNW pch L=4e-08 W=3.5e-07 
M8 2 B1 4 VNW pch L=4e-08 W=3.5e-07 
M9 Y 4 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO22_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 11 A1 VSS VPW nch L=4e-08 W=3.4e-07 
M1 4 A0 11 VPW nch L=4e-08 W=3.4e-07 
M2 12 B0 4 VPW nch L=4e-08 W=3.4e-07 
M3 VSS B1 12 VPW nch L=4e-08 W=3.4e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=2.2e-07 
M5 VSS 4 Y VPW nch L=4e-08 W=2.2e-07 
M6 VDD A0 1 VNW pch L=4e-08 W=2.85e-07 
M7 1 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M8 VDD A1 1 VNW pch L=4e-08 W=2.85e-07 
M9 1 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M10 4 B0 1 VNW pch L=4e-08 W=2.85e-07 
M11 1 B1 4 VNW pch L=4e-08 W=2.85e-07 
M12 4 B1 1 VNW pch L=4e-08 W=2.85e-07 
M13 1 B0 4 VNW pch L=4e-08 W=2.85e-07 
M14 Y 4 VDD VNW pch L=4e-08 W=2.85e-07 
M15 VDD 4 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AO22_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 10 A1 VSS VPW nch L=4e-08 W=2.15e-07 
M1 4 A0 10 VPW nch L=4e-08 W=2.15e-07 
M2 11 A0 4 VPW nch L=4e-08 W=2.15e-07 
M3 VSS A1 11 VPW nch L=4e-08 W=2.15e-07 
M4 12 B1 VSS VPW nch L=4e-08 W=2.15e-07 
M5 4 B0 12 VPW nch L=4e-08 W=2.15e-07 
M6 13 B0 4 VPW nch L=4e-08 W=2.15e-07 
M7 VSS B1 13 VPW nch L=4e-08 W=2.15e-07 
M8 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M10 VDD A1 2 VNW pch L=4e-08 W=3.55e-07 
M11 2 A0 VDD VNW pch L=4e-08 W=3.55e-07 
M12 VDD A0 2 VNW pch L=4e-08 W=3.55e-07 
M13 2 A1 VDD VNW pch L=4e-08 W=3.55e-07 
M14 4 B1 2 VNW pch L=4e-08 W=3.55e-07 
M15 2 B0 4 VNW pch L=4e-08 W=3.55e-07 
M16 4 B0 2 VNW pch L=4e-08 W=3.55e-07 
M17 2 B1 4 VNW pch L=4e-08 W=3.55e-07 
M18 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO22_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 10 A0 1 VPW nch L=4e-08 W=2.25e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=2.25e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=2.25e-07 
M3 1 A0 11 VPW nch L=4e-08 W=2.25e-07 
M4 12 A0 1 VPW nch L=4e-08 W=2.25e-07 
M5 VSS A1 12 VPW nch L=4e-08 W=2.25e-07 
M6 13 B1 VSS VPW nch L=4e-08 W=2.25e-07 
M7 1 B0 13 VPW nch L=4e-08 W=2.25e-07 
M8 14 B0 1 VPW nch L=4e-08 W=2.25e-07 
M9 VSS B1 14 VPW nch L=4e-08 W=2.25e-07 
M10 15 B1 VSS VPW nch L=4e-08 W=2.25e-07 
M11 1 B0 15 VPW nch L=4e-08 W=2.25e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VDD A0 2 VNW pch L=4e-08 W=3.75e-07 
M16 2 A1 VDD VNW pch L=4e-08 W=3.75e-07 
M17 VDD A1 2 VNW pch L=4e-08 W=3.75e-07 
M18 2 A0 VDD VNW pch L=4e-08 W=3.75e-07 
M19 VDD A0 2 VNW pch L=4e-08 W=3.75e-07 
M20 2 A1 VDD VNW pch L=4e-08 W=3.75e-07 
M21 1 B1 2 VNW pch L=4e-08 W=3.75e-07 
M22 2 B0 1 VNW pch L=4e-08 W=3.75e-07 
M23 1 B0 2 VNW pch L=4e-08 W=3.75e-07 
M24 2 B1 1 VNW pch L=4e-08 W=3.75e-07 
M25 1 B1 2 VNW pch L=4e-08 W=3.75e-07 
M26 2 B0 1 VNW pch L=4e-08 W=3.75e-07 
M27 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M29 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO22_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 10 A0 1 VPW nch L=4e-08 W=2.15e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=2.15e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=2.15e-07 
M3 1 A0 11 VPW nch L=4e-08 W=2.15e-07 
M4 12 A0 1 VPW nch L=4e-08 W=2.15e-07 
M5 VSS A1 12 VPW nch L=4e-08 W=2.15e-07 
M6 13 A1 VSS VPW nch L=4e-08 W=2.15e-07 
M7 1 A0 13 VPW nch L=4e-08 W=2.15e-07 
M8 14 B0 1 VPW nch L=4e-08 W=2.15e-07 
M9 VSS B1 14 VPW nch L=4e-08 W=2.15e-07 
M10 15 B1 VSS VPW nch L=4e-08 W=2.15e-07 
M11 1 B0 15 VPW nch L=4e-08 W=2.15e-07 
M12 16 B0 1 VPW nch L=4e-08 W=2.15e-07 
M13 VSS B1 16 VPW nch L=4e-08 W=2.15e-07 
M14 17 B1 VSS VPW nch L=4e-08 W=2.15e-07 
M15 1 B0 17 VPW nch L=4e-08 W=2.15e-07 
M16 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M18 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M20 VDD A0 2 VNW pch L=4e-08 W=3.6e-07 
M21 2 A1 VDD VNW pch L=4e-08 W=3.6e-07 
M22 VDD A1 2 VNW pch L=4e-08 W=3.6e-07 
M23 2 A0 VDD VNW pch L=4e-08 W=3.6e-07 
M24 VDD A0 2 VNW pch L=4e-08 W=3.6e-07 
M25 2 A1 VDD VNW pch L=4e-08 W=3.6e-07 
M26 VDD A1 2 VNW pch L=4e-08 W=3.6e-07 
M27 2 A0 VDD VNW pch L=4e-08 W=3.6e-07 
M28 1 B0 2 VNW pch L=4e-08 W=3.6e-07 
M29 2 B1 1 VNW pch L=4e-08 W=3.6e-07 
M30 1 B1 2 VNW pch L=4e-08 W=3.6e-07 
M31 2 B0 1 VNW pch L=4e-08 W=3.6e-07 
M32 1 B0 2 VNW pch L=4e-08 W=3.6e-07 
M33 2 B1 1 VNW pch L=4e-08 W=3.6e-07 
M34 1 B1 2 VNW pch L=4e-08 W=3.6e-07 
M35 2 B0 1 VNW pch L=4e-08 W=3.6e-07 
M36 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M38 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AO22_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 10 A0 1 VPW nch L=4e-08 W=2.15e-07 
M1 VSS A1 10 VPW nch L=4e-08 W=2.15e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=2.15e-07 
M3 1 A0 11 VPW nch L=4e-08 W=2.15e-07 
M4 12 A0 1 VPW nch L=4e-08 W=2.15e-07 
M5 VSS A1 12 VPW nch L=4e-08 W=2.15e-07 
M6 13 A1 VSS VPW nch L=4e-08 W=2.15e-07 
M7 1 A0 13 VPW nch L=4e-08 W=2.15e-07 
M8 14 A0 1 VPW nch L=4e-08 W=2.15e-07 
M9 VSS A1 14 VPW nch L=4e-08 W=2.15e-07 
M10 15 A1 VSS VPW nch L=4e-08 W=2.15e-07 
M11 1 A0 15 VPW nch L=4e-08 W=2.15e-07 
M12 16 B0 1 VPW nch L=4e-08 W=2.15e-07 
M13 VSS B1 16 VPW nch L=4e-08 W=2.15e-07 
M14 17 B1 VSS VPW nch L=4e-08 W=2.15e-07 
M15 1 B0 17 VPW nch L=4e-08 W=2.15e-07 
M16 18 B0 1 VPW nch L=4e-08 W=2.15e-07 
M17 VSS B1 18 VPW nch L=4e-08 W=2.15e-07 
M18 19 B1 VSS VPW nch L=4e-08 W=2.15e-07 
M19 1 B0 19 VPW nch L=4e-08 W=2.15e-07 
M20 20 B0 1 VPW nch L=4e-08 W=2.15e-07 
M21 VSS B1 20 VPW nch L=4e-08 W=2.15e-07 
M22 21 B1 VSS VPW nch L=4e-08 W=2.15e-07 
M23 1 B0 21 VPW nch L=4e-08 W=2.15e-07 
M24 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M25 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M26 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M27 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M28 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M29 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M30 VDD A0 2 VNW pch L=4e-08 W=3.55e-07 
M31 2 A1 VDD VNW pch L=4e-08 W=3.55e-07 
M32 VDD A1 2 VNW pch L=4e-08 W=3.55e-07 
M33 2 A0 VDD VNW pch L=4e-08 W=3.55e-07 
M34 VDD A0 2 VNW pch L=4e-08 W=3.55e-07 
M35 2 A1 VDD VNW pch L=4e-08 W=3.55e-07 
M36 VDD A1 2 VNW pch L=4e-08 W=3.55e-07 
M37 2 A0 VDD VNW pch L=4e-08 W=3.55e-07 
M38 VDD A0 2 VNW pch L=4e-08 W=3.55e-07 
M39 2 A1 VDD VNW pch L=4e-08 W=3.55e-07 
M40 VDD A1 2 VNW pch L=4e-08 W=3.55e-07 
M41 2 A0 VDD VNW pch L=4e-08 W=3.55e-07 
M42 1 B0 2 VNW pch L=4e-08 W=3.55e-07 
M43 2 B1 1 VNW pch L=4e-08 W=3.55e-07 
M44 1 B1 2 VNW pch L=4e-08 W=3.55e-07 
M45 2 B0 1 VNW pch L=4e-08 W=3.55e-07 
M46 1 B0 2 VNW pch L=4e-08 W=3.55e-07 
M47 2 B1 1 VNW pch L=4e-08 W=3.55e-07 
M48 1 B1 2 VNW pch L=4e-08 W=3.55e-07 
M49 2 B0 1 VNW pch L=4e-08 W=3.55e-07 
M50 1 B0 2 VNW pch L=4e-08 W=3.55e-07 
M51 2 B1 1 VNW pch L=4e-08 W=3.55e-07 
M52 1 B1 2 VNW pch L=4e-08 W=3.55e-07 
M53 2 B0 1 VNW pch L=4e-08 W=3.55e-07 
M54 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M55 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M56 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M57 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M58 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M59 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI211_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A0 10 VPW nch L=4e-08 W=1.2e-07 
M2 VSS B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 Y C0 VSS VPW nch L=4e-08 W=1.2e-07 
M4 VDD A1 2 VNW pch L=4e-08 W=2e-07 
M5 2 A0 VDD VNW pch L=4e-08 W=2e-07 
M6 9 B0 2 VNW pch L=4e-08 W=2e-07 
M7 Y C0 9 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AOI211_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A0 10 VPW nch L=4e-08 W=1.2e-07 
M2 VSS B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 Y C0 VSS VPW nch L=4e-08 W=1.2e-07 
M4 VDD A1 2 VNW pch L=4e-08 W=2.85e-07 
M5 2 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M6 9 B0 2 VNW pch L=4e-08 W=2.85e-07 
M7 Y C0 9 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI211_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 10 A1 VSS VPW nch L=4e-08 W=1.8e-07 
M1 Y A0 10 VPW nch L=4e-08 W=1.8e-07 
M2 VSS B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 Y C0 VSS VPW nch L=4e-08 W=1.2e-07 
M4 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M5 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M6 9 B0 2 VNW pch L=4e-08 W=4e-07 
M7 Y C0 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI211_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 12 A0 Y VPW nch L=4e-08 W=2.3e-07 
M1 VSS A1 12 VPW nch L=4e-08 W=2.3e-07 
M2 Y B0 VSS VPW nch L=4e-08 W=1.5e-07 
M3 VSS C0 Y VPW nch L=4e-08 W=1.5e-07 
M4 VDD A1 1 VNW pch L=4e-08 W=2.85e-07 
M5 1 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M6 VDD A0 1 VNW pch L=4e-08 W=2.85e-07 
M7 1 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M8 9 B0 1 VNW pch L=4e-08 W=2.85e-07 
M9 Y C0 9 VNW pch L=4e-08 W=2.85e-07 
M10 10 C0 Y VNW pch L=4e-08 W=2.85e-07 
M11 1 B0 10 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI211_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 11 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M1 Y A0 11 VPW nch L=4e-08 W=1.6e-07 
M2 12 A0 Y VPW nch L=4e-08 W=1.6e-07 
M3 VSS A1 12 VPW nch L=4e-08 W=1.6e-07 
M4 Y B0 VSS VPW nch L=4e-08 W=2.1e-07 
M5 VSS C0 Y VPW nch L=4e-08 W=2.1e-07 
M6 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M7 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M8 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M9 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M10 9 B0 2 VNW pch L=4e-08 W=4e-07 
M11 Y C0 9 VNW pch L=4e-08 W=4e-07 
M12 10 C0 Y VNW pch L=4e-08 W=4e-07 
M13 2 B0 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI211_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 13 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M1 Y A0 13 VPW nch L=4e-08 W=2.4e-07 
M2 14 A0 Y VPW nch L=4e-08 W=2.4e-07 
M3 VSS A1 14 VPW nch L=4e-08 W=2.4e-07 
M4 Y B0 VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS C0 Y VPW nch L=4e-08 W=1.6e-07 
M6 Y C0 VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS B0 Y VPW nch L=4e-08 W=1.6e-07 
M8 VDD A0 1 VNW pch L=4e-08 W=4e-07 
M9 1 A1 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A1 1 VNW pch L=4e-08 W=4e-07 
M11 1 A0 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD A0 1 VNW pch L=4e-08 W=4e-07 
M13 1 A1 VDD VNW pch L=4e-08 W=4e-07 
M14 9 B0 1 VNW pch L=4e-08 W=4e-07 
M15 Y C0 9 VNW pch L=4e-08 W=4e-07 
M16 10 C0 Y VNW pch L=4e-08 W=4e-07 
M17 1 B0 10 VNW pch L=4e-08 W=4e-07 
M18 11 B0 1 VNW pch L=4e-08 W=4e-07 
M19 Y C0 11 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI211_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 13 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M1 Y A0 13 VPW nch L=4e-08 W=1.6e-07 
M2 14 A0 Y VPW nch L=4e-08 W=1.6e-07 
M3 VSS A1 14 VPW nch L=4e-08 W=1.6e-07 
M4 15 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M5 Y A0 15 VPW nch L=4e-08 W=1.6e-07 
M6 16 A0 Y VPW nch L=4e-08 W=1.6e-07 
M7 VSS A1 16 VPW nch L=4e-08 W=1.6e-07 
M8 Y B0 VSS VPW nch L=4e-08 W=2.1e-07 
M9 VSS C0 Y VPW nch L=4e-08 W=2.1e-07 
M10 Y C0 VSS VPW nch L=4e-08 W=2.1e-07 
M11 VSS B0 Y VPW nch L=4e-08 W=2.1e-07 
M12 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M13 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M15 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M17 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M19 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M20 9 B0 2 VNW pch L=4e-08 W=4e-07 
M21 Y C0 9 VNW pch L=4e-08 W=4e-07 
M22 10 C0 Y VNW pch L=4e-08 W=4e-07 
M23 2 B0 10 VNW pch L=4e-08 W=4e-07 
M24 11 B0 2 VNW pch L=4e-08 W=4e-07 
M25 Y C0 11 VNW pch L=4e-08 W=4e-07 
M26 12 C0 Y VNW pch L=4e-08 W=4e-07 
M27 2 B0 12 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21B_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 B0N VSS VPW nch L=4e-08 W=1.2e-07 
M1 9 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 Y A0 9 VPW nch L=4e-08 W=1.2e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=1.2e-07 
M4 3 B0N VDD VNW pch L=4e-08 W=1.55e-07 
M5 VDD A1 4 VNW pch L=4e-08 W=2e-07 
M6 4 A0 VDD VNW pch L=4e-08 W=2e-07 
M7 Y 3 4 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AOI21B_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 B0N VSS VPW nch L=4e-08 W=1.2e-07 
M1 9 A1 VSS VPW nch L=4e-08 W=1.8e-07 
M2 Y A0 9 VPW nch L=4e-08 W=1.8e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=1.2e-07 
M4 3 B0N VDD VNW pch L=4e-08 W=1.55e-07 
M5 VDD A1 4 VNW pch L=4e-08 W=3e-07 
M6 4 A0 VDD VNW pch L=4e-08 W=3e-07 
M7 Y 3 4 VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT AOI21B_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 B0N VSS VPW nch L=4e-08 W=1.2e-07 
M1 9 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M2 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M4 3 B0N VDD VNW pch L=4e-08 W=1.55e-07 
M5 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M6 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M7 Y 3 4 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21B_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 B0N VSS VPW nch L=4e-08 W=1.2e-07 
M1 9 A1 VSS VPW nch L=4e-08 W=1.7e-07 
M2 Y A0 9 VPW nch L=4e-08 W=1.7e-07 
M3 10 A0 Y VPW nch L=4e-08 W=1.7e-07 
M4 VSS A1 10 VPW nch L=4e-08 W=1.7e-07 
M5 Y 3 VSS VPW nch L=4e-08 W=2.3e-07 
M6 3 B0N VDD VNW pch L=4e-08 W=1.55e-07 
M7 VDD A1 4 VNW pch L=4e-08 W=2.85e-07 
M8 4 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M9 VDD A0 4 VNW pch L=4e-08 W=2.85e-07 
M10 4 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M11 Y 3 4 VNW pch L=4e-08 W=2.85e-07 
M12 4 3 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI21B_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 B0N VSS VPW nch L=4e-08 W=1.45e-07 
M1 9 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M2 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M3 10 A0 Y VPW nch L=4e-08 W=2.4e-07 
M4 VSS A1 10 VPW nch L=4e-08 W=2.4e-07 
M5 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M6 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M7 3 B0N VDD VNW pch L=4e-08 W=1.9e-07 
M8 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M9 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M11 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M12 Y 3 4 VNW pch L=4e-08 W=4e-07 
M13 4 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21B_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 B0N VSS VPW nch L=4e-08 W=2.15e-07 
M1 Y 3 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS 3 Y VPW nch L=4e-08 W=2.4e-07 
M3 10 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M4 Y A0 10 VPW nch L=4e-08 W=3.6e-07 
M5 11 A0 Y VPW nch L=4e-08 W=3.6e-07 
M6 VSS A1 11 VPW nch L=4e-08 W=3.6e-07 
M7 3 B0N VDD VNW pch L=4e-08 W=2.75e-07 
M8 5 3 Y VNW pch L=4e-08 W=4e-07 
M9 Y 3 5 VNW pch L=4e-08 W=4e-07 
M10 5 3 Y VNW pch L=4e-08 W=4e-07 
M11 VDD A1 5 VNW pch L=4e-08 W=4e-07 
M12 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M13 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M14 5 A1 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD A1 5 VNW pch L=4e-08 W=4e-07 
M16 5 A0 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21B_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 B0N VSS VPW nch L=4e-08 W=2.8e-07 
M1 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M3 10 A0 Y VPW nch L=4e-08 W=3.2e-07 
M4 VSS A1 10 VPW nch L=4e-08 W=3.2e-07 
M5 11 A1 VSS VPW nch L=4e-08 W=3.2e-07 
M6 Y A0 11 VPW nch L=4e-08 W=3.2e-07 
M7 12 A0 Y VPW nch L=4e-08 W=3.2e-07 
M8 VSS A1 12 VPW nch L=4e-08 W=3.2e-07 
M9 3 B0N VDD VNW pch L=4e-08 W=3.6e-07 
M10 Y 3 4 VNW pch L=4e-08 W=4e-07 
M11 4 3 Y VNW pch L=4e-08 W=4e-07 
M12 Y 3 4 VNW pch L=4e-08 W=4e-07 
M13 4 3 Y VNW pch L=4e-08 W=4e-07 
M14 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M15 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M17 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M19 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M21 4 A0 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21B_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 B0N VSS VPW nch L=4e-08 W=2.1e-07 
M1 VSS B0N 3 VPW nch L=4e-08 W=2.1e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M5 10 A0 Y VPW nch L=4e-08 W=3.6e-07 
M6 VSS A1 10 VPW nch L=4e-08 W=3.6e-07 
M7 11 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M8 Y A0 11 VPW nch L=4e-08 W=3.6e-07 
M9 12 A0 Y VPW nch L=4e-08 W=3.6e-07 
M10 VSS A1 12 VPW nch L=4e-08 W=3.6e-07 
M11 13 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M12 Y A0 13 VPW nch L=4e-08 W=3.6e-07 
M13 3 B0N VDD VNW pch L=4e-08 W=2.75e-07 
M14 VDD B0N 3 VNW pch L=4e-08 W=2.75e-07 
M15 Y 3 4 VNW pch L=4e-08 W=4e-07 
M16 4 3 Y VNW pch L=4e-08 W=4e-07 
M17 Y 3 4 VNW pch L=4e-08 W=4e-07 
M18 4 3 Y VNW pch L=4e-08 W=4e-07 
M19 Y 3 4 VNW pch L=4e-08 W=4e-07 
M20 4 3 Y VNW pch L=4e-08 W=4e-07 
M21 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M22 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M24 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M26 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M28 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M30 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M32 4 A0 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21B_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 B0N VSS VPW nch L=4e-08 W=2.8e-07 
M1 VSS B0N 3 VPW nch L=4e-08 W=2.8e-07 
M2 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M3 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M4 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M5 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M6 10 A0 Y VPW nch L=4e-08 W=3.2e-07 
M7 VSS A1 10 VPW nch L=4e-08 W=3.2e-07 
M8 11 A1 VSS VPW nch L=4e-08 W=3.2e-07 
M9 Y A0 11 VPW nch L=4e-08 W=3.2e-07 
M10 12 A0 Y VPW nch L=4e-08 W=3.2e-07 
M11 VSS A1 12 VPW nch L=4e-08 W=3.2e-07 
M12 13 A1 VSS VPW nch L=4e-08 W=3.2e-07 
M13 Y A0 13 VPW nch L=4e-08 W=3.2e-07 
M14 14 A0 Y VPW nch L=4e-08 W=3.2e-07 
M15 VSS A1 14 VPW nch L=4e-08 W=3.2e-07 
M16 15 A1 VSS VPW nch L=4e-08 W=3.2e-07 
M17 Y A0 15 VPW nch L=4e-08 W=3.2e-07 
M18 3 B0N VDD VNW pch L=4e-08 W=3.6e-07 
M19 VDD B0N 3 VNW pch L=4e-08 W=3.6e-07 
M20 Y 3 4 VNW pch L=4e-08 W=4e-07 
M21 4 3 Y VNW pch L=4e-08 W=4e-07 
M22 Y 3 4 VNW pch L=4e-08 W=4e-07 
M23 4 3 Y VNW pch L=4e-08 W=4e-07 
M24 Y 3 4 VNW pch L=4e-08 W=4e-07 
M25 4 3 Y VNW pch L=4e-08 W=4e-07 
M26 Y 3 4 VNW pch L=4e-08 W=4e-07 
M27 4 3 Y VNW pch L=4e-08 W=4e-07 
M28 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M29 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M31 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M33 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M35 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M37 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M39 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M41 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M42 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M43 4 A0 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 8 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A0 8 VPW nch L=4e-08 W=1.2e-07 
M2 VSS B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 VDD A1 2 VNW pch L=4e-08 W=2e-07 
M4 2 A0 VDD VNW pch L=4e-08 W=2e-07 
M5 Y B0 2 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AOI21_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 8 A1 VSS VPW nch L=4e-08 W=1.8e-07 
M1 Y A0 8 VPW nch L=4e-08 W=1.8e-07 
M2 VSS B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 VDD A1 2 VNW pch L=4e-08 W=3e-07 
M4 2 A0 VDD VNW pch L=4e-08 W=3e-07 
M5 Y B0 2 VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT AOI21_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 8 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M1 Y A0 8 VPW nch L=4e-08 W=2.4e-07 
M2 VSS B0 Y VPW nch L=4e-08 W=1.6e-07 
M3 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M4 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M5 Y B0 2 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 9 A1 VSS VPW nch L=4e-08 W=3.4e-07 
M1 Y A0 9 VPW nch L=4e-08 W=3.4e-07 
M2 VSS B0 Y VPW nch L=4e-08 W=2.3e-07 
M3 VDD A0 1 VNW pch L=4e-08 W=2.85e-07 
M4 1 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M5 VDD A1 1 VNW pch L=4e-08 W=2.85e-07 
M6 1 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M7 Y B0 1 VNW pch L=4e-08 W=2.85e-07 
M8 1 B0 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI21_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 8 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M1 Y A0 8 VPW nch L=4e-08 W=2.4e-07 
M2 9 A0 Y VPW nch L=4e-08 W=2.4e-07 
M3 VSS A1 9 VPW nch L=4e-08 W=2.4e-07 
M4 Y B0 VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS B0 Y VPW nch L=4e-08 W=1.6e-07 
M6 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M7 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M8 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M9 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M10 Y B0 2 VNW pch L=4e-08 W=4e-07 
M11 2 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 8 A0 Y VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=2.4e-07 
M2 9 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M4 10 A0 Y VPW nch L=4e-08 W=2.4e-07 
M5 VSS A1 10 VPW nch L=4e-08 W=2.4e-07 
M6 Y B0 VSS VPW nch L=4e-08 W=2.4e-07 
M7 VSS B0 Y VPW nch L=4e-08 W=2.4e-07 
M8 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M9 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M11 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M13 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M14 Y B0 2 VNW pch L=4e-08 W=4e-07 
M15 2 B0 Y VNW pch L=4e-08 W=4e-07 
M16 Y B0 2 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 8 A0 Y VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=2.4e-07 
M2 9 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M4 10 A0 Y VPW nch L=4e-08 W=2.4e-07 
M5 VSS A1 10 VPW nch L=4e-08 W=2.4e-07 
M6 11 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M7 Y A0 11 VPW nch L=4e-08 W=2.4e-07 
M8 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M9 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M10 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M11 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M13 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M15 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M17 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M18 Y B0 2 VNW pch L=4e-08 W=4e-07 
M19 2 B0 Y VNW pch L=4e-08 W=4e-07 
M20 Y B0 2 VNW pch L=4e-08 W=4e-07 
M21 2 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 8 A0 Y VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=2.4e-07 
M2 9 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M4 10 A0 Y VPW nch L=4e-08 W=2.4e-07 
M5 VSS A1 10 VPW nch L=4e-08 W=2.4e-07 
M6 11 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M7 Y A0 11 VPW nch L=4e-08 W=2.4e-07 
M8 12 A0 Y VPW nch L=4e-08 W=2.4e-07 
M9 VSS A1 12 VPW nch L=4e-08 W=2.4e-07 
M10 13 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M11 Y A0 13 VPW nch L=4e-08 W=2.4e-07 
M12 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M13 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M14 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M15 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M16 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M17 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M18 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M20 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M22 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M24 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M26 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M27 Y B0 2 VNW pch L=4e-08 W=4e-07 
M28 2 B0 Y VNW pch L=4e-08 W=4e-07 
M29 Y B0 2 VNW pch L=4e-08 W=4e-07 
M30 2 B0 Y VNW pch L=4e-08 W=4e-07 
M31 Y B0 2 VNW pch L=4e-08 W=4e-07 
M32 2 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI21_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 8 A0 Y VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1 8 VPW nch L=4e-08 W=2.4e-07 
M2 9 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M4 10 A0 Y VPW nch L=4e-08 W=2.4e-07 
M5 VSS A1 10 VPW nch L=4e-08 W=2.4e-07 
M6 11 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M7 Y A0 11 VPW nch L=4e-08 W=2.4e-07 
M8 12 A0 Y VPW nch L=4e-08 W=2.4e-07 
M9 VSS A1 12 VPW nch L=4e-08 W=2.4e-07 
M10 13 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M11 Y A0 13 VPW nch L=4e-08 W=2.4e-07 
M12 14 A0 Y VPW nch L=4e-08 W=2.4e-07 
M13 VSS A1 14 VPW nch L=4e-08 W=2.4e-07 
M14 15 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M15 Y A0 15 VPW nch L=4e-08 W=2.4e-07 
M16 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M17 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M18 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M19 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M20 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M21 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M23 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M25 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M27 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M29 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M31 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M33 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M35 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M36 Y B0 2 VNW pch L=4e-08 W=4e-07 
M37 2 B0 Y VNW pch L=4e-08 W=4e-07 
M38 Y B0 2 VNW pch L=4e-08 W=4e-07 
M39 2 B0 Y VNW pch L=4e-08 W=4e-07 
M40 Y B0 2 VNW pch L=4e-08 W=4e-07 
M41 2 B0 Y VNW pch L=4e-08 W=4e-07 
M42 Y B0 2 VNW pch L=4e-08 W=4e-07 
M43 2 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI221_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 11 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A0 11 VPW nch L=4e-08 W=1.2e-07 
M2 12 B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 VSS B1 12 VPW nch L=4e-08 W=1.2e-07 
M4 Y C0 VSS VPW nch L=4e-08 W=1.2e-07 
M5 VDD A1 2 VNW pch L=4e-08 W=2.1e-07 
M6 2 A0 VDD VNW pch L=4e-08 W=2.1e-07 
M7 5 B0 2 VNW pch L=4e-08 W=2.1e-07 
M8 2 B1 5 VNW pch L=4e-08 W=2.1e-07 
M9 Y C0 5 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AOI221_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 11 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A0 11 VPW nch L=4e-08 W=1.2e-07 
M2 12 B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 VSS B1 12 VPW nch L=4e-08 W=1.2e-07 
M4 Y C0 VSS VPW nch L=4e-08 W=1.2e-07 
M5 VDD A1 2 VNW pch L=4e-08 W=2.85e-07 
M6 2 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M7 5 B0 2 VNW pch L=4e-08 W=2.85e-07 
M8 2 B1 5 VNW pch L=4e-08 W=2.85e-07 
M9 Y C0 5 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI221_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 11 A1 VSS VPW nch L=4e-08 W=1.8e-07 
M1 Y A0 11 VPW nch L=4e-08 W=1.8e-07 
M2 12 B0 Y VPW nch L=4e-08 W=1.8e-07 
M3 VSS B1 12 VPW nch L=4e-08 W=1.8e-07 
M4 Y C0 VSS VPW nch L=4e-08 W=1.2e-07 
M5 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M6 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M7 5 B0 2 VNW pch L=4e-08 W=4e-07 
M8 2 B1 5 VNW pch L=4e-08 W=4e-07 
M9 Y C0 5 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI221_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 12 A1 VSS VPW nch L=4e-08 W=2.3e-07 
M1 Y A0 12 VPW nch L=4e-08 W=2.3e-07 
M2 13 B0 Y VPW nch L=4e-08 W=2.3e-07 
M3 VSS B1 13 VPW nch L=4e-08 W=2.3e-07 
M4 Y C0 VSS VPW nch L=4e-08 W=1.5e-07 
M5 VDD A0 1 VNW pch L=4e-08 W=2.85e-07 
M6 1 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M7 VDD A1 1 VNW pch L=4e-08 W=2.85e-07 
M8 1 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M9 5 B0 1 VNW pch L=4e-08 W=2.85e-07 
M10 1 B1 5 VNW pch L=4e-08 W=2.85e-07 
M11 5 B1 1 VNW pch L=4e-08 W=2.85e-07 
M12 1 B0 5 VNW pch L=4e-08 W=2.85e-07 
M13 Y C0 5 VNW pch L=4e-08 W=2.85e-07 
M14 5 C0 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI221_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 11 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M1 Y A0 11 VPW nch L=4e-08 W=1.6e-07 
M2 12 A0 Y VPW nch L=4e-08 W=1.6e-07 
M3 VSS A1 12 VPW nch L=4e-08 W=1.6e-07 
M4 13 B1 VSS VPW nch L=4e-08 W=1.6e-07 
M5 Y B0 13 VPW nch L=4e-08 W=1.6e-07 
M6 14 B0 Y VPW nch L=4e-08 W=1.6e-07 
M7 VSS B1 14 VPW nch L=4e-08 W=1.6e-07 
M8 Y C0 VSS VPW nch L=4e-08 W=2.1e-07 
M9 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M10 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M12 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 5 B1 2 VNW pch L=4e-08 W=4e-07 
M14 2 B0 5 VNW pch L=4e-08 W=4e-07 
M15 5 B0 2 VNW pch L=4e-08 W=4e-07 
M16 2 B1 5 VNW pch L=4e-08 W=4e-07 
M17 Y C0 5 VNW pch L=4e-08 W=4e-07 
M18 5 C0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI221_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 12 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M1 Y A0 12 VPW nch L=4e-08 W=2.4e-07 
M2 13 A0 Y VPW nch L=4e-08 W=2.4e-07 
M3 VSS A1 13 VPW nch L=4e-08 W=2.4e-07 
M4 14 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M5 Y B0 14 VPW nch L=4e-08 W=2.4e-07 
M6 15 B0 Y VPW nch L=4e-08 W=2.4e-07 
M7 VSS B1 15 VPW nch L=4e-08 W=2.4e-07 
M8 Y C0 VSS VPW nch L=4e-08 W=3.15e-07 
M9 VDD A0 1 VNW pch L=4e-08 W=4e-07 
M10 1 A1 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD A1 1 VNW pch L=4e-08 W=4e-07 
M12 1 A0 VDD VNW pch L=4e-08 W=4e-07 
M13 VDD A0 1 VNW pch L=4e-08 W=4e-07 
M14 1 A1 VDD VNW pch L=4e-08 W=4e-07 
M15 5 B1 1 VNW pch L=4e-08 W=4e-07 
M16 1 B0 5 VNW pch L=4e-08 W=4e-07 
M17 5 B0 1 VNW pch L=4e-08 W=4e-07 
M18 1 B1 5 VNW pch L=4e-08 W=4e-07 
M19 5 B1 1 VNW pch L=4e-08 W=4e-07 
M20 1 B0 5 VNW pch L=4e-08 W=4e-07 
M21 Y C0 5 VNW pch L=4e-08 W=4e-07 
M22 5 C0 Y VNW pch L=4e-08 W=4e-07 
M23 Y C0 5 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI221_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 11 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M1 Y A0 11 VPW nch L=4e-08 W=1.6e-07 
M2 12 A0 Y VPW nch L=4e-08 W=1.6e-07 
M3 VSS A1 12 VPW nch L=4e-08 W=1.6e-07 
M4 13 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M5 Y A0 13 VPW nch L=4e-08 W=1.6e-07 
M6 14 A0 Y VPW nch L=4e-08 W=1.6e-07 
M7 VSS A1 14 VPW nch L=4e-08 W=1.6e-07 
M8 15 B1 VSS VPW nch L=4e-08 W=1.6e-07 
M9 Y B0 15 VPW nch L=4e-08 W=1.6e-07 
M10 16 B0 Y VPW nch L=4e-08 W=1.6e-07 
M11 VSS B1 16 VPW nch L=4e-08 W=1.6e-07 
M12 17 B1 VSS VPW nch L=4e-08 W=1.6e-07 
M13 Y B0 17 VPW nch L=4e-08 W=1.6e-07 
M14 18 B0 Y VPW nch L=4e-08 W=1.6e-07 
M15 VSS B1 18 VPW nch L=4e-08 W=1.6e-07 
M16 Y C0 VSS VPW nch L=4e-08 W=2.1e-07 
M17 VSS C0 Y VPW nch L=4e-08 W=2.1e-07 
M18 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M19 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M21 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M23 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M25 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M26 5 B1 2 VNW pch L=4e-08 W=4e-07 
M27 2 B0 5 VNW pch L=4e-08 W=4e-07 
M28 5 B0 2 VNW pch L=4e-08 W=4e-07 
M29 2 B1 5 VNW pch L=4e-08 W=4e-07 
M30 5 B1 2 VNW pch L=4e-08 W=4e-07 
M31 2 B0 5 VNW pch L=4e-08 W=4e-07 
M32 5 B0 2 VNW pch L=4e-08 W=4e-07 
M33 2 B1 5 VNW pch L=4e-08 W=4e-07 
M34 Y C0 5 VNW pch L=4e-08 W=4e-07 
M35 5 C0 Y VNW pch L=4e-08 W=4e-07 
M36 Y C0 5 VNW pch L=4e-08 W=4e-07 
M37 5 C0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI222_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 12 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A0 12 VPW nch L=4e-08 W=1.2e-07 
M2 13 B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 VSS B1 13 VPW nch L=4e-08 W=1.2e-07 
M4 14 C0 Y VPW nch L=4e-08 W=1.2e-07 
M5 VSS C1 14 VPW nch L=4e-08 W=1.2e-07 
M6 VDD A1 2 VNW pch L=4e-08 W=2.1e-07 
M7 2 A0 VDD VNW pch L=4e-08 W=2.1e-07 
M8 5 B0 2 VNW pch L=4e-08 W=2.1e-07 
M9 2 B1 5 VNW pch L=4e-08 W=2.1e-07 
M10 Y C0 5 VNW pch L=4e-08 W=2.1e-07 
M11 5 C1 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT AOI222_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 12 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A0 12 VPW nch L=4e-08 W=1.2e-07 
M2 13 B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 VSS B1 13 VPW nch L=4e-08 W=1.2e-07 
M4 14 C0 Y VPW nch L=4e-08 W=1.2e-07 
M5 VSS C1 14 VPW nch L=4e-08 W=1.2e-07 
M6 VDD A1 2 VNW pch L=4e-08 W=2.95e-07 
M7 2 A0 VDD VNW pch L=4e-08 W=2.95e-07 
M8 5 B0 2 VNW pch L=4e-08 W=2.95e-07 
M9 2 B1 5 VNW pch L=4e-08 W=2.95e-07 
M10 Y C0 5 VNW pch L=4e-08 W=2.95e-07 
M11 5 C1 Y VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT AOI222_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 12 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M1 Y A0 12 VPW nch L=4e-08 W=1.6e-07 
M2 13 B0 Y VPW nch L=4e-08 W=1.6e-07 
M3 VSS B1 13 VPW nch L=4e-08 W=1.6e-07 
M4 14 C0 Y VPW nch L=4e-08 W=1.6e-07 
M5 VSS C1 14 VPW nch L=4e-08 W=1.6e-07 
M6 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M7 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M8 5 B0 2 VNW pch L=4e-08 W=4e-07 
M9 2 B1 5 VNW pch L=4e-08 W=4e-07 
M10 Y C0 5 VNW pch L=4e-08 W=4e-07 
M11 5 C1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI222_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 13 A1 VSS VPW nch L=4e-08 W=2.3e-07 
M1 Y A0 13 VPW nch L=4e-08 W=2.3e-07 
M2 14 B0 Y VPW nch L=4e-08 W=2.3e-07 
M3 VSS B1 14 VPW nch L=4e-08 W=2.3e-07 
M4 16 C1 VSS VPW nch L=4e-08 W=2.3e-07 
M5 Y C0 16 VPW nch L=4e-08 W=2.3e-07 
M6 VDD A0 1 VNW pch L=4e-08 W=2.85e-07 
M7 1 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M8 VDD A1 1 VNW pch L=4e-08 W=2.85e-07 
M9 1 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M10 5 B0 1 VNW pch L=4e-08 W=2.85e-07 
M11 1 B1 5 VNW pch L=4e-08 W=2.85e-07 
M12 5 B1 1 VNW pch L=4e-08 W=2.85e-07 
M13 1 B0 5 VNW pch L=4e-08 W=2.85e-07 
M14 Y C1 5 VNW pch L=4e-08 W=2.85e-07 
M15 5 C0 Y VNW pch L=4e-08 W=2.85e-07 
M16 Y C0 5 VNW pch L=4e-08 W=2.85e-07 
M17 5 C1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI222_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 12 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M1 Y A0 12 VPW nch L=4e-08 W=1.6e-07 
M2 13 A0 Y VPW nch L=4e-08 W=1.6e-07 
M3 VSS A1 13 VPW nch L=4e-08 W=1.6e-07 
M4 14 B1 VSS VPW nch L=4e-08 W=1.6e-07 
M5 Y B0 14 VPW nch L=4e-08 W=1.6e-07 
M6 15 B0 Y VPW nch L=4e-08 W=1.6e-07 
M7 VSS B1 15 VPW nch L=4e-08 W=1.6e-07 
M8 16 C1 VSS VPW nch L=4e-08 W=1.6e-07 
M9 Y C0 16 VPW nch L=4e-08 W=1.6e-07 
M10 17 C0 Y VPW nch L=4e-08 W=1.6e-07 
M11 VSS C1 17 VPW nch L=4e-08 W=1.6e-07 
M12 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M13 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M15 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M16 5 B1 2 VNW pch L=4e-08 W=4e-07 
M17 2 B0 5 VNW pch L=4e-08 W=4e-07 
M18 5 B0 2 VNW pch L=4e-08 W=4e-07 
M19 2 B1 5 VNW pch L=4e-08 W=4e-07 
M20 Y C1 5 VNW pch L=4e-08 W=4e-07 
M21 5 C0 Y VNW pch L=4e-08 W=4e-07 
M22 Y C0 5 VNW pch L=4e-08 W=4e-07 
M23 5 C1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI222_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 12 A0 Y VPW nch L=4e-08 W=1.6e-07 
M1 VSS A1 12 VPW nch L=4e-08 W=1.6e-07 
M2 13 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M3 Y A0 13 VPW nch L=4e-08 W=1.6e-07 
M4 14 A0 Y VPW nch L=4e-08 W=1.6e-07 
M5 VSS A1 14 VPW nch L=4e-08 W=1.6e-07 
M6 15 B1 VSS VPW nch L=4e-08 W=1.6e-07 
M7 Y B0 15 VPW nch L=4e-08 W=1.6e-07 
M8 16 B0 Y VPW nch L=4e-08 W=1.6e-07 
M9 VSS B1 16 VPW nch L=4e-08 W=1.6e-07 
M10 17 B1 VSS VPW nch L=4e-08 W=1.6e-07 
M11 Y B0 17 VPW nch L=4e-08 W=1.6e-07 
M12 18 C1 VSS VPW nch L=4e-08 W=1.6e-07 
M13 Y C0 18 VPW nch L=4e-08 W=1.6e-07 
M14 19 C0 Y VPW nch L=4e-08 W=1.6e-07 
M15 VSS C1 19 VPW nch L=4e-08 W=1.6e-07 
M16 20 C1 VSS VPW nch L=4e-08 W=1.6e-07 
M17 Y C0 20 VPW nch L=4e-08 W=1.6e-07 
M18 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M19 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M21 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M23 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M24 5 B1 2 VNW pch L=4e-08 W=4e-07 
M25 2 B0 5 VNW pch L=4e-08 W=4e-07 
M26 5 B0 2 VNW pch L=4e-08 W=4e-07 
M27 2 B1 5 VNW pch L=4e-08 W=4e-07 
M28 5 B1 2 VNW pch L=4e-08 W=4e-07 
M29 2 B0 5 VNW pch L=4e-08 W=4e-07 
M30 Y C1 5 VNW pch L=4e-08 W=4e-07 
M31 5 C0 Y VNW pch L=4e-08 W=4e-07 
M32 Y C0 5 VNW pch L=4e-08 W=4e-07 
M33 5 C1 Y VNW pch L=4e-08 W=4e-07 
M34 Y C1 5 VNW pch L=4e-08 W=4e-07 
M35 5 C0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI222_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 12 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M1 Y A0 12 VPW nch L=4e-08 W=1.6e-07 
M2 13 A0 Y VPW nch L=4e-08 W=1.6e-07 
M3 VSS A1 13 VPW nch L=4e-08 W=1.6e-07 
M4 14 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M5 Y A0 14 VPW nch L=4e-08 W=1.6e-07 
M6 15 A0 Y VPW nch L=4e-08 W=1.6e-07 
M7 VSS A1 15 VPW nch L=4e-08 W=1.6e-07 
M8 16 B1 VSS VPW nch L=4e-08 W=1.6e-07 
M9 Y B0 16 VPW nch L=4e-08 W=1.6e-07 
M10 17 B0 Y VPW nch L=4e-08 W=1.6e-07 
M11 VSS B1 17 VPW nch L=4e-08 W=1.6e-07 
M12 18 B1 VSS VPW nch L=4e-08 W=1.6e-07 
M13 Y B0 18 VPW nch L=4e-08 W=1.6e-07 
M14 19 B0 Y VPW nch L=4e-08 W=1.6e-07 
M15 VSS B1 19 VPW nch L=4e-08 W=1.6e-07 
M16 20 C1 VSS VPW nch L=4e-08 W=1.6e-07 
M17 Y C0 20 VPW nch L=4e-08 W=1.6e-07 
M18 21 C0 Y VPW nch L=4e-08 W=1.6e-07 
M19 VSS C1 21 VPW nch L=4e-08 W=1.6e-07 
M20 22 C1 VSS VPW nch L=4e-08 W=1.6e-07 
M21 Y C0 22 VPW nch L=4e-08 W=1.6e-07 
M22 23 C0 Y VPW nch L=4e-08 W=1.6e-07 
M23 VSS C1 23 VPW nch L=4e-08 W=1.6e-07 
M24 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M25 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M27 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M29 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M31 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M32 5 B1 2 VNW pch L=4e-08 W=4e-07 
M33 2 B0 5 VNW pch L=4e-08 W=4e-07 
M34 5 B0 2 VNW pch L=4e-08 W=4e-07 
M35 2 B1 5 VNW pch L=4e-08 W=4e-07 
M36 5 B1 2 VNW pch L=4e-08 W=4e-07 
M37 2 B0 5 VNW pch L=4e-08 W=4e-07 
M38 5 B0 2 VNW pch L=4e-08 W=4e-07 
M39 2 B1 5 VNW pch L=4e-08 W=4e-07 
M40 Y C1 5 VNW pch L=4e-08 W=4e-07 
M41 5 C0 Y VNW pch L=4e-08 W=4e-07 
M42 Y C0 5 VNW pch L=4e-08 W=4e-07 
M43 5 C1 Y VNW pch L=4e-08 W=4e-07 
M44 Y C1 5 VNW pch L=4e-08 W=4e-07 
M45 5 C0 Y VNW pch L=4e-08 W=4e-07 
M46 Y C0 5 VNW pch L=4e-08 W=4e-07 
M47 5 C1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22BB_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 3 B1N VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B0N 3 VPW nch L=4e-08 W=1.2e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M3 Y A0 11 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 3 Y VPW nch L=4e-08 W=1.2e-07 
M5 10 B1N VDD VNW pch L=4e-08 W=2e-07 
M6 3 B0N 10 VNW pch L=4e-08 W=2e-07 
M7 VDD A1 4 VNW pch L=4e-08 W=2e-07 
M8 4 A0 VDD VNW pch L=4e-08 W=2e-07 
M9 Y 3 4 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AOI22BB_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 3 B1N VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B0N 3 VPW nch L=4e-08 W=1.2e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=1.8e-07 
M3 Y A0 11 VPW nch L=4e-08 W=1.8e-07 
M4 VSS 3 Y VPW nch L=4e-08 W=1.2e-07 
M5 10 B1N VDD VNW pch L=4e-08 W=2.3e-07 
M6 3 B0N 10 VNW pch L=4e-08 W=2.3e-07 
M7 VDD A1 4 VNW pch L=4e-08 W=3e-07 
M8 4 A0 VDD VNW pch L=4e-08 W=3e-07 
M9 Y 3 4 VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT AOI22BB_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 3 B1N VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B0N 3 VPW nch L=4e-08 W=1.2e-07 
M2 11 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y A0 11 VPW nch L=4e-08 W=2.4e-07 
M4 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M5 10 B1N VDD VNW pch L=4e-08 W=2.7e-07 
M6 3 B0N 10 VNW pch L=4e-08 W=2.7e-07 
M7 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M8 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M9 Y 3 4 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22BB_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 3 B1N VSS VPW nch L=4e-08 W=1.4e-07 
M1 VSS B0N 3 VPW nch L=4e-08 W=1.4e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=2.3e-07 
M3 12 A0 Y VPW nch L=4e-08 W=3.4e-07 
M4 VSS A1 12 VPW nch L=4e-08 W=3.4e-07 
M5 10 B1N VDD VNW pch L=4e-08 W=3.55e-07 
M6 3 B0N 10 VNW pch L=4e-08 W=3.55e-07 
M7 Y 3 4 VNW pch L=4e-08 W=2.85e-07 
M8 4 3 Y VNW pch L=4e-08 W=2.85e-07 
M9 VDD A0 4 VNW pch L=4e-08 W=2.85e-07 
M10 4 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M11 VDD A1 4 VNW pch L=4e-08 W=2.85e-07 
M12 4 A0 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI22BB_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 3 B1N VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS B0N 3 VPW nch L=4e-08 W=1.6e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M4 11 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M5 Y A0 11 VPW nch L=4e-08 W=2.4e-07 
M6 12 A0 Y VPW nch L=4e-08 W=2.4e-07 
M7 VSS A1 12 VPW nch L=4e-08 W=2.4e-07 
M8 10 B1N VDD VNW pch L=4e-08 W=4e-07 
M9 3 B0N 10 VNW pch L=4e-08 W=4e-07 
M10 Y 3 4 VNW pch L=4e-08 W=4e-07 
M11 4 3 Y VNW pch L=4e-08 W=4e-07 
M12 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M13 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M15 4 A1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22BB_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 3 B0N VSS VPW nch L=4e-08 W=2.8e-07 
M1 VSS B1N 3 VPW nch L=4e-08 W=2.8e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=2.4e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=2.4e-07 
M4 14 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M5 Y A0 14 VPW nch L=4e-08 W=2.4e-07 
M6 15 A0 Y VPW nch L=4e-08 W=2.4e-07 
M7 VSS A1 15 VPW nch L=4e-08 W=2.4e-07 
M8 16 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M9 Y A0 16 VPW nch L=4e-08 W=2.4e-07 
M10 10 B1N VDD VNW pch L=4e-08 W=3.5e-07 
M11 3 B0N 10 VNW pch L=4e-08 W=3.5e-07 
M12 11 B0N 3 VNW pch L=4e-08 W=3.5e-07 
M13 VDD B1N 11 VNW pch L=4e-08 W=3.5e-07 
M14 5 3 Y VNW pch L=4e-08 W=4e-07 
M15 Y 3 5 VNW pch L=4e-08 W=4e-07 
M16 5 3 Y VNW pch L=4e-08 W=4e-07 
M17 VDD A1 5 VNW pch L=4e-08 W=4e-07 
M18 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M20 5 A1 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A1 5 VNW pch L=4e-08 W=4e-07 
M22 5 A0 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22BB_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 3 B0N VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS B1N 3 VPW nch L=4e-08 W=3.2e-07 
M2 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M3 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M4 14 A0 Y VPW nch L=4e-08 W=2.4e-07 
M5 VSS A1 14 VPW nch L=4e-08 W=2.4e-07 
M6 15 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M7 Y A0 15 VPW nch L=4e-08 W=2.4e-07 
M8 16 A0 Y VPW nch L=4e-08 W=2.4e-07 
M9 VSS A1 16 VPW nch L=4e-08 W=2.4e-07 
M10 17 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M11 Y A0 17 VPW nch L=4e-08 W=2.4e-07 
M12 10 B1N VDD VNW pch L=4e-08 W=4e-07 
M13 3 B0N 10 VNW pch L=4e-08 W=4e-07 
M14 11 B0N 3 VNW pch L=4e-08 W=4e-07 
M15 VDD B1N 11 VNW pch L=4e-08 W=4e-07 
M16 Y 3 4 VNW pch L=4e-08 W=4e-07 
M17 4 3 Y VNW pch L=4e-08 W=4e-07 
M18 Y 3 4 VNW pch L=4e-08 W=4e-07 
M19 4 3 Y VNW pch L=4e-08 W=4e-07 
M20 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M21 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M23 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M25 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M27 4 A0 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22BB_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 3 B0N VSS VPW nch L=4e-08 W=2.4e-07 
M1 VSS B1N 3 VPW nch L=4e-08 W=2.4e-07 
M2 3 B1N VSS VPW nch L=4e-08 W=2.4e-07 
M3 VSS B0N 3 VPW nch L=4e-08 W=2.4e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M7 15 A0 Y VPW nch L=4e-08 W=2.4e-07 
M8 VSS A1 15 VPW nch L=4e-08 W=2.4e-07 
M9 16 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M10 Y A0 16 VPW nch L=4e-08 W=2.4e-07 
M11 17 A0 Y VPW nch L=4e-08 W=2.4e-07 
M12 VSS A1 17 VPW nch L=4e-08 W=2.4e-07 
M13 18 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M14 Y A0 18 VPW nch L=4e-08 W=2.4e-07 
M15 19 A0 Y VPW nch L=4e-08 W=2.4e-07 
M16 VSS A1 19 VPW nch L=4e-08 W=2.4e-07 
M17 20 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M18 Y A0 20 VPW nch L=4e-08 W=2.4e-07 
M19 10 B1N VDD VNW pch L=4e-08 W=4e-07 
M20 3 B0N 10 VNW pch L=4e-08 W=4e-07 
M21 11 B0N 3 VNW pch L=4e-08 W=4e-07 
M22 VDD B1N 11 VNW pch L=4e-08 W=4e-07 
M23 12 B1N VDD VNW pch L=4e-08 W=4e-07 
M24 3 B0N 12 VNW pch L=4e-08 W=4e-07 
M25 Y 3 4 VNW pch L=4e-08 W=4e-07 
M26 4 3 Y VNW pch L=4e-08 W=4e-07 
M27 Y 3 4 VNW pch L=4e-08 W=4e-07 
M28 4 3 Y VNW pch L=4e-08 W=4e-07 
M29 Y 3 4 VNW pch L=4e-08 W=4e-07 
M30 4 3 Y VNW pch L=4e-08 W=4e-07 
M31 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M32 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M33 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M34 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M36 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M38 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M40 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M41 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M42 4 A0 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22BB_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 2 B1N VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS B0N 2 VPW nch L=4e-08 W=3.2e-07 
M2 2 B0N VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS B1N 2 VPW nch L=4e-08 W=3.2e-07 
M4 VSS 2 Y VPW nch L=4e-08 W=3.2e-07 
M5 Y 2 VSS VPW nch L=4e-08 W=3.2e-07 
M6 VSS 2 Y VPW nch L=4e-08 W=3.2e-07 
M7 Y 2 VSS VPW nch L=4e-08 W=3.2e-07 
M8 16 A0 Y VPW nch L=4e-08 W=2.4e-07 
M9 VSS A1 16 VPW nch L=4e-08 W=2.4e-07 
M10 17 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M11 Y A0 17 VPW nch L=4e-08 W=2.4e-07 
M12 18 A0 Y VPW nch L=4e-08 W=2.4e-07 
M13 VSS A1 18 VPW nch L=4e-08 W=2.4e-07 
M14 19 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M15 Y A0 19 VPW nch L=4e-08 W=2.4e-07 
M16 20 A0 Y VPW nch L=4e-08 W=2.4e-07 
M17 VSS A1 20 VPW nch L=4e-08 W=2.4e-07 
M18 21 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M19 Y A0 21 VPW nch L=4e-08 W=2.4e-07 
M20 22 A0 Y VPW nch L=4e-08 W=2.4e-07 
M21 VSS A1 22 VPW nch L=4e-08 W=2.4e-07 
M22 23 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M23 Y A0 23 VPW nch L=4e-08 W=2.4e-07 
M24 10 B1N VDD VNW pch L=4e-08 W=4e-07 
M25 2 B0N 10 VNW pch L=4e-08 W=4e-07 
M26 11 B0N 2 VNW pch L=4e-08 W=4e-07 
M27 VDD B1N 11 VNW pch L=4e-08 W=4e-07 
M28 12 B1N VDD VNW pch L=4e-08 W=4e-07 
M29 2 B0N 12 VNW pch L=4e-08 W=4e-07 
M30 13 B0N 2 VNW pch L=4e-08 W=4e-07 
M31 VDD B1N 13 VNW pch L=4e-08 W=4e-07 
M32 Y 2 4 VNW pch L=4e-08 W=4e-07 
M33 4 2 Y VNW pch L=4e-08 W=4e-07 
M34 Y 2 4 VNW pch L=4e-08 W=4e-07 
M35 4 2 Y VNW pch L=4e-08 W=4e-07 
M36 Y 2 4 VNW pch L=4e-08 W=4e-07 
M37 4 2 Y VNW pch L=4e-08 W=4e-07 
M38 Y 2 4 VNW pch L=4e-08 W=4e-07 
M39 4 2 Y VNW pch L=4e-08 W=4e-07 
M40 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M41 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M42 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M43 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M44 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M45 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M46 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M47 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M48 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M49 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M50 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M51 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M52 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M53 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M54 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M55 4 A0 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 9 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A0 9 VPW nch L=4e-08 W=1.2e-07 
M2 10 B0 Y VPW nch L=4e-08 W=1.2e-07 
M3 VSS B1 10 VPW nch L=4e-08 W=1.2e-07 
M4 VDD A1 2 VNW pch L=4e-08 W=2.1e-07 
M5 2 A0 VDD VNW pch L=4e-08 W=2.1e-07 
M6 Y B0 2 VNW pch L=4e-08 W=2.1e-07 
M7 2 B1 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT AOI22_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 9 A1 VSS VPW nch L=4e-08 W=1.7e-07 
M1 Y A0 9 VPW nch L=4e-08 W=1.7e-07 
M2 10 B0 Y VPW nch L=4e-08 W=1.7e-07 
M3 VSS B1 10 VPW nch L=4e-08 W=1.7e-07 
M4 VDD A1 2 VNW pch L=4e-08 W=2.85e-07 
M5 2 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M6 Y B0 2 VNW pch L=4e-08 W=2.85e-07 
M7 2 B1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI22_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 9 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M1 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M2 10 B0 Y VPW nch L=4e-08 W=2.4e-07 
M3 VSS B1 10 VPW nch L=4e-08 W=2.4e-07 
M4 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M5 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M6 Y B0 2 VNW pch L=4e-08 W=4e-07 
M7 2 B1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 10 A1 VSS VPW nch L=4e-08 W=3.4e-07 
M1 Y A0 10 VPW nch L=4e-08 W=3.4e-07 
M2 11 B0 Y VPW nch L=4e-08 W=3.4e-07 
M3 VSS B1 11 VPW nch L=4e-08 W=3.4e-07 
M4 VDD A0 1 VNW pch L=4e-08 W=2.85e-07 
M5 1 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M6 VDD A1 1 VNW pch L=4e-08 W=2.85e-07 
M7 1 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M8 Y B0 1 VNW pch L=4e-08 W=2.85e-07 
M9 1 B1 Y VNW pch L=4e-08 W=2.85e-07 
M10 Y B1 1 VNW pch L=4e-08 W=2.85e-07 
M11 1 B0 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI22_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 9 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M1 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M2 10 A0 Y VPW nch L=4e-08 W=2.4e-07 
M3 VSS A1 10 VPW nch L=4e-08 W=2.4e-07 
M4 11 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M5 Y B0 11 VPW nch L=4e-08 W=2.4e-07 
M6 12 B0 Y VPW nch L=4e-08 W=2.4e-07 
M7 VSS B1 12 VPW nch L=4e-08 W=2.4e-07 
M8 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M9 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M11 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M12 Y B1 2 VNW pch L=4e-08 W=4e-07 
M13 2 B0 Y VNW pch L=4e-08 W=4e-07 
M14 Y B0 2 VNW pch L=4e-08 W=4e-07 
M15 2 B1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 9 A0 Y VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1 9 VPW nch L=4e-08 W=2.4e-07 
M2 10 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y A0 10 VPW nch L=4e-08 W=2.4e-07 
M4 11 A0 Y VPW nch L=4e-08 W=2.4e-07 
M5 VSS A1 11 VPW nch L=4e-08 W=2.4e-07 
M6 12 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M7 Y B0 12 VPW nch L=4e-08 W=2.4e-07 
M8 13 B0 Y VPW nch L=4e-08 W=2.4e-07 
M9 VSS B1 13 VPW nch L=4e-08 W=2.4e-07 
M10 14 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M11 Y B0 14 VPW nch L=4e-08 W=2.4e-07 
M12 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M13 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M15 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M17 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M18 Y B1 2 VNW pch L=4e-08 W=4e-07 
M19 2 B0 Y VNW pch L=4e-08 W=4e-07 
M20 Y B0 2 VNW pch L=4e-08 W=4e-07 
M21 2 B1 Y VNW pch L=4e-08 W=4e-07 
M22 Y B1 2 VNW pch L=4e-08 W=4e-07 
M23 2 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 9 A0 Y VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1 9 VPW nch L=4e-08 W=2.4e-07 
M2 10 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y A0 10 VPW nch L=4e-08 W=2.4e-07 
M4 11 A0 Y VPW nch L=4e-08 W=2.4e-07 
M5 VSS A1 11 VPW nch L=4e-08 W=2.4e-07 
M6 12 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M7 Y A0 12 VPW nch L=4e-08 W=2.4e-07 
M8 13 B0 Y VPW nch L=4e-08 W=2.4e-07 
M9 VSS B1 13 VPW nch L=4e-08 W=2.4e-07 
M10 14 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M11 Y B0 14 VPW nch L=4e-08 W=2.4e-07 
M12 15 B0 Y VPW nch L=4e-08 W=2.4e-07 
M13 VSS B1 15 VPW nch L=4e-08 W=2.4e-07 
M14 16 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M15 Y B0 16 VPW nch L=4e-08 W=2.4e-07 
M16 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M17 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M19 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M21 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M23 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M24 Y B0 2 VNW pch L=4e-08 W=4e-07 
M25 2 B1 Y VNW pch L=4e-08 W=4e-07 
M26 Y B1 2 VNW pch L=4e-08 W=4e-07 
M27 2 B0 Y VNW pch L=4e-08 W=4e-07 
M28 Y B0 2 VNW pch L=4e-08 W=4e-07 
M29 2 B1 Y VNW pch L=4e-08 W=4e-07 
M30 Y B1 2 VNW pch L=4e-08 W=4e-07 
M31 2 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 9 A0 Y VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1 9 VPW nch L=4e-08 W=2.4e-07 
M2 10 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y A0 10 VPW nch L=4e-08 W=2.4e-07 
M4 11 A0 Y VPW nch L=4e-08 W=2.4e-07 
M5 VSS A1 11 VPW nch L=4e-08 W=2.4e-07 
M6 12 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M7 Y A0 12 VPW nch L=4e-08 W=2.4e-07 
M8 13 A0 Y VPW nch L=4e-08 W=2.4e-07 
M9 VSS A1 13 VPW nch L=4e-08 W=2.4e-07 
M10 14 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M11 Y A0 14 VPW nch L=4e-08 W=2.4e-07 
M12 15 B0 Y VPW nch L=4e-08 W=2.4e-07 
M13 VSS B1 15 VPW nch L=4e-08 W=2.4e-07 
M14 16 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M15 Y B0 16 VPW nch L=4e-08 W=2.4e-07 
M16 17 B0 Y VPW nch L=4e-08 W=2.4e-07 
M17 VSS B1 17 VPW nch L=4e-08 W=2.4e-07 
M18 18 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M19 Y B0 18 VPW nch L=4e-08 W=2.4e-07 
M20 19 B0 Y VPW nch L=4e-08 W=2.4e-07 
M21 VSS B1 19 VPW nch L=4e-08 W=2.4e-07 
M22 20 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M23 Y B0 20 VPW nch L=4e-08 W=2.4e-07 
M24 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M25 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M27 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M29 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M31 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M33 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M35 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M36 Y B0 2 VNW pch L=4e-08 W=4e-07 
M37 2 B1 Y VNW pch L=4e-08 W=4e-07 
M38 Y B1 2 VNW pch L=4e-08 W=4e-07 
M39 2 B0 Y VNW pch L=4e-08 W=4e-07 
M40 Y B0 2 VNW pch L=4e-08 W=4e-07 
M41 2 B1 Y VNW pch L=4e-08 W=4e-07 
M42 Y B1 2 VNW pch L=4e-08 W=4e-07 
M43 2 B0 Y VNW pch L=4e-08 W=4e-07 
M44 Y B0 2 VNW pch L=4e-08 W=4e-07 
M45 2 B1 Y VNW pch L=4e-08 W=4e-07 
M46 Y B1 2 VNW pch L=4e-08 W=4e-07 
M47 2 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI22_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 9 A0 Y VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1 9 VPW nch L=4e-08 W=2.4e-07 
M2 10 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y A0 10 VPW nch L=4e-08 W=2.4e-07 
M4 11 A0 Y VPW nch L=4e-08 W=2.4e-07 
M5 VSS A1 11 VPW nch L=4e-08 W=2.4e-07 
M6 12 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M7 Y A0 12 VPW nch L=4e-08 W=2.4e-07 
M8 13 A0 Y VPW nch L=4e-08 W=2.4e-07 
M9 VSS A1 13 VPW nch L=4e-08 W=2.4e-07 
M10 14 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M11 Y A0 14 VPW nch L=4e-08 W=2.4e-07 
M12 15 A0 Y VPW nch L=4e-08 W=2.4e-07 
M13 VSS A1 15 VPW nch L=4e-08 W=2.4e-07 
M14 16 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M15 Y A0 16 VPW nch L=4e-08 W=2.4e-07 
M16 17 B0 Y VPW nch L=4e-08 W=2.4e-07 
M17 VSS B1 17 VPW nch L=4e-08 W=2.4e-07 
M18 18 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M19 Y B0 18 VPW nch L=4e-08 W=2.4e-07 
M20 19 B0 Y VPW nch L=4e-08 W=2.4e-07 
M21 VSS B1 19 VPW nch L=4e-08 W=2.4e-07 
M22 20 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M23 Y B0 20 VPW nch L=4e-08 W=2.4e-07 
M24 21 B0 Y VPW nch L=4e-08 W=2.4e-07 
M25 VSS B1 21 VPW nch L=4e-08 W=2.4e-07 
M26 22 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M27 Y B0 22 VPW nch L=4e-08 W=2.4e-07 
M28 23 B0 Y VPW nch L=4e-08 W=2.4e-07 
M29 VSS B1 23 VPW nch L=4e-08 W=2.4e-07 
M30 24 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M31 Y B0 24 VPW nch L=4e-08 W=2.4e-07 
M32 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M33 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M35 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M37 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M39 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M41 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M42 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M43 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M44 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M45 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M46 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M47 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M48 Y B0 2 VNW pch L=4e-08 W=4e-07 
M49 2 B1 Y VNW pch L=4e-08 W=4e-07 
M50 Y B1 2 VNW pch L=4e-08 W=4e-07 
M51 2 B0 Y VNW pch L=4e-08 W=4e-07 
M52 Y B0 2 VNW pch L=4e-08 W=4e-07 
M53 2 B1 Y VNW pch L=4e-08 W=4e-07 
M54 Y B1 2 VNW pch L=4e-08 W=4e-07 
M55 2 B0 Y VNW pch L=4e-08 W=4e-07 
M56 Y B0 2 VNW pch L=4e-08 W=4e-07 
M57 2 B1 Y VNW pch L=4e-08 W=4e-07 
M58 Y B1 2 VNW pch L=4e-08 W=4e-07 
M59 2 B0 Y VNW pch L=4e-08 W=4e-07 
M60 Y B0 2 VNW pch L=4e-08 W=4e-07 
M61 2 B1 Y VNW pch L=4e-08 W=4e-07 
M62 Y B1 2 VNW pch L=4e-08 W=4e-07 
M63 2 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI2XB1_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=1.2e-07 
M1 9 3 VSS VPW nch L=4e-08 W=1.2e-07 
M2 Y A0 9 VPW nch L=4e-08 W=1.2e-07 
M3 VSS B0 Y VPW nch L=4e-08 W=1.2e-07 
M4 3 A1N VDD VNW pch L=4e-08 W=1.55e-07 
M5 VDD 3 4 VNW pch L=4e-08 W=2e-07 
M6 4 A0 VDD VNW pch L=4e-08 W=2e-07 
M7 Y B0 4 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AOI2XB1_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=1.2e-07 
M1 9 3 VSS VPW nch L=4e-08 W=1.8e-07 
M2 Y A0 9 VPW nch L=4e-08 W=1.8e-07 
M3 VSS B0 Y VPW nch L=4e-08 W=1.2e-07 
M4 3 A1N VDD VNW pch L=4e-08 W=1.55e-07 
M5 VDD 3 4 VNW pch L=4e-08 W=3e-07 
M6 4 A0 VDD VNW pch L=4e-08 W=3e-07 
M7 Y B0 4 VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT AOI2XB1_X1M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=1.2e-07 
M1 9 3 VSS VPW nch L=4e-08 W=2.4e-07 
M2 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M3 VSS B0 Y VPW nch L=4e-08 W=1.6e-07 
M4 3 A1N VDD VNW pch L=4e-08 W=1.55e-07 
M5 VDD 3 4 VNW pch L=4e-08 W=4e-07 
M6 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M7 Y B0 4 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI2XB1_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=1.25e-07 
M1 10 3 VSS VPW nch L=4e-08 W=3.4e-07 
M2 Y A0 10 VPW nch L=4e-08 W=3.4e-07 
M3 VSS B0 Y VPW nch L=4e-08 W=2.3e-07 
M4 3 A1N VDD VNW pch L=4e-08 W=1.6e-07 
M5 VDD A0 4 VNW pch L=4e-08 W=2.85e-07 
M6 4 3 VDD VNW pch L=4e-08 W=2.85e-07 
M7 VDD 3 4 VNW pch L=4e-08 W=2.85e-07 
M8 4 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M9 Y B0 4 VNW pch L=4e-08 W=2.85e-07 
M10 4 B0 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI2XB1_X2M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=1.65e-07 
M1 9 3 VSS VPW nch L=4e-08 W=2.4e-07 
M2 Y A0 9 VPW nch L=4e-08 W=2.4e-07 
M3 10 A0 Y VPW nch L=4e-08 W=2.4e-07 
M4 VSS 3 10 VPW nch L=4e-08 W=2.4e-07 
M5 Y B0 VSS VPW nch L=4e-08 W=1.6e-07 
M6 VSS B0 Y VPW nch L=4e-08 W=1.6e-07 
M7 3 A1N VDD VNW pch L=4e-08 W=2.1e-07 
M8 VDD 3 4 VNW pch L=4e-08 W=4e-07 
M9 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M11 4 3 VDD VNW pch L=4e-08 W=4e-07 
M12 Y B0 4 VNW pch L=4e-08 W=4e-07 
M13 4 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI2XB1_X3M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=2.4e-07 
M1 9 A0 Y VPW nch L=4e-08 W=2.4e-07 
M2 VSS 3 9 VPW nch L=4e-08 W=2.4e-07 
M3 10 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 Y A0 10 VPW nch L=4e-08 W=2.4e-07 
M5 11 A0 Y VPW nch L=4e-08 W=2.4e-07 
M6 VSS 3 11 VPW nch L=4e-08 W=2.4e-07 
M7 Y B0 VSS VPW nch L=4e-08 W=2.4e-07 
M8 VSS B0 Y VPW nch L=4e-08 W=2.4e-07 
M9 3 A1N VDD VNW pch L=4e-08 W=3.1e-07 
M10 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M11 5 3 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M13 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M15 5 3 VDD VNW pch L=4e-08 W=4e-07 
M16 Y B0 5 VNW pch L=4e-08 W=4e-07 
M17 5 B0 Y VNW pch L=4e-08 W=4e-07 
M18 Y B0 5 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI2XB1_X4M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=3.1e-07 
M1 9 A0 Y VPW nch L=4e-08 W=2.4e-07 
M2 VSS 3 9 VPW nch L=4e-08 W=2.4e-07 
M3 10 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 Y A0 10 VPW nch L=4e-08 W=2.4e-07 
M5 11 A0 Y VPW nch L=4e-08 W=2.4e-07 
M6 VSS 3 11 VPW nch L=4e-08 W=2.4e-07 
M7 12 3 VSS VPW nch L=4e-08 W=2.4e-07 
M8 Y A0 12 VPW nch L=4e-08 W=2.4e-07 
M9 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M10 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M11 3 A1N VDD VNW pch L=4e-08 W=4e-07 
M12 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M13 5 3 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M15 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M17 5 3 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M19 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M20 Y B0 5 VNW pch L=4e-08 W=4e-07 
M21 5 B0 Y VNW pch L=4e-08 W=4e-07 
M22 Y B0 5 VNW pch L=4e-08 W=4e-07 
M23 5 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI2XB1_X6M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1N 3 VPW nch L=4e-08 W=2.4e-07 
M2 9 A0 Y VPW nch L=4e-08 W=2.4e-07 
M3 VSS 3 9 VPW nch L=4e-08 W=2.4e-07 
M4 10 3 VSS VPW nch L=4e-08 W=2.4e-07 
M5 Y A0 10 VPW nch L=4e-08 W=2.4e-07 
M6 11 A0 Y VPW nch L=4e-08 W=2.4e-07 
M7 VSS 3 11 VPW nch L=4e-08 W=2.4e-07 
M8 12 3 VSS VPW nch L=4e-08 W=2.4e-07 
M9 Y A0 12 VPW nch L=4e-08 W=2.4e-07 
M10 13 A0 Y VPW nch L=4e-08 W=2.4e-07 
M11 VSS 3 13 VPW nch L=4e-08 W=2.4e-07 
M12 14 3 VSS VPW nch L=4e-08 W=2.4e-07 
M13 Y A0 14 VPW nch L=4e-08 W=2.4e-07 
M14 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M15 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M16 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M17 3 A1N VDD VNW pch L=4e-08 W=3.05e-07 
M18 VDD A1N 3 VNW pch L=4e-08 W=3.05e-07 
M19 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M20 5 3 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M22 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M24 5 3 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M26 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M28 5 3 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M30 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M31 Y B0 5 VNW pch L=4e-08 W=4e-07 
M32 5 B0 Y VNW pch L=4e-08 W=4e-07 
M33 Y B0 5 VNW pch L=4e-08 W=4e-07 
M34 5 B0 Y VNW pch L=4e-08 W=4e-07 
M35 Y B0 5 VNW pch L=4e-08 W=4e-07 
M36 5 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI2XB1_X8M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A1N 3 VPW nch L=4e-08 W=3.1e-07 
M2 9 A0 Y VPW nch L=4e-08 W=2.4e-07 
M3 VSS 3 9 VPW nch L=4e-08 W=2.4e-07 
M4 10 3 VSS VPW nch L=4e-08 W=2.4e-07 
M5 Y A0 10 VPW nch L=4e-08 W=2.4e-07 
M6 11 A0 Y VPW nch L=4e-08 W=2.4e-07 
M7 VSS 3 11 VPW nch L=4e-08 W=2.4e-07 
M8 12 3 VSS VPW nch L=4e-08 W=2.4e-07 
M9 Y A0 12 VPW nch L=4e-08 W=2.4e-07 
M10 13 A0 Y VPW nch L=4e-08 W=2.4e-07 
M11 VSS 3 13 VPW nch L=4e-08 W=2.4e-07 
M12 14 3 VSS VPW nch L=4e-08 W=2.4e-07 
M13 Y A0 14 VPW nch L=4e-08 W=2.4e-07 
M14 15 A0 Y VPW nch L=4e-08 W=2.4e-07 
M15 VSS 3 15 VPW nch L=4e-08 W=2.4e-07 
M16 16 3 VSS VPW nch L=4e-08 W=2.4e-07 
M17 Y A0 16 VPW nch L=4e-08 W=2.4e-07 
M18 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M19 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M20 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M21 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M22 3 A1N VDD VNW pch L=4e-08 W=4e-07 
M23 VDD A1N 3 VNW pch L=4e-08 W=4e-07 
M24 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M25 5 3 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M27 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M29 5 3 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M31 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M33 5 3 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M35 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD A0 5 VNW pch L=4e-08 W=4e-07 
M37 5 3 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 3 5 VNW pch L=4e-08 W=4e-07 
M39 5 A0 VDD VNW pch L=4e-08 W=4e-07 
M40 Y B0 5 VNW pch L=4e-08 W=4e-07 
M41 5 B0 Y VNW pch L=4e-08 W=4e-07 
M42 Y B0 5 VNW pch L=4e-08 W=4e-07 
M43 5 B0 Y VNW pch L=4e-08 W=4e-07 
M44 Y B0 5 VNW pch L=4e-08 W=4e-07 
M45 5 B0 Y VNW pch L=4e-08 W=4e-07 
M46 Y B0 5 VNW pch L=4e-08 W=4e-07 
M47 5 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI31_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 9 A2 VSS VPW nch L=4e-08 W=1.55e-07 
M1 10 A1 9 VPW nch L=4e-08 W=1.55e-07 
M2 Y A0 10 VPW nch L=4e-08 W=1.55e-07 
M3 VSS B0 Y VPW nch L=4e-08 W=1.2e-07 
M4 3 A2 VDD VNW pch L=4e-08 W=2e-07 
M5 VDD A1 3 VNW pch L=4e-08 W=2e-07 
M6 3 A0 VDD VNW pch L=4e-08 W=2e-07 
M7 Y B0 3 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT AOI31_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 9 A2 VSS VPW nch L=4e-08 W=2.3e-07 
M1 10 A1 9 VPW nch L=4e-08 W=2.3e-07 
M2 Y A0 10 VPW nch L=4e-08 W=2.3e-07 
M3 VSS B0 Y VPW nch L=4e-08 W=1.2e-07 
M4 3 A2 VDD VNW pch L=4e-08 W=2.95e-07 
M5 VDD A1 3 VNW pch L=4e-08 W=2.95e-07 
M6 3 A0 VDD VNW pch L=4e-08 W=2.95e-07 
M7 Y B0 3 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT AOI31_X1M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 9 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M1 10 A1 9 VPW nch L=4e-08 W=3.1e-07 
M2 Y A0 10 VPW nch L=4e-08 W=3.1e-07 
M3 VSS B0 Y VPW nch L=4e-08 W=1.6e-07 
M4 3 A2 VDD VNW pch L=4e-08 W=4e-07 
M5 VDD A1 3 VNW pch L=4e-08 W=4e-07 
M6 3 A0 VDD VNW pch L=4e-08 W=4e-07 
M7 Y B0 3 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI31_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 VSS A2 1 VPW nch L=4e-08 W=2.2e-07 
M1 1 A2 VSS VPW nch L=4e-08 W=2.2e-07 
M2 10 A1 1 VPW nch L=4e-08 W=2.2e-07 
M3 Y A0 10 VPW nch L=4e-08 W=2.2e-07 
M4 11 A0 Y VPW nch L=4e-08 W=2.2e-07 
M5 1 A1 11 VPW nch L=4e-08 W=2.2e-07 
M6 Y B0 VSS VPW nch L=4e-08 W=2.3e-07 
M7 VDD A2 2 VNW pch L=4e-08 W=2.85e-07 
M8 2 A2 VDD VNW pch L=4e-08 W=2.85e-07 
M9 VDD A1 2 VNW pch L=4e-08 W=2.85e-07 
M10 2 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M11 VDD A0 2 VNW pch L=4e-08 W=2.85e-07 
M12 2 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M13 Y B0 2 VNW pch L=4e-08 W=2.85e-07 
M14 2 B0 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI31_X2M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M2 10 A1 1 VPW nch L=4e-08 W=3.1e-07 
M3 Y A0 10 VPW nch L=4e-08 W=3.1e-07 
M4 11 A0 Y VPW nch L=4e-08 W=3.1e-07 
M5 1 A1 11 VPW nch L=4e-08 W=3.1e-07 
M6 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M7 VDD A2 2 VNW pch L=4e-08 W=4e-07 
M8 2 A2 VDD VNW pch L=4e-08 W=4e-07 
M9 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M10 2 A0 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD A0 2 VNW pch L=4e-08 W=4e-07 
M12 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y B0 2 VNW pch L=4e-08 W=4e-07 
M14 2 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI31_X3M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 3 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A2 3 VPW nch L=4e-08 W=3.1e-07 
M2 3 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M3 10 A1 3 VPW nch L=4e-08 W=3.1e-07 
M4 Y A0 10 VPW nch L=4e-08 W=3.1e-07 
M5 11 A0 Y VPW nch L=4e-08 W=3.1e-07 
M6 3 A1 11 VPW nch L=4e-08 W=3.1e-07 
M7 12 A1 3 VPW nch L=4e-08 W=3.1e-07 
M8 Y A0 12 VPW nch L=4e-08 W=3.1e-07 
M9 VSS B0 Y VPW nch L=4e-08 W=2.4e-07 
M10 Y B0 VSS VPW nch L=4e-08 W=2.4e-07 
M11 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M13 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M15 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M17 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M19 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M20 Y B0 4 VNW pch L=4e-08 W=4e-07 
M21 4 B0 Y VNW pch L=4e-08 W=4e-07 
M22 Y B0 4 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI31_X4M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M4 10 A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 Y A0 10 VPW nch L=4e-08 W=3.1e-07 
M6 11 A0 Y VPW nch L=4e-08 W=3.1e-07 
M7 1 A1 11 VPW nch L=4e-08 W=3.1e-07 
M8 12 A1 1 VPW nch L=4e-08 W=3.1e-07 
M9 Y A0 12 VPW nch L=4e-08 W=3.1e-07 
M10 13 A0 Y VPW nch L=4e-08 W=3.1e-07 
M11 1 A1 13 VPW nch L=4e-08 W=3.1e-07 
M12 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M13 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M14 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M16 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M17 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M18 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M20 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M22 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M24 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M26 Y B0 4 VNW pch L=4e-08 W=4e-07 
M27 4 B0 Y VNW pch L=4e-08 W=4e-07 
M28 Y B0 4 VNW pch L=4e-08 W=4e-07 
M29 4 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI31_X6M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M6 10 A1 1 VPW nch L=4e-08 W=3.1e-07 
M7 Y A0 10 VPW nch L=4e-08 W=3.1e-07 
M8 11 A0 Y VPW nch L=4e-08 W=3.1e-07 
M9 1 A1 11 VPW nch L=4e-08 W=3.1e-07 
M10 12 A1 1 VPW nch L=4e-08 W=3.1e-07 
M11 Y A0 12 VPW nch L=4e-08 W=3.1e-07 
M12 13 A0 Y VPW nch L=4e-08 W=3.1e-07 
M13 1 A1 13 VPW nch L=4e-08 W=3.1e-07 
M14 14 A1 1 VPW nch L=4e-08 W=3.1e-07 
M15 Y A0 14 VPW nch L=4e-08 W=3.1e-07 
M16 15 A0 Y VPW nch L=4e-08 W=3.1e-07 
M17 1 A1 15 VPW nch L=4e-08 W=3.1e-07 
M18 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M19 VSS B0 Y VPW nch L=4e-08 W=3.2e-07 
M20 Y B0 VSS VPW nch L=4e-08 W=3.2e-07 
M21 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M23 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M25 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M27 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M29 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M31 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M33 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M35 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M37 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M39 Y B0 4 VNW pch L=4e-08 W=4e-07 
M40 4 B0 Y VNW pch L=4e-08 W=4e-07 
M41 Y B0 4 VNW pch L=4e-08 W=4e-07 
M42 4 B0 Y VNW pch L=4e-08 W=4e-07 
M43 Y B0 4 VNW pch L=4e-08 W=4e-07 
M44 4 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI32_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
M0 10 A2 VSS VPW nch L=4e-08 W=1.55e-07 
M1 11 A1 10 VPW nch L=4e-08 W=1.55e-07 
M2 Y A0 11 VPW nch L=4e-08 W=1.55e-07 
M3 12 B0 Y VPW nch L=4e-08 W=1.2e-07 
M4 VSS B1 12 VPW nch L=4e-08 W=1.2e-07 
M5 3 A2 VDD VNW pch L=4e-08 W=2.1e-07 
M6 VDD A1 3 VNW pch L=4e-08 W=2.1e-07 
M7 3 A0 VDD VNW pch L=4e-08 W=2.1e-07 
M8 Y B0 3 VNW pch L=4e-08 W=2.1e-07 
M9 3 B1 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT AOI32_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
M0 10 A2 VSS VPW nch L=4e-08 W=2.2e-07 
M1 11 A1 10 VPW nch L=4e-08 W=2.2e-07 
M2 Y A0 11 VPW nch L=4e-08 W=2.2e-07 
M3 12 B0 Y VPW nch L=4e-08 W=1.7e-07 
M4 VSS B1 12 VPW nch L=4e-08 W=1.7e-07 
M5 3 A2 VDD VNW pch L=4e-08 W=2.85e-07 
M6 VDD A1 3 VNW pch L=4e-08 W=2.85e-07 
M7 3 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M8 Y B0 3 VNW pch L=4e-08 W=2.85e-07 
M9 3 B1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI32_X1M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
M0 10 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M1 11 A1 10 VPW nch L=4e-08 W=3.1e-07 
M2 Y A0 11 VPW nch L=4e-08 W=3.1e-07 
M3 12 B0 Y VPW nch L=4e-08 W=2.4e-07 
M4 VSS B1 12 VPW nch L=4e-08 W=2.4e-07 
M5 3 A2 VDD VNW pch L=4e-08 W=4e-07 
M6 VDD A1 3 VNW pch L=4e-08 W=4e-07 
M7 3 A0 VDD VNW pch L=4e-08 W=4e-07 
M8 Y B0 3 VNW pch L=4e-08 W=4e-07 
M9 3 B1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI32_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
M0 VSS A2 1 VPW nch L=4e-08 W=2.2e-07 
M1 1 A2 VSS VPW nch L=4e-08 W=2.2e-07 
M2 11 A1 1 VPW nch L=4e-08 W=2.2e-07 
M3 Y A0 11 VPW nch L=4e-08 W=2.2e-07 
M4 12 A0 Y VPW nch L=4e-08 W=2.2e-07 
M5 1 A1 12 VPW nch L=4e-08 W=2.2e-07 
M6 13 B1 VSS VPW nch L=4e-08 W=1.7e-07 
M7 Y B0 13 VPW nch L=4e-08 W=1.7e-07 
M8 14 B0 Y VPW nch L=4e-08 W=1.7e-07 
M9 VSS B1 14 VPW nch L=4e-08 W=1.7e-07 
M10 4 A2 VDD VNW pch L=4e-08 W=2.85e-07 
M11 VDD A2 4 VNW pch L=4e-08 W=2.85e-07 
M12 4 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M13 VDD A0 4 VNW pch L=4e-08 W=2.85e-07 
M14 4 A0 VDD VNW pch L=4e-08 W=2.85e-07 
M15 VDD A1 4 VNW pch L=4e-08 W=2.85e-07 
M16 Y B1 4 VNW pch L=4e-08 W=2.85e-07 
M17 4 B0 Y VNW pch L=4e-08 W=2.85e-07 
M18 Y B0 4 VNW pch L=4e-08 W=2.85e-07 
M19 4 B1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT AOI32_X2M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
M0 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M2 11 A1 1 VPW nch L=4e-08 W=3.1e-07 
M3 Y A0 11 VPW nch L=4e-08 W=3.1e-07 
M4 12 A0 Y VPW nch L=4e-08 W=3.1e-07 
M5 1 A1 12 VPW nch L=4e-08 W=3.1e-07 
M6 13 B1 VSS VPW nch L=4e-08 W=2.4e-07 
M7 Y B0 13 VPW nch L=4e-08 W=2.4e-07 
M8 14 B0 Y VPW nch L=4e-08 W=2.4e-07 
M9 VSS B1 14 VPW nch L=4e-08 W=2.4e-07 
M10 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M12 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M14 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M16 Y B1 4 VNW pch L=4e-08 W=4e-07 
M17 4 B0 Y VNW pch L=4e-08 W=4e-07 
M18 Y B0 4 VNW pch L=4e-08 W=4e-07 
M19 4 B1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI32_X3M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
M0 3 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A2 3 VPW nch L=4e-08 W=3.1e-07 
M2 3 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M3 11 A1 3 VPW nch L=4e-08 W=3.1e-07 
M4 Y A0 11 VPW nch L=4e-08 W=3.1e-07 
M5 12 A0 Y VPW nch L=4e-08 W=3.1e-07 
M6 3 A1 12 VPW nch L=4e-08 W=3.1e-07 
M7 13 A1 3 VPW nch L=4e-08 W=3.1e-07 
M8 Y A0 13 VPW nch L=4e-08 W=3.1e-07 
M9 14 B0 Y VPW nch L=4e-08 W=3.6e-07 
M10 VSS B1 14 VPW nch L=4e-08 W=3.6e-07 
M11 15 B1 VSS VPW nch L=4e-08 W=3.6e-07 
M12 Y B0 15 VPW nch L=4e-08 W=3.6e-07 
M13 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M15 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M17 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M19 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M21 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M22 Y B0 4 VNW pch L=4e-08 W=4e-07 
M23 4 B1 Y VNW pch L=4e-08 W=4e-07 
M24 Y B1 4 VNW pch L=4e-08 W=4e-07 
M25 4 B0 Y VNW pch L=4e-08 W=4e-07 
M26 Y B0 4 VNW pch L=4e-08 W=4e-07 
M27 4 B1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI32_X4M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
M0 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M4 11 A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 Y A0 11 VPW nch L=4e-08 W=3.1e-07 
M6 12 A0 Y VPW nch L=4e-08 W=3.1e-07 
M7 1 A1 12 VPW nch L=4e-08 W=3.1e-07 
M8 13 A1 1 VPW nch L=4e-08 W=3.1e-07 
M9 Y A0 13 VPW nch L=4e-08 W=3.1e-07 
M10 14 A0 Y VPW nch L=4e-08 W=3.1e-07 
M11 1 A1 14 VPW nch L=4e-08 W=3.1e-07 
M12 16 B1 VSS VPW nch L=4e-08 W=3.2e-07 
M13 Y B0 16 VPW nch L=4e-08 W=3.2e-07 
M14 17 B0 Y VPW nch L=4e-08 W=3.2e-07 
M15 VSS B1 17 VPW nch L=4e-08 W=3.2e-07 
M16 18 B1 VSS VPW nch L=4e-08 W=3.2e-07 
M17 Y B0 18 VPW nch L=4e-08 W=3.2e-07 
M18 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M20 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M22 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M24 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M26 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M28 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M30 Y B0 4 VNW pch L=4e-08 W=4e-07 
M31 4 B1 Y VNW pch L=4e-08 W=4e-07 
M32 Y B1 4 VNW pch L=4e-08 W=4e-07 
M33 4 B0 Y VNW pch L=4e-08 W=4e-07 
M34 Y B0 4 VNW pch L=4e-08 W=4e-07 
M35 4 B1 Y VNW pch L=4e-08 W=4e-07 
M36 Y B1 4 VNW pch L=4e-08 W=4e-07 
M37 4 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT AOI32_X6M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
M0 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A2 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A2 VSS VPW nch L=4e-08 W=3.1e-07 
M6 11 A1 1 VPW nch L=4e-08 W=3.1e-07 
M7 Y A0 11 VPW nch L=4e-08 W=3.1e-07 
M8 12 A0 Y VPW nch L=4e-08 W=3.1e-07 
M9 1 A1 12 VPW nch L=4e-08 W=3.1e-07 
M10 13 A1 1 VPW nch L=4e-08 W=3.1e-07 
M11 Y A0 13 VPW nch L=4e-08 W=3.1e-07 
M12 14 A0 Y VPW nch L=4e-08 W=3.1e-07 
M13 1 A1 14 VPW nch L=4e-08 W=3.1e-07 
M14 15 A1 1 VPW nch L=4e-08 W=3.1e-07 
M15 Y A0 15 VPW nch L=4e-08 W=3.1e-07 
M16 16 A0 Y VPW nch L=4e-08 W=3.1e-07 
M17 1 A1 16 VPW nch L=4e-08 W=3.1e-07 
M18 18 B1 VSS VPW nch L=4e-08 W=3.6e-07 
M19 Y B0 18 VPW nch L=4e-08 W=3.6e-07 
M20 19 B0 Y VPW nch L=4e-08 W=3.6e-07 
M21 VSS B1 19 VPW nch L=4e-08 W=3.6e-07 
M22 20 B1 VSS VPW nch L=4e-08 W=3.6e-07 
M23 Y B0 20 VPW nch L=4e-08 W=3.6e-07 
M24 21 B0 Y VPW nch L=4e-08 W=3.6e-07 
M25 VSS B1 21 VPW nch L=4e-08 W=3.6e-07 
M26 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M28 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M30 4 A2 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD A2 4 VNW pch L=4e-08 W=4e-07 
M32 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M33 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M34 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M36 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M38 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M40 4 A1 VDD VNW pch L=4e-08 W=4e-07 
M41 VDD A0 4 VNW pch L=4e-08 W=4e-07 
M42 4 A0 VDD VNW pch L=4e-08 W=4e-07 
M43 VDD A1 4 VNW pch L=4e-08 W=4e-07 
M44 Y B0 4 VNW pch L=4e-08 W=4e-07 
M45 4 B1 Y VNW pch L=4e-08 W=4e-07 
M46 Y B1 4 VNW pch L=4e-08 W=4e-07 
M47 4 B0 Y VNW pch L=4e-08 W=4e-07 
M48 Y B0 4 VNW pch L=4e-08 W=4e-07 
M49 4 B1 Y VNW pch L=4e-08 W=4e-07 
M50 Y B1 4 VNW pch L=4e-08 W=4e-07 
M51 4 B0 Y VNW pch L=4e-08 W=4e-07 
M52 Y B0 4 VNW pch L=4e-08 W=4e-07 
M53 4 B1 Y VNW pch L=4e-08 W=4e-07 
M54 Y B1 4 VNW pch L=4e-08 W=4e-07 
M55 4 B0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BENC_X11M_A9TR AN SN X2 VDD VNW VPW VSS M0 M1 M2
M0 VSS 4 1 VPW nch L=4e-08 W=2.95e-07 
M1 4 M0 VSS VPW nch L=4e-08 W=2.95e-07 
M2 5 6 4 VPW nch L=4e-08 W=2.95e-07 
M3 1 M1 5 VPW nch L=4e-08 W=2.95e-07 
M4 VSS M1 6 VPW nch L=4e-08 W=2.95e-07 
M5 7 5 VSS VPW nch L=4e-08 W=2.95e-07 
M6 VSS 5 7 VPW nch L=4e-08 W=2.95e-07 
M7 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M8 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M9 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M10 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M11 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M12 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M13 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M14 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M15 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M16 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M17 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M18 9 M2 VSS VPW nch L=4e-08 W=1.75e-07 
M19 VSS M1 10 VPW nch L=4e-08 W=2.45e-07 
M20 10 M0 VSS VPW nch L=4e-08 W=2.45e-07 
M21 11 9 10 VPW nch L=4e-08 W=2.45e-07 
M22 12 11 VSS VPW nch L=4e-08 W=2.95e-07 
M23 VSS 11 12 VPW nch L=4e-08 W=2.95e-07 
M24 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M25 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M26 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M27 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M28 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M29 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M30 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M31 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M32 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M33 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M34 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M35 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M36 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M37 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M38 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M39 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M40 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M41 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M42 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M43 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M44 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M45 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M46 15 16 VSS VPW nch L=4e-08 W=2.95e-07 
M47 VSS 16 15 VPW nch L=4e-08 W=2.95e-07 
M48 17 M2 16 VPW nch L=4e-08 W=2.3e-07 
M49 VSS 4 17 VPW nch L=4e-08 W=2.3e-07 
M50 17 6 VSS VPW nch L=4e-08 W=2.3e-07 
M51 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M52 4 M0 VDD VNW pch L=4e-08 W=3.8e-07 
M53 5 6 1 VNW pch L=4e-08 W=3.8e-07 
M54 4 M1 5 VNW pch L=4e-08 W=3.8e-07 
M55 VDD M1 6 VNW pch L=4e-08 W=3.8e-07 
M56 7 5 VDD VNW pch L=4e-08 W=3.8e-07 
M57 VDD 5 7 VNW pch L=4e-08 W=3.8e-07 
M58 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M59 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M60 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M61 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M62 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M63 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M64 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M65 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M66 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M67 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M68 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M69 9 M2 VDD VNW pch L=4e-08 W=2.25e-07 
M70 21 M1 VDD VNW pch L=4e-08 W=3.8e-07 
M71 11 M0 21 VNW pch L=4e-08 W=3.8e-07 
M72 VDD 9 11 VNW pch L=4e-08 W=2e-07 
M73 12 11 VDD VNW pch L=4e-08 W=3.8e-07 
M74 VDD 11 12 VNW pch L=4e-08 W=3.8e-07 
M75 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M76 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M77 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M78 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M79 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M80 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M81 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M82 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M83 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M84 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M85 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M86 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M87 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M88 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M89 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M90 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M91 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M92 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M93 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M94 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M95 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M96 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M97 15 16 VDD VNW pch L=4e-08 W=3.8e-07 
M98 VDD 16 15 VNW pch L=4e-08 W=3.8e-07 
M99 16 M2 VDD VNW pch L=4e-08 W=2e-07 
M100 22 4 16 VNW pch L=4e-08 W=3.5e-07 
M101 VDD 6 22 VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT BENC_X16M_A9TR AN SN X2 VDD VNW VPW VSS M0 M1 M2
M0 VSS 4 1 VPW nch L=4e-08 W=2.95e-07 
M1 4 M0 VSS VPW nch L=4e-08 W=2.95e-07 
M2 5 6 4 VPW nch L=4e-08 W=2.95e-07 
M3 1 M1 5 VPW nch L=4e-08 W=2.95e-07 
M4 VSS M1 6 VPW nch L=4e-08 W=2.95e-07 
M5 7 5 VSS VPW nch L=4e-08 W=2.95e-07 
M6 VSS 5 7 VPW nch L=4e-08 W=2.95e-07 
M7 7 5 VSS VPW nch L=4e-08 W=2.95e-07 
M8 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M9 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M10 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M11 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M12 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M13 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M14 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M15 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M16 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M17 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M18 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M19 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M20 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M21 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M22 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M23 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M24 9 M2 VSS VPW nch L=4e-08 W=2.95e-07 
M25 VSS M1 10 VPW nch L=4e-08 W=2.35e-07 
M26 10 M0 VSS VPW nch L=4e-08 W=2.35e-07 
M27 VSS M0 10 VPW nch L=4e-08 W=2.35e-07 
M28 10 M1 VSS VPW nch L=4e-08 W=2.35e-07 
M29 11 9 10 VPW nch L=4e-08 W=2.35e-07 
M30 10 9 11 VPW nch L=4e-08 W=2.35e-07 
M31 VSS 11 12 VPW nch L=4e-08 W=2.95e-07 
M32 12 11 VSS VPW nch L=4e-08 W=2.95e-07 
M33 VSS 11 12 VPW nch L=4e-08 W=2.95e-07 
M34 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M35 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M36 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M37 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M38 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M39 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M40 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M41 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M42 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M43 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M44 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M45 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M46 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M47 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M48 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M49 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M50 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M51 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M52 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M53 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M54 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M55 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M56 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M57 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M58 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M59 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M60 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M61 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M62 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M63 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M64 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M65 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M66 15 17 VSS VPW nch L=4e-08 W=2.95e-07 
M67 VSS 17 15 VPW nch L=4e-08 W=2.95e-07 
M68 15 17 VSS VPW nch L=4e-08 W=2.95e-07 
M69 17 M2 16 VPW nch L=4e-08 W=2.2e-07 
M70 16 M2 17 VPW nch L=4e-08 W=2.2e-07 
M71 VSS 6 16 VPW nch L=4e-08 W=2.2e-07 
M72 16 4 VSS VPW nch L=4e-08 W=2.2e-07 
M73 VSS 4 16 VPW nch L=4e-08 W=2.2e-07 
M74 16 6 VSS VPW nch L=4e-08 W=2.2e-07 
M75 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M76 4 M0 VDD VNW pch L=4e-08 W=3.8e-07 
M77 5 6 1 VNW pch L=4e-08 W=3.8e-07 
M78 4 M1 5 VNW pch L=4e-08 W=3.8e-07 
M79 VDD M1 6 VNW pch L=4e-08 W=3.8e-07 
M80 7 5 VDD VNW pch L=4e-08 W=3.8e-07 
M81 VDD 5 7 VNW pch L=4e-08 W=3.8e-07 
M82 7 5 VDD VNW pch L=4e-08 W=3.8e-07 
M83 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M84 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M85 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M86 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M87 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M88 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M89 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M90 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M91 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M92 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M93 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M94 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M95 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M96 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M97 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M98 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M99 9 M2 VDD VNW pch L=4e-08 W=3.8e-07 
M100 21 M1 VDD VNW pch L=4e-08 W=3.8e-07 
M101 11 M0 21 VNW pch L=4e-08 W=3.8e-07 
M102 22 M0 11 VNW pch L=4e-08 W=3.8e-07 
M103 VDD M1 22 VNW pch L=4e-08 W=3.8e-07 
M104 11 9 VDD VNW pch L=4e-08 W=3.8e-07 
M105 VDD 11 12 VNW pch L=4e-08 W=3.8e-07 
M106 12 11 VDD VNW pch L=4e-08 W=3.8e-07 
M107 VDD 11 12 VNW pch L=4e-08 W=3.8e-07 
M108 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M109 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M110 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M111 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M112 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M113 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M114 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M115 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M116 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M117 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M118 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M119 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M120 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M121 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M122 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M123 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M124 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M125 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M126 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M127 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M128 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M129 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M130 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M131 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M132 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M133 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M134 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M135 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M136 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M137 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M138 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M139 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M140 15 17 VDD VNW pch L=4e-08 W=3.8e-07 
M141 VDD 17 15 VNW pch L=4e-08 W=3.8e-07 
M142 15 17 VDD VNW pch L=4e-08 W=3.8e-07 
M143 17 M2 VDD VNW pch L=4e-08 W=1.9e-07 
M144 VDD M2 17 VNW pch L=4e-08 W=1.9e-07 
M145 23 6 VDD VNW pch L=4e-08 W=3.35e-07 
M146 17 4 23 VNW pch L=4e-08 W=3.35e-07 
M147 24 4 17 VNW pch L=4e-08 W=3.35e-07 
M148 VDD 6 24 VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BENC_X2M_A9TR AN SN X2 VDD VNW VPW VSS M0 M1 M2
M0 VSS 4 1 VPW nch L=4e-08 W=2.95e-07 
M1 4 M0 VSS VPW nch L=4e-08 W=2.95e-07 
M2 5 M1 4 VPW nch L=4e-08 W=2.95e-07 
M3 1 6 5 VPW nch L=4e-08 W=2.95e-07 
M4 VSS M1 6 VPW nch L=4e-08 W=2.95e-07 
M5 X2 5 VSS VPW nch L=4e-08 W=2.95e-07 
M6 VSS 5 X2 VPW nch L=4e-08 W=2.95e-07 
M7 8 M2 VSS VPW nch L=4e-08 W=2.05e-07 
M8 18 M1 VSS VPW nch L=4e-08 W=2e-07 
M9 10 M0 18 VPW nch L=4e-08 W=2e-07 
M10 VSS 8 10 VPW nch L=4e-08 W=1.5e-07 
M11 SN 10 VSS VPW nch L=4e-08 W=2.95e-07 
M12 VSS 10 SN VPW nch L=4e-08 W=2.95e-07 
M13 AN 13 VSS VPW nch L=4e-08 W=2.95e-07 
M14 VSS 13 AN VPW nch L=4e-08 W=2.95e-07 
M15 13 M2 VSS VPW nch L=4e-08 W=1.5e-07 
M16 19 4 13 VPW nch L=4e-08 W=2.55e-07 
M17 VSS 6 19 VPW nch L=4e-08 W=2.55e-07 
M18 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M19 4 M0 VDD VNW pch L=4e-08 W=3.8e-07 
M20 5 M1 1 VNW pch L=4e-08 W=3.8e-07 
M21 4 6 5 VNW pch L=4e-08 W=3.8e-07 
M22 VDD M1 6 VNW pch L=4e-08 W=3.8e-07 
M23 X2 5 VDD VNW pch L=4e-08 W=3.8e-07 
M24 VDD 5 X2 VNW pch L=4e-08 W=3.8e-07 
M25 8 M2 VDD VNW pch L=4e-08 W=2.6e-07 
M26 VDD M1 9 VNW pch L=4e-08 W=3.8e-07 
M27 9 M0 VDD VNW pch L=4e-08 W=3.8e-07 
M28 10 8 9 VNW pch L=4e-08 W=3.8e-07 
M29 SN 10 VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD 10 SN VNW pch L=4e-08 W=3.8e-07 
M31 AN 13 VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD 13 AN VNW pch L=4e-08 W=3.8e-07 
M33 14 M2 13 VNW pch L=4e-08 W=3.8e-07 
M34 VDD 4 14 VNW pch L=4e-08 W=3.8e-07 
M35 14 6 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT BENC_X3M_A9TR AN SN X2 VDD VNW VPW VSS M0 M1 M2
M0 VSS 4 1 VPW nch L=4e-08 W=1.55e-07 
M1 4 M0 VSS VPW nch L=4e-08 W=1.55e-07 
M2 5 6 4 VPW nch L=4e-08 W=1.55e-07 
M3 1 M1 5 VPW nch L=4e-08 W=1.55e-07 
M4 VSS M1 6 VPW nch L=4e-08 W=2.8e-07 
M5 VSS 5 7 VPW nch L=4e-08 W=2.4e-07 
M6 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M7 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M8 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M9 9 M2 VSS VPW nch L=4e-08 W=1.5e-07 
M10 VSS M1 10 VPW nch L=4e-08 W=1.8e-07 
M11 10 M0 VSS VPW nch L=4e-08 W=1.8e-07 
M12 11 9 10 VPW nch L=4e-08 W=1.8e-07 
M13 VSS 11 12 VPW nch L=4e-08 W=2.4e-07 
M14 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M15 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M16 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M17 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M18 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M19 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M20 15 16 VSS VPW nch L=4e-08 W=2.4e-07 
M21 17 M2 16 VPW nch L=4e-08 W=1.7e-07 
M22 VSS 4 17 VPW nch L=4e-08 W=1.7e-07 
M23 17 6 VSS VPW nch L=4e-08 W=1.7e-07 
M24 VDD 4 1 VNW pch L=4e-08 W=2e-07 
M25 4 M0 VDD VNW pch L=4e-08 W=2e-07 
M26 5 6 1 VNW pch L=4e-08 W=2e-07 
M27 4 M1 5 VNW pch L=4e-08 W=2e-07 
M28 VDD M1 6 VNW pch L=4e-08 W=3.7e-07 
M29 VDD 5 7 VNW pch L=4e-08 W=3.15e-07 
M30 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M32 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M33 9 M2 VDD VNW pch L=4e-08 W=1.95e-07 
M34 21 M1 VDD VNW pch L=4e-08 W=3e-07 
M35 11 M0 21 VNW pch L=4e-08 W=3e-07 
M36 VDD 9 11 VNW pch L=4e-08 W=1.5e-07 
M37 VDD 11 12 VNW pch L=4e-08 W=3.15e-07 
M38 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M39 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M40 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M41 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M42 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M43 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M44 15 16 VDD VNW pch L=4e-08 W=3.15e-07 
M45 16 M2 VDD VNW pch L=4e-08 W=1.5e-07 
M46 22 4 16 VNW pch L=4e-08 W=2.6e-07 
M47 VDD 6 22 VNW pch L=4e-08 W=2.6e-07 
.ENDS


.SUBCKT BENC_X4M_A9TR AN SN X2 VDD VNW VPW VSS M0 M1 M2
M0 VSS 4 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 M0 VSS VPW nch L=4e-08 W=1.8e-07 
M2 5 6 4 VPW nch L=4e-08 W=1.8e-07 
M3 1 M1 5 VPW nch L=4e-08 W=1.8e-07 
M4 VSS M1 6 VPW nch L=4e-08 W=2.95e-07 
M5 VSS 5 7 VPW nch L=4e-08 W=2.95e-07 
M6 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M7 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M8 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M9 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M10 9 M2 VSS VPW nch L=4e-08 W=1.65e-07 
M11 VSS M1 10 VPW nch L=4e-08 W=2.1e-07 
M12 10 M0 VSS VPW nch L=4e-08 W=2.1e-07 
M13 11 9 10 VPW nch L=4e-08 W=2.1e-07 
M14 VSS 11 12 VPW nch L=4e-08 W=2.95e-07 
M15 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M16 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M17 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M18 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M19 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M20 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M21 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M22 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M23 15 16 VSS VPW nch L=4e-08 W=2.95e-07 
M24 17 M2 16 VPW nch L=4e-08 W=1.95e-07 
M25 VSS 4 17 VPW nch L=4e-08 W=1.95e-07 
M26 17 6 VSS VPW nch L=4e-08 W=1.95e-07 
M27 VDD 4 1 VNW pch L=4e-08 W=2.3e-07 
M28 4 M0 VDD VNW pch L=4e-08 W=2.3e-07 
M29 5 6 1 VNW pch L=4e-08 W=2.3e-07 
M30 4 M1 5 VNW pch L=4e-08 W=2.3e-07 
M31 VDD M1 6 VNW pch L=4e-08 W=3.8e-07 
M32 VDD 5 7 VNW pch L=4e-08 W=3.8e-07 
M33 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M35 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M37 9 M2 VDD VNW pch L=4e-08 W=2.1e-07 
M38 21 M1 VDD VNW pch L=4e-08 W=3.4e-07 
M39 11 M0 21 VNW pch L=4e-08 W=3.4e-07 
M40 VDD 9 11 VNW pch L=4e-08 W=1.7e-07 
M41 VDD 11 12 VNW pch L=4e-08 W=3.8e-07 
M42 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M43 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M44 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M45 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M46 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M47 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M48 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M49 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M50 15 16 VDD VNW pch L=4e-08 W=3.8e-07 
M51 16 M2 VDD VNW pch L=4e-08 W=1.7e-07 
M52 22 4 16 VNW pch L=4e-08 W=2.95e-07 
M53 VDD 6 22 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT BENC_X6M_A9TR AN SN X2 VDD VNW VPW VSS M0 M1 M2
M0 VSS 4 1 VPW nch L=4e-08 W=2.5e-07 
M1 4 M0 VSS VPW nch L=4e-08 W=2.5e-07 
M2 5 6 4 VPW nch L=4e-08 W=2.5e-07 
M3 1 M1 5 VPW nch L=4e-08 W=2.5e-07 
M4 VSS M1 6 VPW nch L=4e-08 W=2.95e-07 
M5 7 5 VSS VPW nch L=4e-08 W=2.25e-07 
M6 VSS 5 7 VPW nch L=4e-08 W=2.25e-07 
M7 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M8 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M9 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M10 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M11 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M12 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M13 9 M2 VSS VPW nch L=4e-08 W=1.75e-07 
M14 VSS M1 10 VPW nch L=4e-08 W=2.45e-07 
M15 10 M0 VSS VPW nch L=4e-08 W=2.45e-07 
M16 11 9 10 VPW nch L=4e-08 W=2.45e-07 
M17 12 11 VSS VPW nch L=4e-08 W=2.25e-07 
M18 VSS 11 12 VPW nch L=4e-08 W=2.25e-07 
M19 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M20 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M21 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M22 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M23 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M24 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M25 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M26 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M27 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M28 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M29 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M30 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M31 15 16 VSS VPW nch L=4e-08 W=2.25e-07 
M32 VSS 16 15 VPW nch L=4e-08 W=2.25e-07 
M33 17 M2 16 VPW nch L=4e-08 W=2.3e-07 
M34 VSS 4 17 VPW nch L=4e-08 W=2.3e-07 
M35 17 6 VSS VPW nch L=4e-08 W=2.3e-07 
M36 VDD 4 1 VNW pch L=4e-08 W=3.2e-07 
M37 4 M0 VDD VNW pch L=4e-08 W=3.2e-07 
M38 5 6 1 VNW pch L=4e-08 W=3.2e-07 
M39 4 M1 5 VNW pch L=4e-08 W=3.2e-07 
M40 VDD M1 6 VNW pch L=4e-08 W=3.8e-07 
M41 7 5 VDD VNW pch L=4e-08 W=2.9e-07 
M42 VDD 5 7 VNW pch L=4e-08 W=2.9e-07 
M43 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M44 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M45 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M46 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M47 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M48 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M49 9 M2 VDD VNW pch L=4e-08 W=2.25e-07 
M50 21 M1 VDD VNW pch L=4e-08 W=3.8e-07 
M51 11 M0 21 VNW pch L=4e-08 W=3.8e-07 
M52 VDD 9 11 VNW pch L=4e-08 W=2e-07 
M53 12 11 VDD VNW pch L=4e-08 W=2.9e-07 
M54 VDD 11 12 VNW pch L=4e-08 W=2.9e-07 
M55 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M56 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M57 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M58 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M59 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M60 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M61 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M62 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M63 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M64 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M65 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M66 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M67 15 16 VDD VNW pch L=4e-08 W=2.9e-07 
M68 VDD 16 15 VNW pch L=4e-08 W=2.9e-07 
M69 16 M2 VDD VNW pch L=4e-08 W=2e-07 
M70 22 4 16 VNW pch L=4e-08 W=3.5e-07 
M71 VDD 6 22 VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT BENC_X8M_A9TR AN SN X2 VDD VNW VPW VSS M0 M1 M2
M0 VSS 4 1 VPW nch L=4e-08 W=2.8e-07 
M1 4 M0 VSS VPW nch L=4e-08 W=2.8e-07 
M2 5 6 4 VPW nch L=4e-08 W=2.8e-07 
M3 1 M1 5 VPW nch L=4e-08 W=2.8e-07 
M4 VSS M1 6 VPW nch L=4e-08 W=2.95e-07 
M5 7 5 VSS VPW nch L=4e-08 W=2.7e-07 
M6 VSS 5 7 VPW nch L=4e-08 W=2.7e-07 
M7 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M8 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M9 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M10 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M11 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M12 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M13 X2 7 VSS VPW nch L=4e-08 W=2.95e-07 
M14 VSS 7 X2 VPW nch L=4e-08 W=2.95e-07 
M15 9 M2 VSS VPW nch L=4e-08 W=1.75e-07 
M16 VSS M1 10 VPW nch L=4e-08 W=2.45e-07 
M17 10 M0 VSS VPW nch L=4e-08 W=2.45e-07 
M18 11 9 10 VPW nch L=4e-08 W=2.45e-07 
M19 12 11 VSS VPW nch L=4e-08 W=2.7e-07 
M20 VSS 11 12 VPW nch L=4e-08 W=2.7e-07 
M21 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M22 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M23 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M24 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M25 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M26 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M27 AN 12 VSS VPW nch L=4e-08 W=2.95e-07 
M28 VSS 12 AN VPW nch L=4e-08 W=2.95e-07 
M29 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M30 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M31 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M32 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M33 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M34 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M35 SN 15 VSS VPW nch L=4e-08 W=2.95e-07 
M36 VSS 15 SN VPW nch L=4e-08 W=2.95e-07 
M37 15 16 VSS VPW nch L=4e-08 W=2.7e-07 
M38 VSS 16 15 VPW nch L=4e-08 W=2.7e-07 
M39 17 M2 16 VPW nch L=4e-08 W=2.3e-07 
M40 VSS 4 17 VPW nch L=4e-08 W=2.3e-07 
M41 17 6 VSS VPW nch L=4e-08 W=2.3e-07 
M42 VDD 4 1 VNW pch L=4e-08 W=3.6e-07 
M43 4 M0 VDD VNW pch L=4e-08 W=3.6e-07 
M44 5 6 1 VNW pch L=4e-08 W=3.6e-07 
M45 4 M1 5 VNW pch L=4e-08 W=3.6e-07 
M46 VDD M1 6 VNW pch L=4e-08 W=3.8e-07 
M47 7 5 VDD VNW pch L=4e-08 W=3.5e-07 
M48 VDD 5 7 VNW pch L=4e-08 W=3.5e-07 
M49 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M50 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M51 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M52 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M53 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M54 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M55 X2 7 VDD VNW pch L=4e-08 W=3.8e-07 
M56 VDD 7 X2 VNW pch L=4e-08 W=3.8e-07 
M57 9 M2 VDD VNW pch L=4e-08 W=2.25e-07 
M58 21 M1 VDD VNW pch L=4e-08 W=3.8e-07 
M59 11 M0 21 VNW pch L=4e-08 W=3.8e-07 
M60 VDD 9 11 VNW pch L=4e-08 W=2e-07 
M61 12 11 VDD VNW pch L=4e-08 W=3.5e-07 
M62 VDD 11 12 VNW pch L=4e-08 W=3.5e-07 
M63 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M64 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M65 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M66 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M67 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M68 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M69 AN 12 VDD VNW pch L=4e-08 W=3.8e-07 
M70 VDD 12 AN VNW pch L=4e-08 W=3.8e-07 
M71 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M72 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M73 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M74 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M75 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M76 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M77 SN 15 VDD VNW pch L=4e-08 W=3.8e-07 
M78 VDD 15 SN VNW pch L=4e-08 W=3.8e-07 
M79 15 16 VDD VNW pch L=4e-08 W=3.5e-07 
M80 VDD 16 15 VNW pch L=4e-08 W=3.5e-07 
M81 16 M2 VDD VNW pch L=4e-08 W=2e-07 
M82 22 4 16 VNW pch L=4e-08 W=3.5e-07 
M83 VDD 6 22 VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT BMXIT_X0P7M_A9TR PPN VDD VNW VPW VSS AN D0 D1 SN X2
M0 3 SN VSS VPW nch L=4e-08 W=1.35e-07 
M1 5 6 3 VPW nch L=4e-08 W=1.35e-07 
M2 4 D1 5 VPW nch L=4e-08 W=1.35e-07 
M3 VSS D1 6 VPW nch L=4e-08 W=1.35e-07 
M4 7 D0 VSS VPW nch L=4e-08 W=1.35e-07 
M5 8 D0 4 VPW nch L=4e-08 W=1.35e-07 
M6 3 7 8 VPW nch L=4e-08 W=1.35e-07 
M7 4 AN VSS VPW nch L=4e-08 W=1.35e-07 
M8 9 X2 VSS VPW nch L=4e-08 W=1.35e-07 
M9 10 X2 8 VPW nch L=4e-08 W=1.35e-07 
M10 5 9 10 VPW nch L=4e-08 W=1.35e-07 
M11 PPN 10 VSS VPW nch L=4e-08 W=2.6e-07 
M12 3 SN VDD VNW pch L=4e-08 W=2.6e-07 
M13 5 6 4 VNW pch L=4e-08 W=2.6e-07 
M14 3 D1 5 VNW pch L=4e-08 W=2.6e-07 
M15 VDD D1 6 VNW pch L=4e-08 W=2.6e-07 
M16 7 D0 VDD VNW pch L=4e-08 W=2.6e-07 
M17 8 D0 3 VNW pch L=4e-08 W=2.6e-07 
M18 4 7 8 VNW pch L=4e-08 W=2.6e-07 
M19 4 AN VDD VNW pch L=4e-08 W=2.6e-07 
M20 9 X2 VDD VNW pch L=4e-08 W=2.6e-07 
M21 10 X2 5 VNW pch L=4e-08 W=2.6e-07 
M22 8 9 10 VNW pch L=4e-08 W=2.6e-07 
M23 PPN 10 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BMXIT_X1M_A9TR PPN VDD VNW VPW VSS AN D0 D1 SN X2
M0 3 SN VSS VPW nch L=4e-08 W=1.7e-07 
M1 5 6 3 VPW nch L=4e-08 W=1.7e-07 
M2 4 D1 5 VPW nch L=4e-08 W=1.7e-07 
M3 VSS D1 6 VPW nch L=4e-08 W=1.7e-07 
M4 7 D0 VSS VPW nch L=4e-08 W=1.7e-07 
M5 8 D0 4 VPW nch L=4e-08 W=1.7e-07 
M6 3 7 8 VPW nch L=4e-08 W=1.7e-07 
M7 4 AN VSS VPW nch L=4e-08 W=1.7e-07 
M8 9 X2 VSS VPW nch L=4e-08 W=1.7e-07 
M9 10 X2 8 VPW nch L=4e-08 W=1.7e-07 
M10 5 9 10 VPW nch L=4e-08 W=1.7e-07 
M11 PPN 10 VSS VPW nch L=4e-08 W=3.65e-07 
M12 3 SN VDD VNW pch L=4e-08 W=3.3e-07 
M13 5 6 4 VNW pch L=4e-08 W=3.3e-07 
M14 3 D1 5 VNW pch L=4e-08 W=3.3e-07 
M15 VDD D1 6 VNW pch L=4e-08 W=3.3e-07 
M16 7 D0 VDD VNW pch L=4e-08 W=3.3e-07 
M17 8 D0 3 VNW pch L=4e-08 W=3.3e-07 
M18 4 7 8 VNW pch L=4e-08 W=3.3e-07 
M19 4 AN VDD VNW pch L=4e-08 W=3.3e-07 
M20 9 X2 VDD VNW pch L=4e-08 W=3.3e-07 
M21 10 X2 5 VNW pch L=4e-08 W=3.3e-07 
M22 8 9 10 VNW pch L=4e-08 W=3.3e-07 
M23 PPN 10 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT BMXIT_X1P4M_A9TR PPN VDD VNW VPW VSS AN D0 D1 SN X2
M0 3 SN VSS VPW nch L=4e-08 W=1.9e-07 
M1 5 6 3 VPW nch L=4e-08 W=1.9e-07 
M2 4 D1 5 VPW nch L=4e-08 W=1.9e-07 
M3 VSS D1 6 VPW nch L=4e-08 W=1.9e-07 
M4 7 D0 VSS VPW nch L=4e-08 W=1.9e-07 
M5 8 D0 4 VPW nch L=4e-08 W=1.9e-07 
M6 3 7 8 VPW nch L=4e-08 W=1.9e-07 
M7 4 AN VSS VPW nch L=4e-08 W=1.9e-07 
M8 9 X2 VSS VPW nch L=4e-08 W=1.9e-07 
M9 10 X2 8 VPW nch L=4e-08 W=1.9e-07 
M10 5 9 10 VPW nch L=4e-08 W=1.9e-07 
M11 PPN 10 VSS VPW nch L=4e-08 W=2.6e-07 
M12 VSS 10 PPN VPW nch L=4e-08 W=2.6e-07 
M13 3 SN VDD VNW pch L=4e-08 W=3.8e-07 
M14 5 6 4 VNW pch L=4e-08 W=3.8e-07 
M15 3 D1 5 VNW pch L=4e-08 W=3.8e-07 
M16 VDD D1 6 VNW pch L=4e-08 W=3.8e-07 
M17 7 D0 VDD VNW pch L=4e-08 W=3.8e-07 
M18 8 D0 3 VNW pch L=4e-08 W=3.8e-07 
M19 4 7 8 VNW pch L=4e-08 W=3.8e-07 
M20 4 AN VDD VNW pch L=4e-08 W=3.8e-07 
M21 9 X2 VDD VNW pch L=4e-08 W=3.8e-07 
M22 10 X2 5 VNW pch L=4e-08 W=3.8e-07 
M23 8 9 10 VNW pch L=4e-08 W=3.8e-07 
M24 PPN 10 VDD VNW pch L=4e-08 W=2.85e-07 
M25 VDD 10 PPN VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BMXIT_X2M_A9TR PPN VDD VNW VPW VSS AN D0 D1 SN X2
M0 3 SN VSS VPW nch L=4e-08 W=1.9e-07 
M1 5 6 3 VPW nch L=4e-08 W=1.9e-07 
M2 4 D1 5 VPW nch L=4e-08 W=1.9e-07 
M3 VSS D1 6 VPW nch L=4e-08 W=1.9e-07 
M4 7 D0 VSS VPW nch L=4e-08 W=1.9e-07 
M5 8 D0 4 VPW nch L=4e-08 W=1.9e-07 
M6 3 7 8 VPW nch L=4e-08 W=1.9e-07 
M7 4 AN VSS VPW nch L=4e-08 W=1.9e-07 
M8 9 X2 VSS VPW nch L=4e-08 W=1.9e-07 
M9 10 X2 8 VPW nch L=4e-08 W=1.9e-07 
M10 5 9 10 VPW nch L=4e-08 W=1.9e-07 
M11 PPN 10 VSS VPW nch L=4e-08 W=3.65e-07 
M12 VSS 10 PPN VPW nch L=4e-08 W=3.65e-07 
M13 3 SN VDD VNW pch L=4e-08 W=3.8e-07 
M14 5 6 4 VNW pch L=4e-08 W=3.8e-07 
M15 3 D1 5 VNW pch L=4e-08 W=3.8e-07 
M16 VDD D1 6 VNW pch L=4e-08 W=3.8e-07 
M17 7 D0 VDD VNW pch L=4e-08 W=3.8e-07 
M18 8 D0 3 VNW pch L=4e-08 W=3.8e-07 
M19 4 7 8 VNW pch L=4e-08 W=3.8e-07 
M20 4 AN VDD VNW pch L=4e-08 W=3.8e-07 
M21 9 X2 VDD VNW pch L=4e-08 W=3.8e-07 
M22 10 X2 5 VNW pch L=4e-08 W=3.8e-07 
M23 8 9 10 VNW pch L=4e-08 W=3.8e-07 
M24 PPN 10 VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD 10 PPN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT BMXT_X0P7M_A9TR PP VDD VNW VPW VSS AN D0 D1 SN X2
M0 VSS SN 1 VPW nch L=4e-08 W=1.6e-07 
M1 4 6 VSS VPW nch L=4e-08 W=1.6e-07 
M2 6 7 1 VPW nch L=4e-08 W=1.6e-07 
M3 5 D1 6 VPW nch L=4e-08 W=1.6e-07 
M4 VSS D1 7 VPW nch L=4e-08 W=1.6e-07 
M5 8 D0 VSS VPW nch L=4e-08 W=1.6e-07 
M6 9 D0 5 VPW nch L=4e-08 W=1.6e-07 
M7 1 8 9 VPW nch L=4e-08 W=1.6e-07 
M8 10 9 VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS AN 5 VPW nch L=4e-08 W=1.6e-07 
M10 11 X2 VSS VPW nch L=4e-08 W=1.6e-07 
M11 12 X2 10 VPW nch L=4e-08 W=1.6e-07 
M12 4 11 12 VPW nch L=4e-08 W=1.6e-07 
M13 PP 12 VSS VPW nch L=4e-08 W=2.2e-07 
M14 VDD SN 1 VNW pch L=4e-08 W=2.65e-07 
M15 4 6 VDD VNW pch L=4e-08 W=2.05e-07 
M16 6 7 5 VNW pch L=4e-08 W=2.65e-07 
M17 1 D1 6 VNW pch L=4e-08 W=2.65e-07 
M18 VDD D1 7 VNW pch L=4e-08 W=2.65e-07 
M19 8 D0 VDD VNW pch L=4e-08 W=2.65e-07 
M20 9 D0 1 VNW pch L=4e-08 W=2.65e-07 
M21 5 8 9 VNW pch L=4e-08 W=2.65e-07 
M22 10 9 VDD VNW pch L=4e-08 W=2.05e-07 
M23 VDD AN 5 VNW pch L=4e-08 W=2.65e-07 
M24 11 X2 VDD VNW pch L=4e-08 W=2.05e-07 
M25 12 X2 4 VNW pch L=4e-08 W=2.05e-07 
M26 10 11 12 VNW pch L=4e-08 W=2.05e-07 
M27 PP 12 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BMXT_X1M_A9TR PP VDD VNW VPW VSS AN D0 D1 SN X2
M0 VSS SN 1 VPW nch L=4e-08 W=1.9e-07 
M1 4 6 VSS VPW nch L=4e-08 W=1.9e-07 
M2 6 7 1 VPW nch L=4e-08 W=1.9e-07 
M3 5 D1 6 VPW nch L=4e-08 W=1.9e-07 
M4 VSS D1 7 VPW nch L=4e-08 W=1.9e-07 
M5 8 D0 VSS VPW nch L=4e-08 W=1.9e-07 
M6 9 D0 5 VPW nch L=4e-08 W=1.9e-07 
M7 1 8 9 VPW nch L=4e-08 W=1.9e-07 
M8 10 9 VSS VPW nch L=4e-08 W=1.9e-07 
M9 VSS AN 5 VPW nch L=4e-08 W=1.9e-07 
M10 11 X2 VSS VPW nch L=4e-08 W=1.9e-07 
M11 12 X2 10 VPW nch L=4e-08 W=1.9e-07 
M12 4 11 12 VPW nch L=4e-08 W=1.9e-07 
M13 PP 12 VSS VPW nch L=4e-08 W=2.95e-07 
M14 VDD SN 1 VNW pch L=4e-08 W=3.15e-07 
M15 4 6 VDD VNW pch L=4e-08 W=2.5e-07 
M16 6 7 5 VNW pch L=4e-08 W=3.15e-07 
M17 1 D1 6 VNW pch L=4e-08 W=3.15e-07 
M18 VDD D1 7 VNW pch L=4e-08 W=3.15e-07 
M19 8 D0 VDD VNW pch L=4e-08 W=3.15e-07 
M20 9 D0 1 VNW pch L=4e-08 W=3.15e-07 
M21 5 8 9 VNW pch L=4e-08 W=3.15e-07 
M22 10 9 VDD VNW pch L=4e-08 W=2.5e-07 
M23 VDD AN 5 VNW pch L=4e-08 W=3.15e-07 
M24 11 X2 VDD VNW pch L=4e-08 W=2.5e-07 
M25 12 X2 4 VNW pch L=4e-08 W=2.5e-07 
M26 10 11 12 VNW pch L=4e-08 W=2.5e-07 
M27 PP 12 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT BMXT_X1P4M_A9TR PP VDD VNW VPW VSS AN D0 D1 SN X2
M0 VSS SN 1 VPW nch L=4e-08 W=2.4e-07 
M1 4 6 VSS VPW nch L=4e-08 W=2.4e-07 
M2 6 7 1 VPW nch L=4e-08 W=2.4e-07 
M3 5 D1 6 VPW nch L=4e-08 W=2.4e-07 
M4 VSS D1 7 VPW nch L=4e-08 W=2.4e-07 
M5 8 D0 VSS VPW nch L=4e-08 W=2.4e-07 
M6 9 D0 5 VPW nch L=4e-08 W=2.4e-07 
M7 1 8 9 VPW nch L=4e-08 W=2.4e-07 
M8 10 9 VSS VPW nch L=4e-08 W=2.4e-07 
M9 VSS AN 5 VPW nch L=4e-08 W=2.4e-07 
M10 11 X2 VSS VPW nch L=4e-08 W=2.4e-07 
M11 12 X2 10 VPW nch L=4e-08 W=2.4e-07 
M12 4 11 12 VPW nch L=4e-08 W=2.4e-07 
M13 PP 12 VSS VPW nch L=4e-08 W=2.2e-07 
M14 VSS 12 PP VPW nch L=4e-08 W=2.2e-07 
M15 VDD SN 1 VNW pch L=4e-08 W=3.8e-07 
M16 4 6 VDD VNW pch L=4e-08 W=3.1e-07 
M17 6 7 5 VNW pch L=4e-08 W=3.8e-07 
M18 1 D1 6 VNW pch L=4e-08 W=3.8e-07 
M19 VDD D1 7 VNW pch L=4e-08 W=3.8e-07 
M20 8 D0 VDD VNW pch L=4e-08 W=3.8e-07 
M21 9 D0 1 VNW pch L=4e-08 W=3.8e-07 
M22 5 8 9 VNW pch L=4e-08 W=3.8e-07 
M23 10 9 VDD VNW pch L=4e-08 W=3.1e-07 
M24 VDD AN 5 VNW pch L=4e-08 W=3.8e-07 
M25 11 X2 VDD VNW pch L=4e-08 W=3.1e-07 
M26 12 X2 4 VNW pch L=4e-08 W=3.1e-07 
M27 10 11 12 VNW pch L=4e-08 W=3.1e-07 
M28 PP 12 VDD VNW pch L=4e-08 W=2.85e-07 
M29 VDD 12 PP VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BMXT_X2M_A9TR PP VDD VNW VPW VSS AN D0 D1 SN X2
M0 VSS SN 1 VPW nch L=4e-08 W=2.4e-07 
M1 4 6 VSS VPW nch L=4e-08 W=2.4e-07 
M2 6 7 1 VPW nch L=4e-08 W=2.4e-07 
M3 5 D1 6 VPW nch L=4e-08 W=2.4e-07 
M4 VSS D1 7 VPW nch L=4e-08 W=2.4e-07 
M5 8 D0 VSS VPW nch L=4e-08 W=2.4e-07 
M6 9 D0 5 VPW nch L=4e-08 W=2.4e-07 
M7 1 8 9 VPW nch L=4e-08 W=2.4e-07 
M8 10 9 VSS VPW nch L=4e-08 W=2.4e-07 
M9 VSS AN 5 VPW nch L=4e-08 W=2.4e-07 
M10 11 X2 VSS VPW nch L=4e-08 W=2.4e-07 
M11 12 X2 10 VPW nch L=4e-08 W=2.4e-07 
M12 4 11 12 VPW nch L=4e-08 W=2.4e-07 
M13 PP 12 VSS VPW nch L=4e-08 W=2.95e-07 
M14 VSS 12 PP VPW nch L=4e-08 W=2.95e-07 
M15 VDD SN 1 VNW pch L=4e-08 W=3.8e-07 
M16 4 6 VDD VNW pch L=4e-08 W=3.1e-07 
M17 6 7 5 VNW pch L=4e-08 W=3.8e-07 
M18 1 D1 6 VNW pch L=4e-08 W=3.8e-07 
M19 VDD D1 7 VNW pch L=4e-08 W=3.8e-07 
M20 8 D0 VDD VNW pch L=4e-08 W=3.8e-07 
M21 9 D0 1 VNW pch L=4e-08 W=3.8e-07 
M22 5 8 9 VNW pch L=4e-08 W=3.8e-07 
M23 10 9 VDD VNW pch L=4e-08 W=3.1e-07 
M24 VDD AN 5 VNW pch L=4e-08 W=3.8e-07 
M25 11 X2 VDD VNW pch L=4e-08 W=3.1e-07 
M26 12 X2 4 VNW pch L=4e-08 W=3.1e-07 
M27 10 11 12 VNW pch L=4e-08 W=3.1e-07 
M28 PP 12 VDD VNW pch L=4e-08 W=3.8e-07 
M29 VDD 12 PP VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT BUFH_X0P7M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.5e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M2 VDD A 1 VNW pch L=4e-08 W=1.95e-07 
M3 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BUFH_X0P8M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.7e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M2 VDD A 1 VNW pch L=4e-08 W=2.2e-07 
M3 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BUFH_X11M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.85e-07 
M1 1 A VSS VPW nch L=4e-08 W=2.85e-07 
M2 VSS A 1 VPW nch L=4e-08 W=2.85e-07 
M3 1 A VSS VPW nch L=4e-08 W=2.85e-07 
M4 VSS A 1 VPW nch L=4e-08 W=2.85e-07 
M5 1 A VSS VPW nch L=4e-08 W=2.85e-07 
M6 VSS A 1 VPW nch L=4e-08 W=2.85e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M13 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M15 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M17 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M18 VDD A 1 VNW pch L=4e-08 W=3.7e-07 
M19 1 A VDD VNW pch L=4e-08 W=3.7e-07 
M20 VDD A 1 VNW pch L=4e-08 W=3.7e-07 
M21 1 A VDD VNW pch L=4e-08 W=3.7e-07 
M22 VDD A 1 VNW pch L=4e-08 W=3.7e-07 
M23 1 A VDD VNW pch L=4e-08 W=3.7e-07 
M24 VDD A 1 VNW pch L=4e-08 W=3.7e-07 
M25 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M27 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M29 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M31 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M33 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M35 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFH_X13M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.95e-07 
M1 VSS A 3 VPW nch L=4e-08 W=2.95e-07 
M2 3 A VSS VPW nch L=4e-08 W=2.95e-07 
M3 VSS A 3 VPW nch L=4e-08 W=2.95e-07 
M4 3 A VSS VPW nch L=4e-08 W=2.95e-07 
M5 VSS A 3 VPW nch L=4e-08 W=2.95e-07 
M6 3 A VSS VPW nch L=4e-08 W=2.95e-07 
M7 VSS A 3 VPW nch L=4e-08 W=2.95e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M10 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M12 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M16 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M18 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M20 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M21 3 A VDD VNW pch L=4e-08 W=3.8e-07 
M22 VDD A 3 VNW pch L=4e-08 W=3.8e-07 
M23 3 A VDD VNW pch L=4e-08 W=3.8e-07 
M24 VDD A 3 VNW pch L=4e-08 W=3.8e-07 
M25 3 A VDD VNW pch L=4e-08 W=3.8e-07 
M26 VDD A 3 VNW pch L=4e-08 W=3.8e-07 
M27 3 A VDD VNW pch L=4e-08 W=3.8e-07 
M28 VDD A 3 VNW pch L=4e-08 W=3.8e-07 
M29 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M31 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M33 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M35 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M37 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M39 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M41 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFH_X16M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M13 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M15 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M17 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M18 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M19 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M20 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M21 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M22 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M23 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M24 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M25 VDD A 1 VNW pch L=4e-08 W=4e-07 
M26 1 A VDD VNW pch L=4e-08 W=4e-07 
M27 VDD A 1 VNW pch L=4e-08 W=4e-07 
M28 1 A VDD VNW pch L=4e-08 W=4e-07 
M29 VDD A 1 VNW pch L=4e-08 W=4e-07 
M30 1 A VDD VNW pch L=4e-08 W=4e-07 
M31 VDD A 1 VNW pch L=4e-08 W=4e-07 
M32 1 A VDD VNW pch L=4e-08 W=4e-07 
M33 VDD A 1 VNW pch L=4e-08 W=4e-07 
M34 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M36 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M38 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M40 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M41 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M42 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M43 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M44 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M45 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M46 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M47 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M48 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M49 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFH_X1M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.95e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VDD A 1 VNW pch L=4e-08 W=2.55e-07 
M3 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFH_X1P2M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.35e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.85e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=1.85e-07 
M3 VDD A 1 VNW pch L=4e-08 W=3e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=2.4e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT BUFH_X1P4M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.7e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.2e-07 
M3 VDD A 1 VNW pch L=4e-08 W=3.45e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BUFH_X1P7M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M3 VDD A 1 VNW pch L=4e-08 W=3.95e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BUFH_X2M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=1.85e-07 
M1 VSS A 3 VPW nch L=4e-08 W=1.85e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M4 3 A VDD VNW pch L=4e-08 W=2.4e-07 
M5 VDD A 3 VNW pch L=4e-08 W=2.4e-07 
M6 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M7 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFH_X2P5M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.3e-07 
M1 VSS A 3 VPW nch L=4e-08 W=2.3e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=2.6e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=2.6e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=2.6e-07 
M5 3 A VDD VNW pch L=4e-08 W=3e-07 
M6 VDD A 3 VNW pch L=4e-08 W=3e-07 
M7 Y 3 VDD VNW pch L=4e-08 W=3.35e-07 
M8 VDD 3 Y VNW pch L=4e-08 W=3.35e-07 
M9 Y 3 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BUFH_X3M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.7e-07 
M1 VSS A 3 VPW nch L=4e-08 W=2.7e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M5 3 A VDD VNW pch L=4e-08 W=3.45e-07 
M6 VDD A 3 VNW pch L=4e-08 W=3.45e-07 
M7 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M8 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M9 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFH_X3P5M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A 3 VPW nch L=4e-08 W=3.1e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=2.7e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=2.7e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=2.7e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=2.7e-07 
M6 3 A VDD VNW pch L=4e-08 W=4e-07 
M7 VDD A 3 VNW pch L=4e-08 W=4e-07 
M8 Y 3 VDD VNW pch L=4e-08 W=3.5e-07 
M9 VDD 3 Y VNW pch L=4e-08 W=3.5e-07 
M10 Y 3 VDD VNW pch L=4e-08 W=3.5e-07 
M11 VDD 3 Y VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT BUFH_X4M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.45e-07 
M1 1 A VSS VPW nch L=4e-08 W=2.45e-07 
M2 VSS A 1 VPW nch L=4e-08 W=2.45e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M7 VDD A 1 VNW pch L=4e-08 W=3.2e-07 
M8 1 A VDD VNW pch L=4e-08 W=3.2e-07 
M9 VDD A 1 VNW pch L=4e-08 W=3.2e-07 
M10 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M12 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M13 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFH_X5M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=3.05e-07 
M1 1 A VSS VPW nch L=4e-08 W=3.05e-07 
M2 VSS A 1 VPW nch L=4e-08 W=3.05e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VDD A 1 VNW pch L=4e-08 W=3.9e-07 
M9 1 A VDD VNW pch L=4e-08 W=3.9e-07 
M10 VDD A 1 VNW pch L=4e-08 W=3.9e-07 
M11 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M13 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M15 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFH_X6M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.75e-07 
M1 VSS A 3 VPW nch L=4e-08 W=2.75e-07 
M2 3 A VSS VPW nch L=4e-08 W=2.75e-07 
M3 VSS A 3 VPW nch L=4e-08 W=2.75e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M10 3 A VDD VNW pch L=4e-08 W=3.5e-07 
M11 VDD A 3 VNW pch L=4e-08 W=3.5e-07 
M12 3 A VDD VNW pch L=4e-08 W=3.5e-07 
M13 VDD A 3 VNW pch L=4e-08 W=3.5e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M16 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M17 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M18 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFH_X7P5M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.75e-07 
M1 1 A VSS VPW nch L=4e-08 W=2.75e-07 
M2 VSS A 1 VPW nch L=4e-08 W=2.75e-07 
M3 1 A VSS VPW nch L=4e-08 W=2.75e-07 
M4 VSS A 1 VPW nch L=4e-08 W=2.75e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=2.9e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=2.9e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=2.9e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=2.9e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=2.9e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=2.9e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=2.9e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=2.9e-07 
M13 VDD A 1 VNW pch L=4e-08 W=3.55e-07 
M14 1 A VDD VNW pch L=4e-08 W=3.55e-07 
M15 VDD A 1 VNW pch L=4e-08 W=3.55e-07 
M16 1 A VDD VNW pch L=4e-08 W=3.55e-07 
M17 VDD A 1 VNW pch L=4e-08 W=3.55e-07 
M18 Y 1 VDD VNW pch L=4e-08 W=3.75e-07 
M19 VDD 1 Y VNW pch L=4e-08 W=3.75e-07 
M20 Y 1 VDD VNW pch L=4e-08 W=3.75e-07 
M21 VDD 1 Y VNW pch L=4e-08 W=3.75e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=3.75e-07 
M23 VDD 1 Y VNW pch L=4e-08 W=3.75e-07 
M24 Y 1 VDD VNW pch L=4e-08 W=3.75e-07 
M25 VDD 1 Y VNW pch L=4e-08 W=3.75e-07 
.ENDS


.SUBCKT BUFH_X9M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 2 VPW nch L=4e-08 W=3.3e-07 
M1 2 A VSS VPW nch L=4e-08 W=3.3e-07 
M2 VSS A 2 VPW nch L=4e-08 W=3.3e-07 
M3 2 A VSS VPW nch L=4e-08 W=3.3e-07 
M4 VSS A 2 VPW nch L=4e-08 W=3.3e-07 
M5 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M7 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M9 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M13 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M14 2 A VDD VNW pch L=4e-08 W=3.55e-07 
M15 VDD A 2 VNW pch L=4e-08 W=3.55e-07 
M16 2 A VDD VNW pch L=4e-08 W=3.55e-07 
M17 VDD A 2 VNW pch L=4e-08 W=3.55e-07 
M18 2 A VDD VNW pch L=4e-08 W=3.55e-07 
M19 VDD A 2 VNW pch L=4e-08 W=3.55e-07 
M20 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M22 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M24 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M26 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M28 Y 2 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUFZ_X11M_A9TR Y VDD VNW VPW VSS A OE
M0 2 OE 1 VPW nch L=4e-08 W=2.5e-07 
M1 1 OE 2 VPW nch L=4e-08 W=2.5e-07 
M2 2 OE 1 VPW nch L=4e-08 W=2.5e-07 
M3 1 A VSS VPW nch L=4e-08 W=2.85e-07 
M4 VSS A 1 VPW nch L=4e-08 W=2.85e-07 
M5 1 A VSS VPW nch L=4e-08 W=2.85e-07 
M6 VSS A 1 VPW nch L=4e-08 W=2.85e-07 
M7 1 A VSS VPW nch L=4e-08 W=2.85e-07 
M8 VSS A 1 VPW nch L=4e-08 W=2.85e-07 
M9 5 OE VSS VPW nch L=4e-08 W=2.85e-07 
M10 VSS OE 5 VPW nch L=4e-08 W=2.85e-07 
M11 5 OE VSS VPW nch L=4e-08 W=2.85e-07 
M12 VSS 5 1 VPW nch L=4e-08 W=2.4e-07 
M13 1 5 VSS VPW nch L=4e-08 W=2.4e-07 
M14 VSS 5 1 VPW nch L=4e-08 W=2.4e-07 
M15 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M16 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M17 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M18 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M19 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M20 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M21 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M22 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M23 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M24 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M25 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M26 2 5 1 VNW pch L=4e-08 W=3.15e-07 
M27 1 5 2 VNW pch L=4e-08 W=3.15e-07 
M28 2 5 1 VNW pch L=4e-08 W=3.15e-07 
M29 2 A VDD VNW pch L=4e-08 W=3.65e-07 
M30 VDD A 2 VNW pch L=4e-08 W=3.65e-07 
M31 2 A VDD VNW pch L=4e-08 W=3.65e-07 
M32 VDD A 2 VNW pch L=4e-08 W=3.65e-07 
M33 2 A VDD VNW pch L=4e-08 W=3.65e-07 
M34 VDD A 2 VNW pch L=4e-08 W=3.65e-07 
M35 5 OE VDD VNW pch L=4e-08 W=3.65e-07 
M36 VDD OE 5 VNW pch L=4e-08 W=3.65e-07 
M37 5 OE VDD VNW pch L=4e-08 W=3.65e-07 
M38 VDD OE 2 VNW pch L=4e-08 W=3.65e-07 
M39 2 OE VDD VNW pch L=4e-08 W=3.65e-07 
M40 VDD OE 2 VNW pch L=4e-08 W=3.65e-07 
M41 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
M42 VDD 2 Y VNW pch L=4e-08 W=3.4e-07 
M43 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
M44 VDD 2 Y VNW pch L=4e-08 W=3.4e-07 
M45 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
M46 VDD 2 Y VNW pch L=4e-08 W=3.4e-07 
M47 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
M48 VDD 2 Y VNW pch L=4e-08 W=3.4e-07 
M49 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
M50 VDD 2 Y VNW pch L=4e-08 W=3.4e-07 
M51 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
.ENDS


.SUBCKT BUFZ_X16M_A9TR Y VDD VNW VPW VSS A OE
M0 2 OE 1 VPW nch L=4e-08 W=2.5e-07 
M1 1 OE 2 VPW nch L=4e-08 W=2.5e-07 
M2 2 OE 1 VPW nch L=4e-08 W=2.5e-07 
M3 1 OE 2 VPW nch L=4e-08 W=2.5e-07 
M4 2 OE 1 VPW nch L=4e-08 W=2.5e-07 
M5 VSS OE 3 VPW nch L=4e-08 W=3.8e-07 
M6 3 OE VSS VPW nch L=4e-08 W=3.8e-07 
M7 VSS OE 3 VPW nch L=4e-08 W=3.8e-07 
M8 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M10 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M12 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M14 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M16 1 3 VSS VPW nch L=4e-08 W=2.4e-07 
M17 VSS 3 1 VPW nch L=4e-08 W=2.4e-07 
M18 1 3 VSS VPW nch L=4e-08 W=2.4e-07 
M19 VSS 3 1 VPW nch L=4e-08 W=2.4e-07 
M20 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M21 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M22 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M23 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M24 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M25 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M26 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M27 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M28 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M29 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M30 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M31 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M32 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M33 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M34 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M35 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M36 2 3 1 VNW pch L=4e-08 W=3.15e-07 
M37 1 3 2 VNW pch L=4e-08 W=3.15e-07 
M38 2 3 1 VNW pch L=4e-08 W=3.15e-07 
M39 1 3 2 VNW pch L=4e-08 W=3.15e-07 
M40 2 3 1 VNW pch L=4e-08 W=3.15e-07 
M41 VDD OE 3 VNW pch L=4e-08 W=3.8e-07 
M42 3 OE VDD VNW pch L=4e-08 W=3.8e-07 
M43 VDD OE 3 VNW pch L=4e-08 W=3.8e-07 
M44 2 A VDD VNW pch L=4e-08 W=3.8e-07 
M45 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M46 2 A VDD VNW pch L=4e-08 W=3.8e-07 
M47 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M48 2 A VDD VNW pch L=4e-08 W=3.8e-07 
M49 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M50 2 A VDD VNW pch L=4e-08 W=3.8e-07 
M51 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M52 2 OE VDD VNW pch L=4e-08 W=3.8e-07 
M53 VDD OE 2 VNW pch L=4e-08 W=3.8e-07 
M54 2 OE VDD VNW pch L=4e-08 W=3.8e-07 
M55 VDD OE 2 VNW pch L=4e-08 W=3.8e-07 
M56 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M57 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M58 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M59 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M60 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M61 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M62 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M63 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M64 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M65 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M66 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M67 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M68 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M69 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M70 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M71 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
.ENDS


.SUBCKT BUFZ_X1M_A9TR Y VDD VNW VPW VSS A OE
M0 2 OE 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A 1 VPW nch L=4e-08 W=1.55e-07 
M2 5 OE VSS VPW nch L=4e-08 W=2.25e-07 
M3 VSS 5 1 VPW nch L=4e-08 W=1.2e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.55e-07 
M5 VSS 1 Y VPW nch L=4e-08 W=1.55e-07 
M6 2 5 1 VNW pch L=4e-08 W=1.55e-07 
M7 VDD A 2 VNW pch L=4e-08 W=2e-07 
M8 5 OE VDD VNW pch L=4e-08 W=2.95e-07 
M9 VDD OE 2 VNW pch L=4e-08 W=1.55e-07 
M10 Y 2 VDD VNW pch L=4e-08 W=2e-07 
M11 VDD 2 Y VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT BUFZ_X1P4M_A9TR Y VDD VNW VPW VSS A OE
M0 2 OE 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A 1 VPW nch L=4e-08 W=2.2e-07 
M2 5 OE VSS VPW nch L=4e-08 W=2.25e-07 
M3 VSS 5 1 VPW nch L=4e-08 W=1.2e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M5 VSS 1 Y VPW nch L=4e-08 W=2.2e-07 
M6 2 5 1 VNW pch L=4e-08 W=1.55e-07 
M7 VDD A 2 VNW pch L=4e-08 W=2.85e-07 
M8 5 OE VDD VNW pch L=4e-08 W=2.95e-07 
M9 VDD OE 2 VNW pch L=4e-08 W=1.55e-07 
M10 Y 2 VDD VNW pch L=4e-08 W=2.85e-07 
M11 VDD 2 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BUFZ_X2M_A9TR Y VDD VNW VPW VSS A OE
M0 2 OE 1 VPW nch L=4e-08 W=1.55e-07 
M1 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M2 5 OE VSS VPW nch L=4e-08 W=2.4e-07 
M3 VSS 5 1 VPW nch L=4e-08 W=1.55e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M5 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M6 2 5 1 VNW pch L=4e-08 W=2e-07 
M7 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M8 5 OE VDD VNW pch L=4e-08 W=3.1e-07 
M9 VDD OE 2 VNW pch L=4e-08 W=2e-07 
M10 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M11 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
.ENDS


.SUBCKT BUFZ_X3M_A9TR Y VDD VNW VPW VSS A OE
M0 2 OE 1 VPW nch L=4e-08 W=2.35e-07 
M1 1 A VSS VPW nch L=4e-08 W=2.35e-07 
M2 VSS A 1 VPW nch L=4e-08 W=2.35e-07 
M3 5 OE VSS VPW nch L=4e-08 W=2.8e-07 
M4 VSS 5 1 VPW nch L=4e-08 W=2.35e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M8 2 5 1 VNW pch L=4e-08 W=3e-07 
M9 2 A VDD VNW pch L=4e-08 W=3e-07 
M10 VDD A 2 VNW pch L=4e-08 W=3e-07 
M11 5 OE VDD VNW pch L=4e-08 W=3.6e-07 
M12 VDD OE 2 VNW pch L=4e-08 W=3e-07 
M13 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M14 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M15 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
.ENDS


.SUBCKT BUFZ_X4M_A9TR Y VDD VNW VPW VSS A OE
M0 2 OE 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M3 5 OE VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS 5 1 VPW nch L=4e-08 W=2.6e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M9 2 5 1 VNW pch L=4e-08 W=3.1e-07 
M10 2 A VDD VNW pch L=4e-08 W=3.8e-07 
M11 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M12 5 OE VDD VNW pch L=4e-08 W=3.8e-07 
M13 VDD OE 2 VNW pch L=4e-08 W=4e-07 
M14 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M15 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M16 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M17 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
.ENDS


.SUBCKT BUFZ_X6M_A9TR Y VDD VNW VPW VSS A OE
M0 2 OE 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 OE 2 VPW nch L=4e-08 W=2.4e-07 
M2 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M5 5 OE VSS VPW nch L=4e-08 W=2.35e-07 
M6 VSS OE 5 VPW nch L=4e-08 W=2.35e-07 
M7 1 5 VSS VPW nch L=4e-08 W=2.35e-07 
M8 VSS 5 1 VPW nch L=4e-08 W=2.35e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M13 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M14 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M15 2 5 1 VNW pch L=4e-08 W=3e-07 
M16 1 5 2 VNW pch L=4e-08 W=3e-07 
M17 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M18 2 A VDD VNW pch L=4e-08 W=3.8e-07 
M19 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M20 5 OE VDD VNW pch L=4e-08 W=3e-07 
M21 VDD OE 5 VNW pch L=4e-08 W=3e-07 
M22 2 OE VDD VNW pch L=4e-08 W=3e-07 
M23 VDD OE 2 VNW pch L=4e-08 W=3e-07 
M24 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M25 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M26 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M27 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
M28 Y 2 VDD VNW pch L=4e-08 W=3.6e-07 
M29 VDD 2 Y VNW pch L=4e-08 W=3.6e-07 
.ENDS


.SUBCKT BUFZ_X8M_A9TR Y VDD VNW VPW VSS A OE
M0 2 OE 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 OE 2 VPW nch L=4e-08 W=3.1e-07 
M2 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M4 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M5 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M6 5 OE VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS OE 5 VPW nch L=4e-08 W=3.1e-07 
M8 1 5 VSS VPW nch L=4e-08 W=2.6e-07 
M9 VSS 5 1 VPW nch L=4e-08 W=2.6e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M11 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M13 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M14 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M15 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M16 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M17 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M18 2 5 1 VNW pch L=4e-08 W=3.1e-07 
M19 1 5 2 VNW pch L=4e-08 W=3.1e-07 
M20 2 A VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M22 2 A VDD VNW pch L=4e-08 W=3.8e-07 
M23 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M24 5 OE VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD OE 5 VNW pch L=4e-08 W=3.8e-07 
M26 2 OE VDD VNW pch L=4e-08 W=4e-07 
M27 VDD OE 2 VNW pch L=4e-08 W=4e-07 
M28 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
M29 VDD 2 Y VNW pch L=4e-08 W=3.4e-07 
M30 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
M31 VDD 2 Y VNW pch L=4e-08 W=3.4e-07 
M32 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
M33 VDD 2 Y VNW pch L=4e-08 W=3.4e-07 
M34 Y 2 VDD VNW pch L=4e-08 W=3.4e-07 
M35 VDD 2 Y VNW pch L=4e-08 W=3.4e-07 
.ENDS


.SUBCKT BUF_X0P7B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M2 VDD A 1 VNW pch L=4e-08 W=2.1e-07 
M3 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BUF_X0P7M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M2 VDD A 1 VNW pch L=4e-08 W=1.55e-07 
M3 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BUF_X0P8B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.9e-07 
M2 VDD A 1 VNW pch L=4e-08 W=2.1e-07 
M3 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BUF_X0P8M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M2 VDD A 1 VNW pch L=4e-08 W=1.55e-07 
M3 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BUF_X11B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.25e-07 
M1 1 A VSS VPW nch L=4e-08 W=2.25e-07 
M2 VSS A 1 VPW nch L=4e-08 W=2.25e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M13 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M14 VDD A 1 VNW pch L=4e-08 W=4e-07 
M15 1 A VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A 1 VNW pch L=4e-08 W=4e-07 
M17 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M19 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M21 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M23 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M25 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M27 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X11M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A 1 VPW nch L=4e-08 W=3.1e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M13 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VDD A 1 VNW pch L=4e-08 W=4e-07 
M15 1 A VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A 1 VNW pch L=4e-08 W=4e-07 
M17 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M19 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M21 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M23 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M25 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M27 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X13B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 2 VPW nch L=4e-08 W=2.8e-07 
M1 2 A VSS VPW nch L=4e-08 W=2.8e-07 
M2 VSS A 2 VPW nch L=4e-08 W=2.8e-07 
M3 Y 2 VSS VPW nch L=4e-08 W=2.25e-07 
M4 VSS 2 Y VPW nch L=4e-08 W=2.25e-07 
M5 Y 2 VSS VPW nch L=4e-08 W=2.25e-07 
M6 VSS 2 Y VPW nch L=4e-08 W=2.25e-07 
M7 Y 2 VSS VPW nch L=4e-08 W=2.25e-07 
M8 VSS 2 Y VPW nch L=4e-08 W=2.25e-07 
M9 Y 2 VSS VPW nch L=4e-08 W=2.25e-07 
M10 VSS 2 Y VPW nch L=4e-08 W=2.25e-07 
M11 Y 2 VSS VPW nch L=4e-08 W=2.25e-07 
M12 VSS 2 Y VPW nch L=4e-08 W=2.25e-07 
M13 Y 2 VSS VPW nch L=4e-08 W=2.25e-07 
M14 VSS 2 Y VPW nch L=4e-08 W=2.25e-07 
M15 Y 2 VSS VPW nch L=4e-08 W=2.25e-07 
M16 2 A VDD VNW pch L=4e-08 W=3.7e-07 
M17 VDD A 2 VNW pch L=4e-08 W=3.7e-07 
M18 2 A VDD VNW pch L=4e-08 W=3.7e-07 
M19 VDD A 2 VNW pch L=4e-08 W=3.7e-07 
M20 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M22 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M24 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M26 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M28 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M30 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M32 Y 2 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X13M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 2 VPW nch L=4e-08 W=3.8e-07 
M1 2 A VSS VPW nch L=4e-08 W=3.8e-07 
M2 VSS A 2 VPW nch L=4e-08 W=3.8e-07 
M3 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M5 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M7 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M9 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M13 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M15 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M16 2 A VDD VNW pch L=4e-08 W=3.65e-07 
M17 VDD A 2 VNW pch L=4e-08 W=3.65e-07 
M18 2 A VDD VNW pch L=4e-08 W=3.65e-07 
M19 VDD A 2 VNW pch L=4e-08 W=3.65e-07 
M20 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M22 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M24 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M26 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M28 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M30 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M32 Y 2 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X16B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=3.5e-07 
M1 1 A VSS VPW nch L=4e-08 W=3.5e-07 
M2 VSS A 1 VPW nch L=4e-08 W=3.5e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M13 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M14 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M15 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M16 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M17 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M18 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M19 VDD A 1 VNW pch L=4e-08 W=3.65e-07 
M20 1 A VDD VNW pch L=4e-08 W=3.65e-07 
M21 VDD A 1 VNW pch L=4e-08 W=3.65e-07 
M22 1 A VDD VNW pch L=4e-08 W=3.65e-07 
M23 VDD A 1 VNW pch L=4e-08 W=3.65e-07 
M24 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M26 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M28 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M30 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M32 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M33 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M34 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M36 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M38 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X16M_A9TR Y VDD VNW VPW VSS A
M0 1 A VSS VPW nch L=4e-08 W=3.5e-07 
M1 VSS A 1 VPW nch L=4e-08 W=3.5e-07 
M2 1 A VSS VPW nch L=4e-08 W=3.5e-07 
M3 VSS A 1 VPW nch L=4e-08 W=3.5e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M5 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M16 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M18 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M20 VDD A 1 VNW pch L=4e-08 W=3.6e-07 
M21 1 A VDD VNW pch L=4e-08 W=3.6e-07 
M22 VDD A 1 VNW pch L=4e-08 W=3.6e-07 
M23 1 A VDD VNW pch L=4e-08 W=3.6e-07 
M24 VDD A 1 VNW pch L=4e-08 W=3.6e-07 
M25 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M27 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M29 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M31 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M33 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M35 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M37 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M39 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X1B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M2 VDD A 1 VNW pch L=4e-08 W=2.1e-07 
M3 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X1M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VDD A 1 VNW pch L=4e-08 W=1.55e-07 
M3 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X1P2B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.35e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=1.35e-07 
M3 VDD A 1 VNW pch L=4e-08 W=2.1e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=2.4e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT BUF_X1P2M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.85e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=1.85e-07 
M3 VDD A 1 VNW pch L=4e-08 W=1.55e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=2.4e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT BUF_X1P4B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M3 VDD A 1 VNW pch L=4e-08 W=2.1e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BUF_X1P4M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.35e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.2e-07 
M3 VDD A 1 VNW pch L=4e-08 W=1.75e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT BUF_X1P7B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.9e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=1.9e-07 
M3 VDD A 1 VNW pch L=4e-08 W=2.1e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BUF_X1P7M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.55e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M3 VDD A 1 VNW pch L=4e-08 W=2e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BUF_X2B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.35e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M3 VDD A 1 VNW pch L=4e-08 W=2.35e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X2M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.8e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M3 VDD A 1 VNW pch L=4e-08 W=2.3e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X2P5B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.65e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.9e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=1.9e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=1.9e-07 
M4 VDD A 1 VNW pch L=4e-08 W=2.95e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
M6 VDD 1 Y VNW pch L=4e-08 W=3.35e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BUF_X2P5M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.25e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.6e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.6e-07 
M4 VDD A 1 VNW pch L=4e-08 W=2.9e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
M6 VDD 1 Y VNW pch L=4e-08 W=3.35e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT BUF_X3B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.95e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M4 VDD A 1 VNW pch L=4e-08 W=3.4e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M6 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X3M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.6e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VDD A 1 VNW pch L=4e-08 W=3.4e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M6 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X3P5B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.25e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=2e-07 
M5 VDD A 1 VNW pch L=4e-08 W=4e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=3.5e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=3.5e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=3.5e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT BUF_X3P5M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=3.05e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.7e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.7e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.7e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=2.7e-07 
M5 VDD A 1 VNW pch L=4e-08 W=3.95e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=3.5e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=3.5e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=3.5e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT BUF_X4B_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=1.3e-07 
M1 VSS A 3 VPW nch L=4e-08 W=1.3e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=2.25e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=2.25e-07 
M6 3 A VDD VNW pch L=4e-08 W=2.3e-07 
M7 VDD A 3 VNW pch L=4e-08 W=2.3e-07 
M8 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M9 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M10 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X4M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=1.75e-07 
M1 VSS A 3 VPW nch L=4e-08 W=1.75e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M6 3 A VDD VNW pch L=4e-08 W=2.3e-07 
M7 VDD A 3 VNW pch L=4e-08 W=2.3e-07 
M8 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M9 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M10 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X5B_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS A 3 VPW nch L=4e-08 W=1.6e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=2.25e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=2.25e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M7 3 A VDD VNW pch L=4e-08 W=2.85e-07 
M8 VDD A 3 VNW pch L=4e-08 W=2.85e-07 
M9 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M11 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M13 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X5M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS A 3 VPW nch L=4e-08 W=2.2e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M7 3 A VDD VNW pch L=4e-08 W=2.8e-07 
M8 VDD A 3 VNW pch L=4e-08 W=2.8e-07 
M9 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M11 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M13 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X6B_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=1.95e-07 
M1 VSS A 3 VPW nch L=4e-08 W=1.95e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=2.25e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=2.25e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=2.25e-07 
M8 3 A VDD VNW pch L=4e-08 W=3.4e-07 
M9 VDD A 3 VNW pch L=4e-08 W=3.4e-07 
M10 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M12 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M13 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X6M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.6e-07 
M1 VSS A 3 VPW nch L=4e-08 W=2.6e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M8 3 A VDD VNW pch L=4e-08 W=3.35e-07 
M9 VDD A 3 VNW pch L=4e-08 W=3.35e-07 
M10 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M11 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M12 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M13 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X7P5B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.65e-07 
M1 1 A VSS VPW nch L=4e-08 W=1.65e-07 
M2 VSS A 1 VPW nch L=4e-08 W=1.65e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.15e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=2.15e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=2.15e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=2.15e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=2.15e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=2.15e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=2.15e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=2.15e-07 
M11 VDD A 1 VNW pch L=4e-08 W=2.95e-07 
M12 1 A VDD VNW pch L=4e-08 W=2.95e-07 
M13 VDD A 1 VNW pch L=4e-08 W=2.95e-07 
M14 Y 1 VDD VNW pch L=4e-08 W=3.75e-07 
M15 VDD 1 Y VNW pch L=4e-08 W=3.75e-07 
M16 Y 1 VDD VNW pch L=4e-08 W=3.75e-07 
M17 VDD 1 Y VNW pch L=4e-08 W=3.75e-07 
M18 Y 1 VDD VNW pch L=4e-08 W=3.75e-07 
M19 VDD 1 Y VNW pch L=4e-08 W=3.75e-07 
M20 Y 1 VDD VNW pch L=4e-08 W=3.75e-07 
M21 VDD 1 Y VNW pch L=4e-08 W=3.75e-07 
.ENDS


.SUBCKT BUF_X7P5M_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A 3 VPW nch L=4e-08 W=3.1e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=2.9e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=2.9e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=2.9e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=2.9e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=2.9e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=2.9e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=2.9e-07 
M9 VSS 3 Y VPW nch L=4e-08 W=2.9e-07 
M10 3 A VDD VNW pch L=4e-08 W=4e-07 
M11 VDD A 3 VNW pch L=4e-08 W=4e-07 
M12 Y 3 VDD VNW pch L=4e-08 W=3.75e-07 
M13 VDD 3 Y VNW pch L=4e-08 W=3.75e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=3.75e-07 
M15 VDD 3 Y VNW pch L=4e-08 W=3.75e-07 
M16 Y 3 VDD VNW pch L=4e-08 W=3.75e-07 
M17 VDD 3 Y VNW pch L=4e-08 W=3.75e-07 
M18 Y 3 VDD VNW pch L=4e-08 W=3.75e-07 
M19 VDD 3 Y VNW pch L=4e-08 W=3.75e-07 
.ENDS


.SUBCKT BUF_X9B_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=1.95e-07 
M1 1 A VSS VPW nch L=4e-08 W=1.95e-07 
M2 VSS A 1 VPW nch L=4e-08 W=1.95e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=2.25e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=2.25e-07 
M12 VDD A 1 VNW pch L=4e-08 W=3.45e-07 
M13 1 A VDD VNW pch L=4e-08 W=3.45e-07 
M14 VDD A 1 VNW pch L=4e-08 W=3.45e-07 
M15 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M17 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M19 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M21 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M23 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT BUF_X9M_A9TR Y VDD VNW VPW VSS A
M0 VSS A 1 VPW nch L=4e-08 W=2.65e-07 
M1 1 A VSS VPW nch L=4e-08 W=2.65e-07 
M2 VSS A 1 VPW nch L=4e-08 W=2.65e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VDD A 1 VNW pch L=4e-08 W=3.4e-07 
M13 1 A VDD VNW pch L=4e-08 W=3.4e-07 
M14 VDD A 1 VNW pch L=4e-08 W=3.4e-07 
M15 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M17 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M19 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M21 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M23 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT CGENCIN_X1M_A9TR CO VDD VNW VPW VSS A B CIN
M0 VSS 4 1 VPW nch L=4e-08 W=2.6e-07 
M1 4 A VSS VPW nch L=4e-08 W=2.6e-07 
M2 5 B 4 VPW nch L=4e-08 W=2.6e-07 
M3 1 7 5 VPW nch L=4e-08 W=2.6e-07 
M4 6 7 4 VPW nch L=4e-08 W=2.6e-07 
M5 1 B 6 VPW nch L=4e-08 W=2.6e-07 
M6 VSS B 7 VPW nch L=4e-08 W=3.6e-07 
M7 8 7 VSS VPW nch L=4e-08 W=2.6e-07 
M8 CO 5 9 VPW nch L=4e-08 W=2.6e-07 
M9 8 6 CO VPW nch L=4e-08 W=2.6e-07 
M10 9 CIN VSS VPW nch L=4e-08 W=2.6e-07 
M11 VDD 4 1 VNW pch L=4e-08 W=3.15e-07 
M12 4 A VDD VNW pch L=4e-08 W=3.15e-07 
M13 5 B 1 VNW pch L=4e-08 W=3.15e-07 
M14 4 7 5 VNW pch L=4e-08 W=3.15e-07 
M15 6 7 1 VNW pch L=4e-08 W=3.15e-07 
M16 4 B 6 VNW pch L=4e-08 W=3.15e-07 
M17 VDD B 7 VNW pch L=4e-08 W=4e-07 
M18 8 7 VDD VNW pch L=4e-08 W=4e-07 
M19 CO 5 8 VNW pch L=4e-08 W=4e-07 
M20 9 6 CO VNW pch L=4e-08 W=4e-07 
M21 9 CIN VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT CGENCIN_X1P4M_A9TR CO VDD VNW VPW VSS A B CIN
M0 VSS 4 1 VPW nch L=4e-08 W=3.3e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.3e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.3e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.3e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.3e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.3e-07 
M6 7 B VSS VPW nch L=4e-08 W=2.75e-07 
M7 VSS B 7 VPW nch L=4e-08 W=2.75e-07 
M8 8 7 VSS VPW nch L=4e-08 W=1.85e-07 
M9 VSS 7 8 VPW nch L=4e-08 W=1.85e-07 
M10 10 5 CO VPW nch L=4e-08 W=1.85e-07 
M11 CO 5 10 VPW nch L=4e-08 W=1.85e-07 
M12 8 6 CO VPW nch L=4e-08 W=2.4e-07 
M13 CO 6 8 VPW nch L=4e-08 W=1.3e-07 
M14 10 CIN VSS VPW nch L=4e-08 W=1.85e-07 
M15 VSS CIN 10 VPW nch L=4e-08 W=1.85e-07 
M16 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M17 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M18 5 B 1 VNW pch L=4e-08 W=4e-07 
M19 4 7 5 VNW pch L=4e-08 W=4e-07 
M20 6 7 1 VNW pch L=4e-08 W=4e-07 
M21 4 B 6 VNW pch L=4e-08 W=4e-07 
M22 7 B VDD VNW pch L=4e-08 W=2.85e-07 
M23 VDD B 7 VNW pch L=4e-08 W=2.85e-07 
M24 8 7 VDD VNW pch L=4e-08 W=2.85e-07 
M25 VDD 7 8 VNW pch L=4e-08 W=2.85e-07 
M26 8 5 CO VNW pch L=4e-08 W=2.85e-07 
M27 CO 5 8 VNW pch L=4e-08 W=2.85e-07 
M28 10 6 CO VNW pch L=4e-08 W=2.85e-07 
M29 CO 6 10 VNW pch L=4e-08 W=2.85e-07 
M30 10 CIN VDD VNW pch L=4e-08 W=2.85e-07 
M31 VDD CIN 10 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT CGENCIN_X2M_A9TR CO VDD VNW VPW VSS A B CIN
M0 VSS 4 1 VPW nch L=4e-08 W=3.3e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.3e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.3e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.3e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.3e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.3e-07 
M6 7 B VSS VPW nch L=4e-08 W=3.8e-07 
M7 VSS B 7 VPW nch L=4e-08 W=3.8e-07 
M8 8 7 VSS VPW nch L=4e-08 W=2.6e-07 
M9 VSS 7 8 VPW nch L=4e-08 W=2.6e-07 
M10 10 5 CO VPW nch L=4e-08 W=2.6e-07 
M11 CO 5 10 VPW nch L=4e-08 W=2.6e-07 
M12 8 6 CO VPW nch L=4e-08 W=3.9e-07 
M13 CO 6 8 VPW nch L=4e-08 W=1.3e-07 
M14 10 CIN VSS VPW nch L=4e-08 W=2.6e-07 
M15 VSS CIN 10 VPW nch L=4e-08 W=2.6e-07 
M16 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M17 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M18 5 B 1 VNW pch L=4e-08 W=4e-07 
M19 4 7 5 VNW pch L=4e-08 W=4e-07 
M20 6 7 1 VNW pch L=4e-08 W=4e-07 
M21 4 B 6 VNW pch L=4e-08 W=4e-07 
M22 7 B VDD VNW pch L=4e-08 W=4e-07 
M23 VDD B 7 VNW pch L=4e-08 W=4e-07 
M24 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD 7 8 VNW pch L=4e-08 W=3.8e-07 
M26 8 5 CO VNW pch L=4e-08 W=4e-07 
M27 CO 5 8 VNW pch L=4e-08 W=4e-07 
M28 10 6 CO VNW pch L=4e-08 W=4e-07 
M29 CO 6 10 VNW pch L=4e-08 W=4e-07 
M30 10 CIN VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD CIN 10 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT CGENCON_X1M_A9TR CON VDD VNW VPW VSS A B CI
M0 VSS 4 1 VPW nch L=4e-08 W=2.6e-07 
M1 4 A VSS VPW nch L=4e-08 W=2.6e-07 
M2 5 B 4 VPW nch L=4e-08 W=2.6e-07 
M3 1 7 5 VPW nch L=4e-08 W=2.6e-07 
M4 6 7 4 VPW nch L=4e-08 W=2.6e-07 
M5 1 B 6 VPW nch L=4e-08 W=2.6e-07 
M6 7 B VSS VPW nch L=4e-08 W=2.6e-07 
M7 CON 5 8 VPW nch L=4e-08 W=2.6e-07 
M8 7 6 CON VPW nch L=4e-08 W=2.6e-07 
M9 8 CI VSS VPW nch L=4e-08 W=2.6e-07 
M10 VDD 4 1 VNW pch L=4e-08 W=3.15e-07 
M11 4 A VDD VNW pch L=4e-08 W=3.15e-07 
M12 5 B 1 VNW pch L=4e-08 W=3.15e-07 
M13 4 7 5 VNW pch L=4e-08 W=3.15e-07 
M14 6 7 1 VNW pch L=4e-08 W=3.15e-07 
M15 4 B 6 VNW pch L=4e-08 W=3.15e-07 
M16 VDD B 7 VNW pch L=4e-08 W=3.8e-07 
M17 CON 5 7 VNW pch L=4e-08 W=4e-07 
M18 8 6 CON VNW pch L=4e-08 W=4e-07 
M19 8 CI VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT CGENCON_X1P4M_A9TR CON VDD VNW VPW VSS A B CI
M0 VSS 4 1 VPW nch L=4e-08 W=3.3e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.3e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.3e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.3e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.3e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.3e-07 
M6 VSS B 7 VPW nch L=4e-08 W=3.7e-07 
M7 CON 5 9 VPW nch L=4e-08 W=3.7e-07 
M8 7 6 CON VPW nch L=4e-08 W=3.7e-07 
M9 9 CI VSS VPW nch L=4e-08 W=1.85e-07 
M10 VSS CI 9 VPW nch L=4e-08 W=1.85e-07 
M11 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M12 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M13 5 B 1 VNW pch L=4e-08 W=4e-07 
M14 4 7 5 VNW pch L=4e-08 W=4e-07 
M15 6 7 1 VNW pch L=4e-08 W=4e-07 
M16 4 B 6 VNW pch L=4e-08 W=4e-07 
M17 7 B VDD VNW pch L=4e-08 W=2.85e-07 
M18 VDD B 7 VNW pch L=4e-08 W=2.85e-07 
M19 7 5 CON VNW pch L=4e-08 W=2.85e-07 
M20 CON 5 7 VNW pch L=4e-08 W=2.85e-07 
M21 9 6 CON VNW pch L=4e-08 W=2.85e-07 
M22 CON 6 9 VNW pch L=4e-08 W=2.85e-07 
M23 9 CI VDD VNW pch L=4e-08 W=2.85e-07 
M24 VDD CI 9 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT CGENCON_X2M_A9TR CON VDD VNW VPW VSS A B CI
M0 VSS 4 1 VPW nch L=4e-08 W=1.9e-07 
M1 4 A VSS VPW nch L=4e-08 W=3.3e-07 
M2 5 B 4 VPW nch L=4e-08 W=3.3e-07 
M3 1 7 5 VPW nch L=4e-08 W=3.3e-07 
M4 6 7 4 VPW nch L=4e-08 W=3.3e-07 
M5 1 B 6 VPW nch L=4e-08 W=3.3e-07 
M6 7 B VSS VPW nch L=4e-08 W=2.6e-07 
M7 VSS B 7 VPW nch L=4e-08 W=2.6e-07 
M8 9 5 CON VPW nch L=4e-08 W=2.6e-07 
M9 CON 5 9 VPW nch L=4e-08 W=2.6e-07 
M10 7 6 CON VPW nch L=4e-08 W=2.6e-07 
M11 CON 6 7 VPW nch L=4e-08 W=2.6e-07 
M12 9 CI VSS VPW nch L=4e-08 W=2.6e-07 
M13 VSS CI 9 VPW nch L=4e-08 W=2.6e-07 
M14 VDD 4 1 VNW pch L=4e-08 W=3.8e-07 
M15 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M16 5 B 1 VNW pch L=4e-08 W=3.9e-07 
M17 4 7 5 VNW pch L=4e-08 W=3.9e-07 
M18 6 7 1 VNW pch L=4e-08 W=3.9e-07 
M19 4 B 6 VNW pch L=4e-08 W=3.9e-07 
M20 7 B VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD B 7 VNW pch L=4e-08 W=3.8e-07 
M22 7 5 CON VNW pch L=4e-08 W=4e-07 
M23 CON 5 7 VNW pch L=4e-08 W=4e-07 
M24 9 6 CON VNW pch L=4e-08 W=4e-07 
M25 CON 6 9 VNW pch L=4e-08 W=4e-07 
M26 9 CI VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD CI 9 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT CGENI_X1M_A9TR CON VDD VNW VPW VSS A B CI
M0 3 A VSS VPW nch L=4e-08 W=2.4e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.4e-07 
M2 10 B VSS VPW nch L=4e-08 W=2.4e-07 
M3 CON A 10 VPW nch L=4e-08 W=2.4e-07 
M4 3 CI CON VPW nch L=4e-08 W=2.4e-07 
M5 4 A VDD VNW pch L=4e-08 W=4e-07 
M6 VDD B 4 VNW pch L=4e-08 W=4e-07 
M7 9 B VDD VNW pch L=4e-08 W=4e-07 
M8 CON A 9 VNW pch L=4e-08 W=4e-07 
M9 4 CI CON VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT CGENI_X1P4M_A9TR CON VDD VNW VPW VSS A B CI
M0 11 A CON VPW nch L=4e-08 W=1.7e-07 
M1 VSS B 11 VPW nch L=4e-08 W=1.7e-07 
M2 4 B VSS VPW nch L=4e-08 W=1.7e-07 
M3 VSS A 4 VPW nch L=4e-08 W=1.7e-07 
M4 4 A VSS VPW nch L=4e-08 W=1.7e-07 
M5 VSS B 4 VPW nch L=4e-08 W=1.7e-07 
M6 12 B VSS VPW nch L=4e-08 W=1.7e-07 
M7 CON A 12 VPW nch L=4e-08 W=1.7e-07 
M8 4 CI CON VPW nch L=4e-08 W=1.7e-07 
M9 CON CI 4 VPW nch L=4e-08 W=1.7e-07 
M10 9 A CON VNW pch L=4e-08 W=2.85e-07 
M11 VDD B 9 VNW pch L=4e-08 W=2.85e-07 
M12 5 B VDD VNW pch L=4e-08 W=2.85e-07 
M13 VDD A 5 VNW pch L=4e-08 W=2.85e-07 
M14 5 A VDD VNW pch L=4e-08 W=2.85e-07 
M15 VDD B 5 VNW pch L=4e-08 W=2.85e-07 
M16 10 B VDD VNW pch L=4e-08 W=2.85e-07 
M17 CON A 10 VNW pch L=4e-08 W=2.85e-07 
M18 5 CI CON VNW pch L=4e-08 W=2.85e-07 
M19 CON CI 5 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT CGENI_X2M_A9TR CON VDD VNW VPW VSS A B CI
M0 11 A CON VPW nch L=4e-08 W=2.3e-07 
M1 VSS B 11 VPW nch L=4e-08 W=2.3e-07 
M2 4 B VSS VPW nch L=4e-08 W=2.3e-07 
M3 VSS A 4 VPW nch L=4e-08 W=2.3e-07 
M4 4 A VSS VPW nch L=4e-08 W=2.3e-07 
M5 VSS B 4 VPW nch L=4e-08 W=2.3e-07 
M6 12 B VSS VPW nch L=4e-08 W=2.3e-07 
M7 CON A 12 VPW nch L=4e-08 W=2.3e-07 
M8 4 CI CON VPW nch L=4e-08 W=2.3e-07 
M9 CON CI 4 VPW nch L=4e-08 W=2.3e-07 
M10 9 A CON VNW pch L=4e-08 W=3.8e-07 
M11 VDD B 9 VNW pch L=4e-08 W=3.8e-07 
M12 5 B VDD VNW pch L=4e-08 W=3.8e-07 
M13 VDD A 5 VNW pch L=4e-08 W=3.8e-07 
M14 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M15 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M16 10 B VDD VNW pch L=4e-08 W=3.8e-07 
M17 CON A 10 VNW pch L=4e-08 W=3.8e-07 
M18 5 CI CON VNW pch L=4e-08 W=3.8e-07 
M19 CON CI 5 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT CGEN_X1M_A9TR CO VDD VNW VPW VSS A B CI
M0 3 CI 1 VPW nch L=4e-08 W=2.3e-07 
M1 11 A 3 VPW nch L=4e-08 W=2.3e-07 
M2 VSS B 11 VPW nch L=4e-08 W=2.3e-07 
M3 1 B VSS VPW nch L=4e-08 W=2.3e-07 
M4 VSS A 1 VPW nch L=4e-08 W=2.3e-07 
M5 CO 3 VSS VPW nch L=4e-08 W=3.1e-07 
M6 3 CI 2 VNW pch L=4e-08 W=3.8e-07 
M7 10 A 3 VNW pch L=4e-08 W=3.8e-07 
M8 VDD B 10 VNW pch L=4e-08 W=3.8e-07 
M9 2 B VDD VNW pch L=4e-08 W=3.8e-07 
M10 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M11 CO 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT CGEN_X1P4M_A9TR CO VDD VNW VPW VSS A B CI
M0 3 CI 1 VPW nch L=4e-08 W=2.3e-07 
M1 11 A 3 VPW nch L=4e-08 W=2.3e-07 
M2 VSS B 11 VPW nch L=4e-08 W=2.3e-07 
M3 1 B VSS VPW nch L=4e-08 W=2.3e-07 
M4 VSS A 1 VPW nch L=4e-08 W=2.3e-07 
M5 CO 3 VSS VPW nch L=4e-08 W=2.2e-07 
M6 VSS 3 CO VPW nch L=4e-08 W=2.2e-07 
M7 3 CI 2 VNW pch L=4e-08 W=3.8e-07 
M8 10 A 3 VNW pch L=4e-08 W=3.8e-07 
M9 VDD B 10 VNW pch L=4e-08 W=3.8e-07 
M10 2 B VDD VNW pch L=4e-08 W=3.8e-07 
M11 VDD A 2 VNW pch L=4e-08 W=3.8e-07 
M12 CO 3 VDD VNW pch L=4e-08 W=2.85e-07 
M13 VDD 3 CO VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT CGEN_X2M_A9TR CO VDD VNW VPW VSS A B CI
M0 12 A 1 VPW nch L=4e-08 W=2.3e-07 
M1 VSS B 12 VPW nch L=4e-08 W=2.3e-07 
M2 4 B VSS VPW nch L=4e-08 W=2.3e-07 
M3 VSS A 4 VPW nch L=4e-08 W=2.3e-07 
M4 4 A VSS VPW nch L=4e-08 W=2.3e-07 
M5 VSS B 4 VPW nch L=4e-08 W=2.3e-07 
M6 13 B VSS VPW nch L=4e-08 W=2.3e-07 
M7 1 A 13 VPW nch L=4e-08 W=2.3e-07 
M8 4 CI 1 VPW nch L=4e-08 W=2.3e-07 
M9 1 CI 4 VPW nch L=4e-08 W=2.3e-07 
M10 CO 1 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 1 CO VPW nch L=4e-08 W=3.1e-07 
M12 10 A 1 VNW pch L=4e-08 W=3.8e-07 
M13 VDD B 10 VNW pch L=4e-08 W=3.8e-07 
M14 5 B VDD VNW pch L=4e-08 W=3.8e-07 
M15 VDD A 5 VNW pch L=4e-08 W=3.8e-07 
M16 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M17 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M18 11 B VDD VNW pch L=4e-08 W=3.8e-07 
M19 1 A 11 VNW pch L=4e-08 W=3.8e-07 
M20 5 CI 1 VNW pch L=4e-08 W=3.8e-07 
M21 1 CI 5 VNW pch L=4e-08 W=3.8e-07 
M22 CO 1 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 1 CO VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT CMPR42_X1M_A9TR CO ICO SUM VDD VNW VPW VSS A B C D ICI
M0 VSS 6 ICO VPW nch L=4e-08 W=3.1e-07 
M1 4 A VSS VPW nch L=4e-08 W=2.2e-07 
M2 VSS B 4 VPW nch L=4e-08 W=2.2e-07 
M3 30 B VSS VPW nch L=4e-08 W=2.2e-07 
M4 6 A 30 VPW nch L=4e-08 W=2.2e-07 
M5 4 C 6 VPW nch L=4e-08 W=2.2e-07 
M6 7 C VSS VPW nch L=4e-08 W=2.35e-07 
M7 VSS A 7 VPW nch L=4e-08 W=2.35e-07 
M8 7 B VSS VPW nch L=4e-08 W=2.35e-07 
M9 9 6 7 VPW nch L=4e-08 W=2.35e-07 
M10 31 C 9 VPW nch L=4e-08 W=1.35e-07 
M11 32 A 31 VPW nch L=4e-08 W=1.35e-07 
M12 VSS B 32 VPW nch L=4e-08 W=1.35e-07 
M13 10 9 VSS VPW nch L=4e-08 W=2.65e-07 
M14 VSS 14 CO VPW nch L=4e-08 W=3.1e-07 
M15 12 ICI VSS VPW nch L=4e-08 W=2.2e-07 
M16 VSS D 12 VPW nch L=4e-08 W=2.2e-07 
M17 33 D VSS VPW nch L=4e-08 W=2.2e-07 
M18 14 ICI 33 VPW nch L=4e-08 W=2.2e-07 
M19 12 10 14 VPW nch L=4e-08 W=2.2e-07 
M20 15 10 VSS VPW nch L=4e-08 W=2.35e-07 
M21 VSS ICI 15 VPW nch L=4e-08 W=2.35e-07 
M22 15 D VSS VPW nch L=4e-08 W=2.35e-07 
M23 17 14 15 VPW nch L=4e-08 W=2.35e-07 
M24 34 10 17 VPW nch L=4e-08 W=1.35e-07 
M25 35 ICI 34 VPW nch L=4e-08 W=1.35e-07 
M26 VSS D 35 VPW nch L=4e-08 W=1.35e-07 
M27 SUM 17 VSS VPW nch L=4e-08 W=3.1e-07 
M28 VDD 6 ICO VNW pch L=4e-08 W=4e-07 
M29 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M31 24 B VDD VNW pch L=4e-08 W=3.8e-07 
M32 6 A 24 VNW pch L=4e-08 W=3.8e-07 
M33 5 C 6 VNW pch L=4e-08 W=3.8e-07 
M34 8 C VDD VNW pch L=4e-08 W=2.55e-07 
M35 VDD A 8 VNW pch L=4e-08 W=2.55e-07 
M36 8 B VDD VNW pch L=4e-08 W=2.55e-07 
M37 9 6 8 VNW pch L=4e-08 W=2.55e-07 
M38 25 C 9 VNW pch L=4e-08 W=2.55e-07 
M39 26 A 25 VNW pch L=4e-08 W=2.55e-07 
M40 VDD B 26 VNW pch L=4e-08 W=2.55e-07 
M41 10 9 VDD VNW pch L=4e-08 W=3.4e-07 
M42 VDD 14 CO VNW pch L=4e-08 W=4e-07 
M43 13 ICI VDD VNW pch L=4e-08 W=3.8e-07 
M44 VDD D 13 VNW pch L=4e-08 W=3.8e-07 
M45 27 D VDD VNW pch L=4e-08 W=3.8e-07 
M46 14 ICI 27 VNW pch L=4e-08 W=3.8e-07 
M47 13 10 14 VNW pch L=4e-08 W=3.8e-07 
M48 16 10 VDD VNW pch L=4e-08 W=2.55e-07 
M49 VDD ICI 16 VNW pch L=4e-08 W=2.55e-07 
M50 16 D VDD VNW pch L=4e-08 W=2.55e-07 
M51 17 14 16 VNW pch L=4e-08 W=2.55e-07 
M52 28 10 17 VNW pch L=4e-08 W=2.55e-07 
M53 29 ICI 28 VNW pch L=4e-08 W=2.55e-07 
M54 VDD D 29 VNW pch L=4e-08 W=2.55e-07 
M55 SUM 17 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT CMPR42_X1P4M_A9TR CO ICO SUM VDD VNW VPW VSS A B C D ICI
M0 ICO 6 VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS 6 ICO VPW nch L=4e-08 W=2.2e-07 
M2 4 A VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS B 4 VPW nch L=4e-08 W=2.2e-07 
M4 30 B VSS VPW nch L=4e-08 W=2.2e-07 
M5 6 A 30 VPW nch L=4e-08 W=2.2e-07 
M6 4 C 6 VPW nch L=4e-08 W=2.2e-07 
M7 7 C VSS VPW nch L=4e-08 W=2.35e-07 
M8 VSS A 7 VPW nch L=4e-08 W=2.35e-07 
M9 7 B VSS VPW nch L=4e-08 W=2.35e-07 
M10 9 6 7 VPW nch L=4e-08 W=2.35e-07 
M11 31 C 9 VPW nch L=4e-08 W=1.35e-07 
M12 32 A 31 VPW nch L=4e-08 W=1.35e-07 
M13 VSS B 32 VPW nch L=4e-08 W=1.35e-07 
M14 10 9 VSS VPW nch L=4e-08 W=2.65e-07 
M15 CO 14 VSS VPW nch L=4e-08 W=2.2e-07 
M16 VSS 14 CO VPW nch L=4e-08 W=2.2e-07 
M17 12 ICI VSS VPW nch L=4e-08 W=2.2e-07 
M18 VSS D 12 VPW nch L=4e-08 W=2.2e-07 
M19 33 D VSS VPW nch L=4e-08 W=2.2e-07 
M20 14 ICI 33 VPW nch L=4e-08 W=2.2e-07 
M21 12 10 14 VPW nch L=4e-08 W=2.2e-07 
M22 15 10 VSS VPW nch L=4e-08 W=2.35e-07 
M23 VSS ICI 15 VPW nch L=4e-08 W=2.35e-07 
M24 15 D VSS VPW nch L=4e-08 W=2.35e-07 
M25 17 14 15 VPW nch L=4e-08 W=2.35e-07 
M26 34 10 17 VPW nch L=4e-08 W=1.35e-07 
M27 35 ICI 34 VPW nch L=4e-08 W=1.35e-07 
M28 VSS D 35 VPW nch L=4e-08 W=1.35e-07 
M29 SUM 17 VSS VPW nch L=4e-08 W=2.2e-07 
M30 VSS 17 SUM VPW nch L=4e-08 W=2.2e-07 
M31 ICO 6 VDD VNW pch L=4e-08 W=2.85e-07 
M32 VDD 6 ICO VNW pch L=4e-08 W=2.85e-07 
M33 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M35 24 B VDD VNW pch L=4e-08 W=3.8e-07 
M36 6 A 24 VNW pch L=4e-08 W=3.8e-07 
M37 5 C 6 VNW pch L=4e-08 W=3.8e-07 
M38 8 C VDD VNW pch L=4e-08 W=2.55e-07 
M39 VDD A 8 VNW pch L=4e-08 W=2.55e-07 
M40 8 B VDD VNW pch L=4e-08 W=2.55e-07 
M41 9 6 8 VNW pch L=4e-08 W=2.55e-07 
M42 25 C 9 VNW pch L=4e-08 W=2.55e-07 
M43 26 A 25 VNW pch L=4e-08 W=2.55e-07 
M44 VDD B 26 VNW pch L=4e-08 W=2.55e-07 
M45 10 9 VDD VNW pch L=4e-08 W=3.4e-07 
M46 CO 14 VDD VNW pch L=4e-08 W=2.85e-07 
M47 VDD 14 CO VNW pch L=4e-08 W=2.85e-07 
M48 13 ICI VDD VNW pch L=4e-08 W=3.8e-07 
M49 VDD D 13 VNW pch L=4e-08 W=3.8e-07 
M50 27 D VDD VNW pch L=4e-08 W=3.8e-07 
M51 14 ICI 27 VNW pch L=4e-08 W=3.8e-07 
M52 13 10 14 VNW pch L=4e-08 W=3.8e-07 
M53 16 10 VDD VNW pch L=4e-08 W=2.55e-07 
M54 VDD ICI 16 VNW pch L=4e-08 W=2.55e-07 
M55 16 D VDD VNW pch L=4e-08 W=2.55e-07 
M56 17 14 16 VNW pch L=4e-08 W=2.55e-07 
M57 28 10 17 VNW pch L=4e-08 W=2.55e-07 
M58 29 ICI 28 VNW pch L=4e-08 W=2.55e-07 
M59 VDD D 29 VNW pch L=4e-08 W=2.55e-07 
M60 SUM 17 VDD VNW pch L=4e-08 W=2.85e-07 
M61 VDD 17 SUM VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT CMPR42_X2M_A9TR CO ICO SUM VDD VNW VPW VSS A B C D ICI
M0 ICO 6 VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS 6 ICO VPW nch L=4e-08 W=3.1e-07 
M2 4 A VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS B 4 VPW nch L=4e-08 W=2.2e-07 
M4 30 B VSS VPW nch L=4e-08 W=2.2e-07 
M5 6 A 30 VPW nch L=4e-08 W=2.2e-07 
M6 4 C 6 VPW nch L=4e-08 W=2.2e-07 
M7 7 C VSS VPW nch L=4e-08 W=2.35e-07 
M8 VSS A 7 VPW nch L=4e-08 W=2.35e-07 
M9 7 B VSS VPW nch L=4e-08 W=2.35e-07 
M10 9 6 7 VPW nch L=4e-08 W=2.35e-07 
M11 31 C 9 VPW nch L=4e-08 W=1.35e-07 
M12 32 A 31 VPW nch L=4e-08 W=1.35e-07 
M13 VSS B 32 VPW nch L=4e-08 W=1.35e-07 
M14 10 9 VSS VPW nch L=4e-08 W=2.65e-07 
M15 CO 14 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 14 CO VPW nch L=4e-08 W=3.1e-07 
M17 12 ICI VSS VPW nch L=4e-08 W=2.2e-07 
M18 VSS D 12 VPW nch L=4e-08 W=2.2e-07 
M19 33 D VSS VPW nch L=4e-08 W=2.2e-07 
M20 14 ICI 33 VPW nch L=4e-08 W=2.2e-07 
M21 12 10 14 VPW nch L=4e-08 W=2.2e-07 
M22 15 10 VSS VPW nch L=4e-08 W=2.35e-07 
M23 VSS ICI 15 VPW nch L=4e-08 W=2.35e-07 
M24 15 D VSS VPW nch L=4e-08 W=2.35e-07 
M25 17 14 15 VPW nch L=4e-08 W=2.35e-07 
M26 34 10 17 VPW nch L=4e-08 W=1.35e-07 
M27 35 ICI 34 VPW nch L=4e-08 W=1.35e-07 
M28 VSS D 35 VPW nch L=4e-08 W=1.35e-07 
M29 SUM 17 VSS VPW nch L=4e-08 W=3.1e-07 
M30 VSS 17 SUM VPW nch L=4e-08 W=3.1e-07 
M31 ICO 6 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 6 ICO VNW pch L=4e-08 W=4e-07 
M33 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M35 24 B VDD VNW pch L=4e-08 W=3.8e-07 
M36 6 A 24 VNW pch L=4e-08 W=3.8e-07 
M37 5 C 6 VNW pch L=4e-08 W=3.8e-07 
M38 8 C VDD VNW pch L=4e-08 W=2.55e-07 
M39 VDD A 8 VNW pch L=4e-08 W=2.55e-07 
M40 8 B VDD VNW pch L=4e-08 W=2.55e-07 
M41 9 6 8 VNW pch L=4e-08 W=2.55e-07 
M42 25 C 9 VNW pch L=4e-08 W=2.55e-07 
M43 26 A 25 VNW pch L=4e-08 W=2.55e-07 
M44 VDD B 26 VNW pch L=4e-08 W=2.55e-07 
M45 10 9 VDD VNW pch L=4e-08 W=3.4e-07 
M46 CO 14 VDD VNW pch L=4e-08 W=4e-07 
M47 VDD 14 CO VNW pch L=4e-08 W=4e-07 
M48 13 ICI VDD VNW pch L=4e-08 W=3.8e-07 
M49 VDD D 13 VNW pch L=4e-08 W=3.8e-07 
M50 27 D VDD VNW pch L=4e-08 W=3.8e-07 
M51 14 ICI 27 VNW pch L=4e-08 W=3.8e-07 
M52 13 10 14 VNW pch L=4e-08 W=3.8e-07 
M53 16 10 VDD VNW pch L=4e-08 W=2.55e-07 
M54 VDD ICI 16 VNW pch L=4e-08 W=2.55e-07 
M55 16 D VDD VNW pch L=4e-08 W=2.55e-07 
M56 17 14 16 VNW pch L=4e-08 W=2.55e-07 
M57 28 10 17 VNW pch L=4e-08 W=2.55e-07 
M58 29 ICI 28 VNW pch L=4e-08 W=2.55e-07 
M59 VDD D 29 VNW pch L=4e-08 W=2.55e-07 
M60 SUM 17 VDD VNW pch L=4e-08 W=4e-07 
M61 VDD 17 SUM VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFNQ_X1M_A9TR Q VDD VNW VPW VSS CKN D
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 CKN VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.2e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.2e-07 
M7 8 4 7 VPW nch L=4e-08 W=1.2e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 8 9 VPW nch L=4e-08 W=2e-07 
M11 Q 9 VSS VPW nch L=4e-08 W=2e-07 
M12 VDD 4 1 VNW pch L=4e-08 W=1.3e-07 
M13 4 CKN VDD VNW pch L=4e-08 W=2.5e-07 
M14 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M15 6 4 5 VNW pch L=4e-08 W=2e-07 
M16 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M18 7 6 VDD VNW pch L=4e-08 W=2e-07 
M19 8 1 7 VNW pch L=4e-08 W=2e-07 
M20 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 8 9 VNW pch L=4e-08 W=2e-07 
M23 Q 9 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFNQ_X2M_A9TR Q VDD VNW VPW VSS CKN D
M0 VSS 4 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 CKN VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.2e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.55e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.55e-07 
M7 8 4 7 VPW nch L=4e-08 W=1.55e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 9 8 VSS VPW nch L=4e-08 W=3.1e-07 
M11 Q 9 VSS VPW nch L=4e-08 W=2e-07 
M12 VSS 9 Q VPW nch L=4e-08 W=2e-07 
M13 VDD 4 1 VNW pch L=4e-08 W=1.4e-07 
M14 4 CKN VDD VNW pch L=4e-08 W=2.7e-07 
M15 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M16 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M17 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M18 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M19 7 6 VDD VNW pch L=4e-08 W=3.1e-07 
M20 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M21 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M23 9 8 VDD VNW pch L=4e-08 W=3.1e-07 
M24 Q 9 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 9 Q VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFNQ_X3M_A9TR Q VDD VNW VPW VSS CKN D
M0 VSS 4 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 CKN VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.2e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.55e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.8e-07 
M7 8 4 7 VPW nch L=4e-08 W=1.55e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 9 8 VSS VPW nch L=4e-08 W=1.9e-07 
M11 VSS 8 9 VPW nch L=4e-08 W=1.9e-07 
M12 Q 9 VSS VPW nch L=4e-08 W=2e-07 
M13 VSS 9 Q VPW nch L=4e-08 W=2e-07 
M14 Q 9 VSS VPW nch L=4e-08 W=2e-07 
M15 VDD 4 1 VNW pch L=4e-08 W=1.4e-07 
M16 4 CKN VDD VNW pch L=4e-08 W=2.7e-07 
M17 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M18 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M19 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M20 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M21 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M22 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M23 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M25 9 8 VDD VNW pch L=4e-08 W=1.9e-07 
M26 VDD 8 9 VNW pch L=4e-08 W=1.9e-07 
M27 Q 9 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 9 Q VNW pch L=4e-08 W=4e-07 
M29 Q 9 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFNSRPQ_X1M_A9TR Q VDD VNW VPW VSS CKN D R SN
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 CKN VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.2e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 20 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 8 20 VPW nch L=4e-08 W=1.2e-07 
M6 7 SN VSS VPW nch L=4e-08 W=1.8e-07 
M7 8 6 7 VPW nch L=4e-08 W=1.8e-07 
M8 7 R 8 VPW nch L=4e-08 W=1.8e-07 
M9 9 4 8 VPW nch L=4e-08 W=1.2e-07 
M10 21 1 9 VPW nch L=4e-08 W=1.6e-07 
M11 22 10 21 VPW nch L=4e-08 W=1.6e-07 
M12 VSS SN 22 VPW nch L=4e-08 W=1.6e-07 
M13 23 R VSS VPW nch L=4e-08 W=1.6e-07 
M14 9 SN 23 VPW nch L=4e-08 W=1.6e-07 
M15 VSS 9 10 VPW nch L=4e-08 W=2e-07 
M16 Q 10 VSS VPW nch L=4e-08 W=2e-07 
M17 VDD 4 1 VNW pch L=4e-08 W=1.3e-07 
M18 4 CKN VDD VNW pch L=4e-08 W=2.5e-07 
M19 5 D VDD VNW pch L=4e-08 W=3.6e-07 
M20 6 4 5 VNW pch L=4e-08 W=2e-07 
M21 16 1 6 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 8 16 VNW pch L=4e-08 W=1.2e-07 
M23 8 SN VDD VNW pch L=4e-08 W=3.6e-07 
M24 17 6 8 VNW pch L=4e-08 W=3.6e-07 
M25 VDD R 17 VNW pch L=4e-08 W=3.6e-07 
M26 9 1 8 VNW pch L=4e-08 W=2e-07 
M27 18 4 9 VNW pch L=4e-08 W=1.6e-07 
M28 19 10 18 VNW pch L=4e-08 W=1.6e-07 
M29 VDD R 19 VNW pch L=4e-08 W=1.6e-07 
M30 9 SN VDD VNW pch L=4e-08 W=1.6e-07 
M31 VDD 9 10 VNW pch L=4e-08 W=2e-07 
M32 Q 10 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFNSRPQ_X2M_A9TR Q VDD VNW VPW VSS CKN D R SN
M0 VSS 4 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 CKN VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.4e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.55e-07 
M4 20 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 8 20 VPW nch L=4e-08 W=1.2e-07 
M6 7 SN VSS VPW nch L=4e-08 W=1.8e-07 
M7 8 6 7 VPW nch L=4e-08 W=1.8e-07 
M8 7 R 8 VPW nch L=4e-08 W=1.8e-07 
M9 9 4 8 VPW nch L=4e-08 W=1.55e-07 
M10 21 1 9 VPW nch L=4e-08 W=1.6e-07 
M11 22 10 21 VPW nch L=4e-08 W=1.6e-07 
M12 VSS SN 22 VPW nch L=4e-08 W=1.6e-07 
M13 23 R VSS VPW nch L=4e-08 W=1.6e-07 
M14 9 SN 23 VPW nch L=4e-08 W=1.6e-07 
M15 VSS 9 10 VPW nch L=4e-08 W=3.1e-07 
M16 Q 10 VSS VPW nch L=4e-08 W=2e-07 
M17 VSS 10 Q VPW nch L=4e-08 W=2e-07 
M18 VDD 4 1 VNW pch L=4e-08 W=1.4e-07 
M19 4 CKN VDD VNW pch L=4e-08 W=2.7e-07 
M20 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M21 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M22 16 1 6 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 8 16 VNW pch L=4e-08 W=1.2e-07 
M24 8 SN VDD VNW pch L=4e-08 W=3.6e-07 
M25 17 6 8 VNW pch L=4e-08 W=3.6e-07 
M26 VDD R 17 VNW pch L=4e-08 W=3.6e-07 
M27 9 1 8 VNW pch L=4e-08 W=3.1e-07 
M28 18 4 9 VNW pch L=4e-08 W=1.6e-07 
M29 19 10 18 VNW pch L=4e-08 W=1.6e-07 
M30 VDD R 19 VNW pch L=4e-08 W=1.6e-07 
M31 9 SN VDD VNW pch L=4e-08 W=1.6e-07 
M32 VDD 9 10 VNW pch L=4e-08 W=3.1e-07 
M33 Q 10 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 10 Q VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFNSRPQ_X3M_A9TR Q VDD VNW VPW VSS CKN D R SN
M0 VSS 4 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 CKN VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.4e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.55e-07 
M4 20 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 8 20 VPW nch L=4e-08 W=1.2e-07 
M6 7 SN VSS VPW nch L=4e-08 W=1.8e-07 
M7 8 6 7 VPW nch L=4e-08 W=1.8e-07 
M8 7 R 8 VPW nch L=4e-08 W=1.8e-07 
M9 9 4 8 VPW nch L=4e-08 W=1.55e-07 
M10 21 1 9 VPW nch L=4e-08 W=1.6e-07 
M11 22 10 21 VPW nch L=4e-08 W=1.6e-07 
M12 VSS SN 22 VPW nch L=4e-08 W=1.6e-07 
M13 23 R VSS VPW nch L=4e-08 W=1.6e-07 
M14 9 SN 23 VPW nch L=4e-08 W=1.6e-07 
M15 VSS 9 10 VPW nch L=4e-08 W=3.8e-07 
M16 Q 10 VSS VPW nch L=4e-08 W=2e-07 
M17 VSS 10 Q VPW nch L=4e-08 W=2e-07 
M18 Q 10 VSS VPW nch L=4e-08 W=2e-07 
M19 VDD 4 1 VNW pch L=4e-08 W=1.4e-07 
M20 4 CKN VDD VNW pch L=4e-08 W=2.7e-07 
M21 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M22 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M23 16 1 6 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 8 16 VNW pch L=4e-08 W=1.2e-07 
M25 8 SN VDD VNW pch L=4e-08 W=3.6e-07 
M26 17 6 8 VNW pch L=4e-08 W=3.6e-07 
M27 VDD R 17 VNW pch L=4e-08 W=3.6e-07 
M28 9 1 8 VNW pch L=4e-08 W=3.1e-07 
M29 18 4 9 VNW pch L=4e-08 W=1.6e-07 
M30 19 10 18 VNW pch L=4e-08 W=1.6e-07 
M31 VDD R 19 VNW pch L=4e-08 W=1.6e-07 
M32 9 SN VDD VNW pch L=4e-08 W=1.6e-07 
M33 VDD 9 10 VNW pch L=4e-08 W=3.8e-07 
M34 Q 10 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 10 Q VNW pch L=4e-08 W=4e-07 
M36 Q 10 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFQN_X0P5M_A9TR QN VDD VNW VPW VSS CK D
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.2e-07 
M7 8 4 7 VPW nch L=4e-08 W=1.2e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M11 QN 8 VSS VPW nch L=4e-08 W=1.55e-07 
M12 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M13 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M14 5 D VDD VNW pch L=4e-08 W=2.6e-07 
M15 6 4 5 VNW pch L=4e-08 W=1.2e-07 
M16 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.8e-07 
M19 8 1 7 VNW pch L=4e-08 W=1.2e-07 
M20 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M23 QN 8 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT DFFQN_X1M_A9TR QN VDD VNW VPW VSS CK D
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.4e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.6e-07 
M7 8 4 7 VPW nch L=4e-08 W=1.6e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M11 QN 8 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M13 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M14 5 D VDD VNW pch L=4e-08 W=3.3e-07 
M15 6 4 5 VNW pch L=4e-08 W=1.6e-07 
M16 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M18 7 6 VDD VNW pch L=4e-08 W=2.3e-07 
M19 8 1 7 VNW pch L=4e-08 W=1.6e-07 
M20 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M23 QN 8 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFQN_X2M_A9TR QN VDD VNW VPW VSS CK D
M0 VSS CK 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=2.5e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2.5e-07 
M7 8 4 7 VPW nch L=4e-08 W=2.5e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M11 QN 8 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 8 QN VPW nch L=4e-08 W=3.1e-07 
M13 VDD CK 1 VNW pch L=4e-08 W=1.4e-07 
M14 4 1 VDD VNW pch L=4e-08 W=2.7e-07 
M15 5 D VDD VNW pch L=4e-08 W=3.2e-07 
M16 6 4 5 VNW pch L=4e-08 W=2.5e-07 
M17 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M18 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M19 7 6 VDD VNW pch L=4e-08 W=3.35e-07 
M20 8 1 7 VNW pch L=4e-08 W=2.5e-07 
M21 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M24 QN 8 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 8 QN VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFQN_X3M_A9TR QN VDD VNW VPW VSS CK D
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=3.1e-07 
M7 8 4 7 VPW nch L=4e-08 W=3.1e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M11 QN 8 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 8 QN VPW nch L=4e-08 W=3.1e-07 
M13 QN 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M16 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M17 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M18 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M20 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M21 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M22 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M25 QN 8 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 8 QN VNW pch L=4e-08 W=4e-07 
M27 QN 8 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.2e-07 
M7 8 4 7 VPW nch L=4e-08 W=1.2e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M11 Q 9 VSS VPW nch L=4e-08 W=1.55e-07 
M12 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M13 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M14 5 D VDD VNW pch L=4e-08 W=2.5e-07 
M15 6 4 5 VNW pch L=4e-08 W=1.2e-07 
M16 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.55e-07 
M19 8 1 7 VNW pch L=4e-08 W=1.2e-07 
M20 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 8 9 VNW pch L=4e-08 W=1.55e-07 
M23 Q 9 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT DFFQ_X1M_A9TR Q VDD VNW VPW VSS CK D
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.4e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.6e-07 
M7 8 4 7 VPW nch L=4e-08 W=1.6e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 8 9 VPW nch L=4e-08 W=1.75e-07 
M11 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M13 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M14 5 D VDD VNW pch L=4e-08 W=3e-07 
M15 6 4 5 VNW pch L=4e-08 W=1.6e-07 
M16 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M18 7 6 VDD VNW pch L=4e-08 W=2.05e-07 
M19 8 1 7 VNW pch L=4e-08 W=1.6e-07 
M20 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 8 9 VNW pch L=4e-08 W=2.45e-07 
M23 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFQ_X2M_A9TR Q VDD VNW VPW VSS CK D
M0 VSS CK 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.5e-07 
M3 6 1 5 VPW nch L=4e-08 W=2.5e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2.5e-07 
M7 8 4 7 VPW nch L=4e-08 W=2.5e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 8 9 VPW nch L=4e-08 W=2.5e-07 
M11 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M13 VDD CK 1 VNW pch L=4e-08 W=1.4e-07 
M14 4 1 VDD VNW pch L=4e-08 W=2.7e-07 
M15 5 D VDD VNW pch L=4e-08 W=3e-07 
M16 6 4 5 VNW pch L=4e-08 W=2.5e-07 
M17 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M18 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M19 7 6 VDD VNW pch L=4e-08 W=3.25e-07 
M20 8 1 7 VNW pch L=4e-08 W=2.5e-07 
M21 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 8 9 VNW pch L=4e-08 W=3.8e-07 
M24 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFQ_X3M_A9TR Q VDD VNW VPW VSS CK D
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=3.1e-07 
M7 8 4 7 VPW nch L=4e-08 W=3.1e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 8 9 VPW nch L=4e-08 W=2.5e-07 
M11 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M13 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M16 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M17 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M18 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M20 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M21 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M22 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 8 9 VNW pch L=4e-08 W=3.8e-07 
M25 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M26 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M27 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFQ_X4M_A9TR Q VDD VNW VPW VSS CK D
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 15 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=3.1e-07 
M7 8 4 7 VPW nch L=4e-08 W=3.1e-07 
M8 16 1 8 VPW nch L=4e-08 W=1.2e-07 
M9 VSS 9 16 VPW nch L=4e-08 W=1.2e-07 
M10 9 8 VSS VPW nch L=4e-08 W=2.5e-07 
M11 VSS 8 9 VPW nch L=4e-08 W=2.5e-07 
M12 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M14 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M16 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M17 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M18 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M19 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M20 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M22 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M23 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M24 14 4 8 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 9 14 VNW pch L=4e-08 W=1.2e-07 
M26 9 8 VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD 8 9 VNW pch L=4e-08 W=3.8e-07 
M28 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M29 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M30 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFRPQN_X0P5M_A9TR QN VDD VNW VPW VSS CK D R
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 18 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 18 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.2e-07 
M7 VSS R 7 VPW nch L=4e-08 W=1.2e-07 
M8 8 4 7 VPW nch L=4e-08 W=1.2e-07 
M9 19 1 8 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 9 19 VPW nch L=4e-08 W=1.2e-07 
M11 8 R VSS VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 QN 8 VSS VPW nch L=4e-08 W=1.65e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M16 5 D VDD VNW pch L=4e-08 W=2.7e-07 
M17 6 4 5 VNW pch L=4e-08 W=1.2e-07 
M18 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M20 15 6 VDD VNW pch L=4e-08 W=2.7e-07 
M21 7 R 15 VNW pch L=4e-08 W=2.7e-07 
M22 8 1 7 VNW pch L=4e-08 W=1.2e-07 
M23 16 4 8 VNW pch L=4e-08 W=1.6e-07 
M24 17 9 16 VNW pch L=4e-08 W=1.6e-07 
M25 VDD R 17 VNW pch L=4e-08 W=1.6e-07 
M26 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M27 QN 8 VDD VNW pch L=4e-08 W=1.8e-07 
.ENDS


.SUBCKT DFFRPQN_X1M_A9TR QN VDD VNW VPW VSS CK D R
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.4e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.5e-07 
M4 18 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 18 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.5e-07 
M7 VSS R 7 VPW nch L=4e-08 W=1.5e-07 
M8 8 4 7 VPW nch L=4e-08 W=1.5e-07 
M9 19 1 8 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 9 19 VPW nch L=4e-08 W=1.2e-07 
M11 8 R VSS VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 QN 8 VSS VPW nch L=4e-08 W=3.3e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M16 5 D VDD VNW pch L=4e-08 W=3.3e-07 
M17 6 4 5 VNW pch L=4e-08 W=1.7e-07 
M18 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M20 15 6 VDD VNW pch L=4e-08 W=3.3e-07 
M21 7 R 15 VNW pch L=4e-08 W=3.3e-07 
M22 8 1 7 VNW pch L=4e-08 W=1.7e-07 
M23 16 4 8 VNW pch L=4e-08 W=1.6e-07 
M24 17 9 16 VNW pch L=4e-08 W=1.6e-07 
M25 VDD R 17 VNW pch L=4e-08 W=1.6e-07 
M26 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M27 QN 8 VDD VNW pch L=4e-08 W=3.6e-07 
.ENDS


.SUBCKT DFFRPQN_X2M_A9TR QN VDD VNW VPW VSS CK D R
M0 VSS CK 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=2e-07 
M4 18 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 18 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2e-07 
M7 VSS R 7 VPW nch L=4e-08 W=2e-07 
M8 8 4 7 VPW nch L=4e-08 W=2e-07 
M9 19 1 8 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 9 19 VPW nch L=4e-08 W=1.2e-07 
M11 8 R VSS VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 QN 8 VSS VPW nch L=4e-08 W=3.3e-07 
M14 VSS 8 QN VPW nch L=4e-08 W=3.3e-07 
M15 VDD CK 1 VNW pch L=4e-08 W=1.4e-07 
M16 4 1 VDD VNW pch L=4e-08 W=2.7e-07 
M17 5 D VDD VNW pch L=4e-08 W=3.2e-07 
M18 6 4 5 VNW pch L=4e-08 W=3e-07 
M19 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M20 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M21 15 6 VDD VNW pch L=4e-08 W=3.8e-07 
M22 7 R 15 VNW pch L=4e-08 W=3.8e-07 
M23 8 1 7 VNW pch L=4e-08 W=3e-07 
M24 16 4 8 VNW pch L=4e-08 W=1.6e-07 
M25 17 9 16 VNW pch L=4e-08 W=1.6e-07 
M26 VDD R 17 VNW pch L=4e-08 W=1.6e-07 
M27 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M28 QN 8 VDD VNW pch L=4e-08 W=3.6e-07 
M29 VDD 8 QN VNW pch L=4e-08 W=3.6e-07 
.ENDS


.SUBCKT DFFRPQN_X3M_A9TR QN VDD VNW VPW VSS CK D R
M0 VSS CK 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.3e-07 
M3 6 1 5 VPW nch L=4e-08 W=2e-07 
M4 18 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 18 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2e-07 
M7 VSS R 7 VPW nch L=4e-08 W=2e-07 
M8 8 4 7 VPW nch L=4e-08 W=2e-07 
M9 19 1 8 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 9 19 VPW nch L=4e-08 W=1.2e-07 
M11 8 R VSS VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 QN 8 VSS VPW nch L=4e-08 W=3.4e-07 
M14 VSS 8 QN VPW nch L=4e-08 W=3.4e-07 
M15 QN 8 VSS VPW nch L=4e-08 W=3.4e-07 
M16 VDD CK 1 VNW pch L=4e-08 W=1.4e-07 
M17 4 1 VDD VNW pch L=4e-08 W=2.7e-07 
M18 5 D VDD VNW pch L=4e-08 W=3.6e-07 
M19 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M20 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M22 15 6 VDD VNW pch L=4e-08 W=3.8e-07 
M23 7 R 15 VNW pch L=4e-08 W=3.8e-07 
M24 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M25 16 4 8 VNW pch L=4e-08 W=1.6e-07 
M26 17 9 16 VNW pch L=4e-08 W=1.6e-07 
M27 VDD R 17 VNW pch L=4e-08 W=1.6e-07 
M28 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M29 QN 8 VDD VNW pch L=4e-08 W=3.5e-07 
M30 VDD 8 QN VNW pch L=4e-08 W=3.5e-07 
M31 QN 8 VDD VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT DFFRPQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D R
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 18 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 18 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.2e-07 
M7 VSS R 7 VPW nch L=4e-08 W=1.2e-07 
M8 8 4 7 VPW nch L=4e-08 W=1.2e-07 
M9 19 1 8 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 9 19 VPW nch L=4e-08 W=1.2e-07 
M11 8 R VSS VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 Q 9 VSS VPW nch L=4e-08 W=1.55e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M16 5 D VDD VNW pch L=4e-08 W=2.5e-07 
M17 6 4 5 VNW pch L=4e-08 W=1.2e-07 
M18 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M20 15 6 VDD VNW pch L=4e-08 W=2.5e-07 
M21 7 R 15 VNW pch L=4e-08 W=2.5e-07 
M22 8 1 7 VNW pch L=4e-08 W=1.2e-07 
M23 16 4 8 VNW pch L=4e-08 W=1.6e-07 
M24 17 9 16 VNW pch L=4e-08 W=1.6e-07 
M25 VDD R 17 VNW pch L=4e-08 W=1.6e-07 
M26 VDD 8 9 VNW pch L=4e-08 W=1.35e-07 
M27 Q 9 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT DFFRPQ_X1M_A9TR Q VDD VNW VPW VSS CK D R
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.4e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 18 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 18 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS R 7 VPW nch L=4e-08 W=1.6e-07 
M8 8 4 7 VPW nch L=4e-08 W=1.6e-07 
M9 19 1 8 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 9 19 VPW nch L=4e-08 W=1.2e-07 
M11 8 R VSS VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.95e-07 
M13 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M16 5 D VDD VNW pch L=4e-08 W=3.1e-07 
M17 6 4 5 VNW pch L=4e-08 W=1.6e-07 
M18 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M20 15 6 VDD VNW pch L=4e-08 W=3.2e-07 
M21 7 R 15 VNW pch L=4e-08 W=3.2e-07 
M22 8 1 7 VNW pch L=4e-08 W=1.6e-07 
M23 16 4 8 VNW pch L=4e-08 W=1.6e-07 
M24 17 9 16 VNW pch L=4e-08 W=1.6e-07 
M25 VDD R 17 VNW pch L=4e-08 W=1.6e-07 
M26 VDD 8 9 VNW pch L=4e-08 W=2.25e-07 
M27 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFRPQ_X2M_A9TR Q VDD VNW VPW VSS CK D R
M0 VSS CK 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=2.5e-07 
M4 18 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 18 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2.5e-07 
M7 VSS R 7 VPW nch L=4e-08 W=2.5e-07 
M8 8 4 7 VPW nch L=4e-08 W=2.5e-07 
M9 19 1 8 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 9 19 VPW nch L=4e-08 W=1.2e-07 
M11 8 R VSS VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=3e-07 
M13 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M15 VDD CK 1 VNW pch L=4e-08 W=1.4e-07 
M16 4 1 VDD VNW pch L=4e-08 W=2.7e-07 
M17 5 D VDD VNW pch L=4e-08 W=3.2e-07 
M18 6 4 5 VNW pch L=4e-08 W=2.5e-07 
M19 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M20 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M21 15 6 VDD VNW pch L=4e-08 W=3.8e-07 
M22 7 R 15 VNW pch L=4e-08 W=3.8e-07 
M23 8 1 7 VNW pch L=4e-08 W=2.5e-07 
M24 16 4 8 VNW pch L=4e-08 W=1.6e-07 
M25 17 9 16 VNW pch L=4e-08 W=1.6e-07 
M26 VDD R 17 VNW pch L=4e-08 W=1.6e-07 
M27 VDD 8 9 VNW pch L=4e-08 W=3.4e-07 
M28 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M29 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFRPQ_X3M_A9TR Q VDD VNW VPW VSS CK D R
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.3e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 18 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 18 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2.5e-07 
M7 VSS R 7 VPW nch L=4e-08 W=2.5e-07 
M8 8 4 7 VPW nch L=4e-08 W=3.1e-07 
M9 19 1 8 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 9 19 VPW nch L=4e-08 W=1.2e-07 
M11 8 R VSS VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=3.4e-07 
M13 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M15 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M17 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M18 5 D VDD VNW pch L=4e-08 W=3.6e-07 
M19 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M20 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M22 15 6 VDD VNW pch L=4e-08 W=3.8e-07 
M23 7 R 15 VNW pch L=4e-08 W=3.8e-07 
M24 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M25 16 4 8 VNW pch L=4e-08 W=1.6e-07 
M26 17 9 16 VNW pch L=4e-08 W=1.6e-07 
M27 VDD R 17 VNW pch L=4e-08 W=1.6e-07 
M28 VDD 8 9 VNW pch L=4e-08 W=3.8e-07 
M29 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M31 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFRPQ_X4M_A9TR Q VDD VNW VPW VSS CK D R
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.3e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 18 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 18 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2.5e-07 
M7 VSS R 7 VPW nch L=4e-08 W=2.5e-07 
M8 8 4 7 VPW nch L=4e-08 W=3.1e-07 
M9 19 1 8 VPW nch L=4e-08 W=1.2e-07 
M10 VSS 9 19 VPW nch L=4e-08 W=1.2e-07 
M11 8 R VSS VPW nch L=4e-08 W=1.2e-07 
M12 9 8 VSS VPW nch L=4e-08 W=3e-07 
M13 VSS 8 9 VPW nch L=4e-08 W=3e-07 
M14 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M16 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M18 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M19 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M20 5 D VDD VNW pch L=4e-08 W=3.6e-07 
M21 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M22 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M24 15 6 VDD VNW pch L=4e-08 W=3.8e-07 
M25 7 R 15 VNW pch L=4e-08 W=3.8e-07 
M26 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M27 16 4 8 VNW pch L=4e-08 W=1.6e-07 
M28 17 9 16 VNW pch L=4e-08 W=1.6e-07 
M29 VDD R 17 VNW pch L=4e-08 W=1.6e-07 
M30 9 8 VDD VNW pch L=4e-08 W=3.2e-07 
M31 VDD 8 9 VNW pch L=4e-08 W=3.2e-07 
M32 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M34 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFSQN_X0P5M_A9TR QN VDD VNW VPW VSS CK D SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 16 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 16 VPW nch L=4e-08 W=1.2e-07 
M6 17 6 VSS VPW nch L=4e-08 W=1.8e-07 
M7 7 SN 17 VPW nch L=4e-08 W=1.8e-07 
M8 8 4 7 VPW nch L=4e-08 W=1.2e-07 
M9 18 1 8 VPW nch L=4e-08 W=1.6e-07 
M10 19 9 18 VPW nch L=4e-08 W=1.6e-07 
M11 VSS SN 19 VPW nch L=4e-08 W=1.6e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 QN 8 VSS VPW nch L=4e-08 W=1.55e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M16 5 D VDD VNW pch L=4e-08 W=2.6e-07 
M17 6 4 5 VNW pch L=4e-08 W=1.2e-07 
M18 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M20 7 6 VDD VNW pch L=4e-08 W=1.55e-07 
M21 VDD SN 7 VNW pch L=4e-08 W=1.55e-07 
M22 8 1 7 VNW pch L=4e-08 W=1.2e-07 
M23 15 4 8 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 9 15 VNW pch L=4e-08 W=1.2e-07 
M25 8 SN VDD VNW pch L=4e-08 W=1.2e-07 
M26 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M27 QN 8 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT DFFSQN_X1M_A9TR QN VDD VNW VPW VSS CK D SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.4e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 16 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 16 VPW nch L=4e-08 W=1.2e-07 
M6 17 6 VSS VPW nch L=4e-08 W=2.45e-07 
M7 7 SN 17 VPW nch L=4e-08 W=2.45e-07 
M8 8 4 7 VPW nch L=4e-08 W=1.6e-07 
M9 18 1 8 VPW nch L=4e-08 W=1.6e-07 
M10 19 9 18 VPW nch L=4e-08 W=1.6e-07 
M11 VSS SN 19 VPW nch L=4e-08 W=1.6e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 QN 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M16 5 D VDD VNW pch L=4e-08 W=3.2e-07 
M17 6 4 5 VNW pch L=4e-08 W=1.6e-07 
M18 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M20 7 6 VDD VNW pch L=4e-08 W=2.05e-07 
M21 VDD SN 7 VNW pch L=4e-08 W=2.05e-07 
M22 8 1 7 VNW pch L=4e-08 W=1.6e-07 
M23 15 4 8 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 9 15 VNW pch L=4e-08 W=1.2e-07 
M25 8 SN VDD VNW pch L=4e-08 W=1.2e-07 
M26 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M27 QN 8 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFSQN_X2M_A9TR QN VDD VNW VPW VSS CK D SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=2.5e-07 
M4 16 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 16 VPW nch L=4e-08 W=1.2e-07 
M6 17 6 VSS VPW nch L=4e-08 W=3.8e-07 
M7 7 SN 17 VPW nch L=4e-08 W=3.8e-07 
M8 8 4 7 VPW nch L=4e-08 W=2.5e-07 
M9 18 1 8 VPW nch L=4e-08 W=1.6e-07 
M10 19 9 18 VPW nch L=4e-08 W=1.6e-07 
M11 VSS SN 19 VPW nch L=4e-08 W=1.6e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 QN 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 8 QN VPW nch L=4e-08 W=3.1e-07 
M15 VDD CK 1 VNW pch L=4e-08 W=1.4e-07 
M16 4 1 VDD VNW pch L=4e-08 W=2.7e-07 
M17 5 D VDD VNW pch L=4e-08 W=3.2e-07 
M18 6 4 5 VNW pch L=4e-08 W=2.5e-07 
M19 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M20 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M21 7 6 VDD VNW pch L=4e-08 W=3.2e-07 
M22 VDD SN 7 VNW pch L=4e-08 W=3.2e-07 
M23 8 1 7 VNW pch L=4e-08 W=2.5e-07 
M24 15 4 8 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 9 15 VNW pch L=4e-08 W=1.2e-07 
M26 8 SN VDD VNW pch L=4e-08 W=1.2e-07 
M27 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M28 QN 8 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 8 QN VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFSQN_X3M_A9TR QN VDD VNW VPW VSS CK D SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 16 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 16 VPW nch L=4e-08 W=1.2e-07 
M6 17 6 VSS VPW nch L=4e-08 W=3.8e-07 
M7 7 SN 17 VPW nch L=4e-08 W=3.8e-07 
M8 8 4 7 VPW nch L=4e-08 W=3.1e-07 
M9 18 1 8 VPW nch L=4e-08 W=1.6e-07 
M10 19 9 18 VPW nch L=4e-08 W=1.6e-07 
M11 VSS SN 19 VPW nch L=4e-08 W=1.6e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 QN 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 8 QN VPW nch L=4e-08 W=3.1e-07 
M15 QN 8 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M17 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M18 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M19 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M20 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M22 7 6 VDD VNW pch L=4e-08 W=3.2e-07 
M23 VDD SN 7 VNW pch L=4e-08 W=3.2e-07 
M24 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M25 15 4 8 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 9 15 VNW pch L=4e-08 W=1.2e-07 
M27 8 SN VDD VNW pch L=4e-08 W=1.2e-07 
M28 VDD 8 9 VNW pch L=4e-08 W=1.2e-07 
M29 QN 8 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 8 QN VNW pch L=4e-08 W=4e-07 
M31 QN 8 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFSQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 16 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 16 VPW nch L=4e-08 W=1.2e-07 
M6 17 SN VSS VPW nch L=4e-08 W=1.8e-07 
M7 7 6 17 VPW nch L=4e-08 W=1.8e-07 
M8 8 4 7 VPW nch L=4e-08 W=1.2e-07 
M9 18 1 8 VPW nch L=4e-08 W=1.6e-07 
M10 19 9 18 VPW nch L=4e-08 W=1.6e-07 
M11 VSS SN 19 VPW nch L=4e-08 W=1.6e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M13 Q 9 VSS VPW nch L=4e-08 W=1.55e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M16 5 D VDD VNW pch L=4e-08 W=2.6e-07 
M17 6 4 5 VNW pch L=4e-08 W=1.2e-07 
M18 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M20 7 SN VDD VNW pch L=4e-08 W=1.55e-07 
M21 VDD 6 7 VNW pch L=4e-08 W=1.55e-07 
M22 8 1 7 VNW pch L=4e-08 W=1.2e-07 
M23 15 4 8 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 9 15 VNW pch L=4e-08 W=1.2e-07 
M25 8 SN VDD VNW pch L=4e-08 W=1.2e-07 
M26 VDD 8 9 VNW pch L=4e-08 W=1.6e-07 
M27 Q 9 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT DFFSQ_X1M_A9TR Q VDD VNW VPW VSS CK D SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.4e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 16 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 16 VPW nch L=4e-08 W=1.2e-07 
M6 17 SN VSS VPW nch L=4e-08 W=2.4e-07 
M7 7 6 17 VPW nch L=4e-08 W=2.4e-07 
M8 8 4 7 VPW nch L=4e-08 W=1.6e-07 
M9 18 1 8 VPW nch L=4e-08 W=1.6e-07 
M10 19 9 18 VPW nch L=4e-08 W=1.6e-07 
M11 VSS SN 19 VPW nch L=4e-08 W=1.6e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=1.65e-07 
M13 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M15 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M16 5 D VDD VNW pch L=4e-08 W=3.2e-07 
M17 6 4 5 VNW pch L=4e-08 W=1.6e-07 
M18 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M20 7 SN VDD VNW pch L=4e-08 W=2.05e-07 
M21 VDD 6 7 VNW pch L=4e-08 W=2.05e-07 
M22 8 1 7 VNW pch L=4e-08 W=1.6e-07 
M23 15 4 8 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 9 15 VNW pch L=4e-08 W=1.2e-07 
M25 8 SN VDD VNW pch L=4e-08 W=1.2e-07 
M26 VDD 8 9 VNW pch L=4e-08 W=2.55e-07 
M27 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFSQ_X2M_A9TR Q VDD VNW VPW VSS CK D SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=2.5e-07 
M4 16 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 16 VPW nch L=4e-08 W=1.2e-07 
M6 17 SN VSS VPW nch L=4e-08 W=3.8e-07 
M7 7 6 17 VPW nch L=4e-08 W=3.8e-07 
M8 8 4 7 VPW nch L=4e-08 W=2.5e-07 
M9 18 1 8 VPW nch L=4e-08 W=1.6e-07 
M10 19 9 18 VPW nch L=4e-08 W=1.6e-07 
M11 VSS SN 19 VPW nch L=4e-08 W=1.6e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=2.5e-07 
M13 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M15 VDD CK 1 VNW pch L=4e-08 W=1.4e-07 
M16 4 1 VDD VNW pch L=4e-08 W=2.7e-07 
M17 5 D VDD VNW pch L=4e-08 W=3.2e-07 
M18 6 4 5 VNW pch L=4e-08 W=2.5e-07 
M19 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M20 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M21 7 SN VDD VNW pch L=4e-08 W=3.25e-07 
M22 VDD 6 7 VNW pch L=4e-08 W=3.25e-07 
M23 8 1 7 VNW pch L=4e-08 W=2.5e-07 
M24 15 4 8 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 9 15 VNW pch L=4e-08 W=1.2e-07 
M26 8 SN VDD VNW pch L=4e-08 W=1.2e-07 
M27 VDD 8 9 VNW pch L=4e-08 W=3.8e-07 
M28 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M29 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFSQ_X3M_A9TR Q VDD VNW VPW VSS CK D SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 16 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 16 VPW nch L=4e-08 W=1.2e-07 
M6 17 SN VSS VPW nch L=4e-08 W=3.8e-07 
M7 7 6 17 VPW nch L=4e-08 W=3.8e-07 
M8 8 4 7 VPW nch L=4e-08 W=3.1e-07 
M9 18 1 8 VPW nch L=4e-08 W=1.6e-07 
M10 19 9 18 VPW nch L=4e-08 W=1.6e-07 
M11 VSS SN 19 VPW nch L=4e-08 W=1.6e-07 
M12 VSS 8 9 VPW nch L=4e-08 W=2.5e-07 
M13 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M15 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M17 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M18 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M19 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M20 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M22 7 SN VDD VNW pch L=4e-08 W=3.25e-07 
M23 VDD 6 7 VNW pch L=4e-08 W=3.25e-07 
M24 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M25 15 4 8 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 9 15 VNW pch L=4e-08 W=1.2e-07 
M27 8 SN VDD VNW pch L=4e-08 W=1.2e-07 
M28 VDD 8 9 VNW pch L=4e-08 W=3.8e-07 
M29 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M31 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFSQ_X4M_A9TR Q VDD VNW VPW VSS CK D SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 16 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 16 VPW nch L=4e-08 W=1.2e-07 
M6 17 SN VSS VPW nch L=4e-08 W=3.8e-07 
M7 7 6 17 VPW nch L=4e-08 W=3.8e-07 
M8 8 4 7 VPW nch L=4e-08 W=3.1e-07 
M9 18 1 8 VPW nch L=4e-08 W=1.6e-07 
M10 19 9 18 VPW nch L=4e-08 W=1.6e-07 
M11 VSS SN 19 VPW nch L=4e-08 W=1.6e-07 
M12 9 8 VSS VPW nch L=4e-08 W=1.9e-07 
M13 VSS 8 9 VPW nch L=4e-08 W=1.9e-07 
M14 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M16 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M18 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M19 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M20 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M21 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M22 14 1 6 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 7 14 VNW pch L=4e-08 W=1.2e-07 
M24 7 SN VDD VNW pch L=4e-08 W=3.25e-07 
M25 VDD 6 7 VNW pch L=4e-08 W=3.25e-07 
M26 8 1 7 VNW pch L=4e-08 W=3.1e-07 
M27 15 4 8 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 9 15 VNW pch L=4e-08 W=1.2e-07 
M29 8 SN VDD VNW pch L=4e-08 W=1.2e-07 
M30 9 8 VDD VNW pch L=4e-08 W=3.4e-07 
M31 VDD 8 9 VNW pch L=4e-08 W=3.4e-07 
M32 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M34 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT DFFSRPQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D R SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=1.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 21 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 8 21 VPW nch L=4e-08 W=1.2e-07 
M6 7 SN VSS VPW nch L=4e-08 W=1.8e-07 
M7 8 6 7 VPW nch L=4e-08 W=1.8e-07 
M8 7 R 8 VPW nch L=4e-08 W=1.8e-07 
M9 9 4 8 VPW nch L=4e-08 W=1.2e-07 
M10 22 1 9 VPW nch L=4e-08 W=1.6e-07 
M11 23 10 22 VPW nch L=4e-08 W=1.6e-07 
M12 VSS SN 23 VPW nch L=4e-08 W=1.6e-07 
M13 24 R VSS VPW nch L=4e-08 W=1.6e-07 
M14 9 SN 24 VPW nch L=4e-08 W=1.6e-07 
M15 VSS 9 10 VPW nch L=4e-08 W=1.2e-07 
M16 Q 10 VSS VPW nch L=4e-08 W=1.55e-07 
M17 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M18 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M19 5 D VDD VNW pch L=4e-08 W=2.6e-07 
M20 6 4 5 VNW pch L=4e-08 W=1.2e-07 
M21 16 1 6 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 8 16 VNW pch L=4e-08 W=1.2e-07 
M23 8 SN VDD VNW pch L=4e-08 W=2.6e-07 
M24 17 6 8 VNW pch L=4e-08 W=2.6e-07 
M25 VDD R 17 VNW pch L=4e-08 W=2.6e-07 
M26 9 1 8 VNW pch L=4e-08 W=1.2e-07 
M27 18 4 9 VNW pch L=4e-08 W=1.6e-07 
M28 19 10 18 VNW pch L=4e-08 W=1.6e-07 
M29 VDD R 19 VNW pch L=4e-08 W=1.6e-07 
M30 9 SN VDD VNW pch L=4e-08 W=1.6e-07 
M31 VDD 9 10 VNW pch L=4e-08 W=1.3e-07 
M32 Q 10 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT DFFSRPQ_X1M_A9TR Q VDD VNW VPW VSS CK D R SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.4e-07 
M3 6 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 21 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 8 21 VPW nch L=4e-08 W=1.2e-07 
M6 7 SN VSS VPW nch L=4e-08 W=2.4e-07 
M7 8 6 7 VPW nch L=4e-08 W=2.4e-07 
M8 7 R 8 VPW nch L=4e-08 W=2.4e-07 
M9 9 4 8 VPW nch L=4e-08 W=1.6e-07 
M10 22 1 9 VPW nch L=4e-08 W=1.6e-07 
M11 23 10 22 VPW nch L=4e-08 W=1.6e-07 
M12 VSS SN 23 VPW nch L=4e-08 W=1.6e-07 
M13 24 R VSS VPW nch L=4e-08 W=1.6e-07 
M14 9 SN 24 VPW nch L=4e-08 W=1.6e-07 
M15 VSS 9 10 VPW nch L=4e-08 W=2e-07 
M16 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VDD CK 1 VNW pch L=4e-08 W=1.3e-07 
M18 4 1 VDD VNW pch L=4e-08 W=2.5e-07 
M19 5 D VDD VNW pch L=4e-08 W=3.1e-07 
M20 6 4 5 VNW pch L=4e-08 W=1.6e-07 
M21 16 1 6 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 8 16 VNW pch L=4e-08 W=1.2e-07 
M23 8 SN VDD VNW pch L=4e-08 W=3.2e-07 
M24 17 6 8 VNW pch L=4e-08 W=3.2e-07 
M25 VDD R 17 VNW pch L=4e-08 W=3.2e-07 
M26 9 1 8 VNW pch L=4e-08 W=1.6e-07 
M27 18 4 9 VNW pch L=4e-08 W=1.6e-07 
M28 19 10 18 VNW pch L=4e-08 W=1.6e-07 
M29 VDD R 19 VNW pch L=4e-08 W=1.6e-07 
M30 9 SN VDD VNW pch L=4e-08 W=1.6e-07 
M31 VDD 9 10 VNW pch L=4e-08 W=2.2e-07 
M32 Q 10 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFSRPQ_X2M_A9TR Q VDD VNW VPW VSS CK D R SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.3e-07 
M2 5 D VSS VPW nch L=4e-08 W=2.8e-07 
M3 6 1 5 VPW nch L=4e-08 W=2.5e-07 
M4 21 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 8 21 VPW nch L=4e-08 W=1.2e-07 
M6 7 SN VSS VPW nch L=4e-08 W=2.95e-07 
M7 8 6 7 VPW nch L=4e-08 W=2.95e-07 
M8 7 R 8 VPW nch L=4e-08 W=2.95e-07 
M9 9 4 8 VPW nch L=4e-08 W=2.5e-07 
M10 22 1 9 VPW nch L=4e-08 W=1.6e-07 
M11 23 10 22 VPW nch L=4e-08 W=1.6e-07 
M12 VSS SN 23 VPW nch L=4e-08 W=1.6e-07 
M13 24 R VSS VPW nch L=4e-08 W=1.6e-07 
M14 9 SN 24 VPW nch L=4e-08 W=1.6e-07 
M15 VSS 9 10 VPW nch L=4e-08 W=3e-07 
M16 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 10 Q VPW nch L=4e-08 W=3.1e-07 
M18 VDD CK 1 VNW pch L=4e-08 W=1.4e-07 
M19 4 1 VDD VNW pch L=4e-08 W=2.7e-07 
M20 5 D VDD VNW pch L=4e-08 W=3.2e-07 
M21 6 4 5 VNW pch L=4e-08 W=2.5e-07 
M22 16 1 6 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 8 16 VNW pch L=4e-08 W=1.2e-07 
M24 8 SN VDD VNW pch L=4e-08 W=3.8e-07 
M25 17 6 8 VNW pch L=4e-08 W=3.8e-07 
M26 VDD R 17 VNW pch L=4e-08 W=3.8e-07 
M27 9 1 8 VNW pch L=4e-08 W=2.5e-07 
M28 18 4 9 VNW pch L=4e-08 W=1.6e-07 
M29 19 10 18 VNW pch L=4e-08 W=1.6e-07 
M30 VDD R 19 VNW pch L=4e-08 W=1.6e-07 
M31 9 SN VDD VNW pch L=4e-08 W=1.6e-07 
M32 VDD 9 10 VNW pch L=4e-08 W=3.35e-07 
M33 Q 10 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 10 Q VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFSRPQ_X3M_A9TR Q VDD VNW VPW VSS CK D R SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 21 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 8 21 VPW nch L=4e-08 W=1.2e-07 
M6 7 SN VSS VPW nch L=4e-08 W=2.95e-07 
M7 8 6 7 VPW nch L=4e-08 W=2.95e-07 
M8 7 R 8 VPW nch L=4e-08 W=2.95e-07 
M9 9 4 8 VPW nch L=4e-08 W=3.1e-07 
M10 22 1 9 VPW nch L=4e-08 W=1.6e-07 
M11 23 10 22 VPW nch L=4e-08 W=1.6e-07 
M12 VSS SN 23 VPW nch L=4e-08 W=1.6e-07 
M13 24 R VSS VPW nch L=4e-08 W=1.6e-07 
M14 9 SN 24 VPW nch L=4e-08 W=1.6e-07 
M15 VSS 9 10 VPW nch L=4e-08 W=3.1e-07 
M16 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 10 Q VPW nch L=4e-08 W=3.1e-07 
M18 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M20 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M21 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M22 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M23 16 1 6 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 8 16 VNW pch L=4e-08 W=1.2e-07 
M25 8 SN VDD VNW pch L=4e-08 W=3.8e-07 
M26 17 6 8 VNW pch L=4e-08 W=3.8e-07 
M27 VDD R 17 VNW pch L=4e-08 W=3.8e-07 
M28 9 1 8 VNW pch L=4e-08 W=3.1e-07 
M29 18 4 9 VNW pch L=4e-08 W=1.6e-07 
M30 19 10 18 VNW pch L=4e-08 W=1.6e-07 
M31 VDD R 19 VNW pch L=4e-08 W=1.6e-07 
M32 9 SN VDD VNW pch L=4e-08 W=1.6e-07 
M33 VDD 9 10 VNW pch L=4e-08 W=3.8e-07 
M34 Q 10 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 10 Q VNW pch L=4e-08 W=4e-07 
M36 Q 10 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DFFSRPQ_X4M_A9TR Q VDD VNW VPW VSS CK D R SN
M0 VSS CK 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 1 VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 D VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 1 5 VPW nch L=4e-08 W=3.1e-07 
M4 21 4 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 8 21 VPW nch L=4e-08 W=1.2e-07 
M6 7 SN VSS VPW nch L=4e-08 W=2.95e-07 
M7 8 6 7 VPW nch L=4e-08 W=2.95e-07 
M8 7 R 8 VPW nch L=4e-08 W=2.95e-07 
M9 9 4 8 VPW nch L=4e-08 W=3.1e-07 
M10 22 1 9 VPW nch L=4e-08 W=1.6e-07 
M11 23 10 22 VPW nch L=4e-08 W=1.6e-07 
M12 VSS SN 23 VPW nch L=4e-08 W=1.6e-07 
M13 24 R VSS VPW nch L=4e-08 W=1.6e-07 
M14 9 SN 24 VPW nch L=4e-08 W=1.6e-07 
M15 10 9 VSS VPW nch L=4e-08 W=3e-07 
M16 VSS 9 10 VPW nch L=4e-08 W=3e-07 
M17 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M18 VSS 10 Q VPW nch L=4e-08 W=3.1e-07 
M19 Q 10 VSS VPW nch L=4e-08 W=3.1e-07 
M20 VSS 10 Q VPW nch L=4e-08 W=3.1e-07 
M21 VDD CK 1 VNW pch L=4e-08 W=1.5e-07 
M22 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M23 5 D VDD VNW pch L=4e-08 W=3.8e-07 
M24 6 4 5 VNW pch L=4e-08 W=3.1e-07 
M25 16 1 6 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 8 16 VNW pch L=4e-08 W=1.2e-07 
M27 8 SN VDD VNW pch L=4e-08 W=3.8e-07 
M28 17 6 8 VNW pch L=4e-08 W=3.8e-07 
M29 VDD R 17 VNW pch L=4e-08 W=3.8e-07 
M30 9 1 8 VNW pch L=4e-08 W=3.1e-07 
M31 18 4 9 VNW pch L=4e-08 W=1.6e-07 
M32 19 10 18 VNW pch L=4e-08 W=1.6e-07 
M33 VDD R 19 VNW pch L=4e-08 W=1.6e-07 
M34 9 SN VDD VNW pch L=4e-08 W=1.6e-07 
M35 10 9 VDD VNW pch L=4e-08 W=3.2e-07 
M36 VDD 9 10 VNW pch L=4e-08 W=3.2e-07 
M37 Q 10 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 10 Q VNW pch L=4e-08 W=4e-07 
M39 Q 10 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD 10 Q VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DLY2_X0P5M_A9TR Y VDD VNW VPW VSS A
M0 7 A 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A 7 VPW nch L=4e-08 W=1.2e-07 
M2 VSS 1 VSS VPW nch L=4e-08 W=1.35e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=1.55e-07 
M4 6 A 1 VNW pch L=4e-08 W=1.55e-07 
M5 VDD A 6 VNW pch L=4e-08 W=1.55e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT DLY2_X1M_A9TR Y VDD VNW VPW VSS A
M0 7 A 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A 7 VPW nch L=4e-08 W=1.2e-07 
M2 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 A 1 VNW pch L=4e-08 W=1.55e-07 
M4 VDD A 6 VNW pch L=4e-08 W=1.55e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DLY4_X0P5M_A9TR Y VDD VNW VPW VSS A
M0 11 A 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A 11 VPW nch L=4e-08 W=1.2e-07 
M2 12 1 VSS VPW nch L=4e-08 W=1.2e-07 
M3 4 1 12 VPW nch L=4e-08 W=1.2e-07 
M4 13 4 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 4 13 VPW nch L=4e-08 W=1.2e-07 
M6 VSS 5 VSS VPW nch L=4e-08 W=1.35e-07 
M7 Y 5 VSS VPW nch L=4e-08 W=1.55e-07 
M8 8 A 1 VNW pch L=4e-08 W=1.55e-07 
M9 VDD A 8 VNW pch L=4e-08 W=1.55e-07 
M10 9 1 VDD VNW pch L=4e-08 W=1.55e-07 
M11 4 1 9 VNW pch L=4e-08 W=1.55e-07 
M12 10 4 5 VNW pch L=4e-08 W=1.55e-07 
M13 VDD 4 10 VNW pch L=4e-08 W=1.55e-07 
M14 Y 5 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT DLY4_X1M_A9TR Y VDD VNW VPW VSS A
M0 11 A 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A 11 VPW nch L=4e-08 W=1.2e-07 
M2 12 1 VSS VPW nch L=4e-08 W=1.2e-07 
M3 4 1 12 VPW nch L=4e-08 W=1.2e-07 
M4 13 4 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 4 13 VPW nch L=4e-08 W=1.2e-07 
M6 Y 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 8 A 1 VNW pch L=4e-08 W=1.55e-07 
M8 VDD A 8 VNW pch L=4e-08 W=1.55e-07 
M9 9 1 VDD VNW pch L=4e-08 W=1.55e-07 
M10 4 1 9 VNW pch L=4e-08 W=1.55e-07 
M11 10 4 5 VNW pch L=4e-08 W=1.55e-07 
M12 VDD 4 10 VNW pch L=4e-08 W=1.55e-07 
M13 Y 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DLYCLK8S2_X1B_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.25e-07 
M1 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M2 3 A VDD VNW pch L=4e-08 W=4e-07 
M3 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DLYCLK8S4_X1B_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.25e-07 
M1 4 3 VSS VPW nch L=4e-08 W=2.25e-07 
M2 5 4 VSS VPW nch L=4e-08 W=2.25e-07 
M3 Y 5 VSS VPW nch L=4e-08 W=2.25e-07 
M4 3 A VDD VNW pch L=4e-08 W=4e-07 
M5 4 3 VDD VNW pch L=4e-08 W=4e-07 
M6 5 4 VDD VNW pch L=4e-08 W=4e-07 
M7 Y 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DLYCLK8S6_X1B_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.25e-07 
M1 4 3 VSS VPW nch L=4e-08 W=2.25e-07 
M2 5 4 VSS VPW nch L=4e-08 W=2.25e-07 
M3 6 5 VSS VPW nch L=4e-08 W=2.25e-07 
M4 7 6 VSS VPW nch L=4e-08 W=2.25e-07 
M5 Y 7 VSS VPW nch L=4e-08 W=2.25e-07 
M6 3 A VDD VNW pch L=4e-08 W=4e-07 
M7 4 3 VDD VNW pch L=4e-08 W=4e-07 
M8 5 4 VDD VNW pch L=4e-08 W=4e-07 
M9 6 5 VDD VNW pch L=4e-08 W=4e-07 
M10 7 6 VDD VNW pch L=4e-08 W=4e-07 
M11 Y 7 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT DLYCLK8S8_X1B_A9TR Y VDD VNW VPW VSS A
M0 3 A VSS VPW nch L=4e-08 W=2.25e-07 
M1 4 3 VSS VPW nch L=4e-08 W=2.25e-07 
M2 5 4 VSS VPW nch L=4e-08 W=2.25e-07 
M3 6 5 VSS VPW nch L=4e-08 W=2.25e-07 
M4 7 6 VSS VPW nch L=4e-08 W=2.25e-07 
M5 8 7 VSS VPW nch L=4e-08 W=2.25e-07 
M6 9 8 VSS VPW nch L=4e-08 W=2.25e-07 
M7 Y 9 VSS VPW nch L=4e-08 W=2.25e-07 
M8 3 A VDD VNW pch L=4e-08 W=4e-07 
M9 4 3 VDD VNW pch L=4e-08 W=4e-07 
M10 5 4 VDD VNW pch L=4e-08 W=4e-07 
M11 6 5 VDD VNW pch L=4e-08 W=4e-07 
M12 7 6 VDD VNW pch L=4e-08 W=4e-07 
M13 8 7 VDD VNW pch L=4e-08 W=4e-07 
M14 9 8 VDD VNW pch L=4e-08 W=4e-07 
M15 Y 9 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT ENDCAPTIE3_A9TR VDD VNW VPW VSS
*.CONNECT VNW VDD
*.CONNECT VPW VSS
.ENDS


.SUBCKT ESDFFQN_X0P5M_A9TR QN VDD VNW VPW VSS CK D E SE SI
M0 VSS D 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.2e-07 
M2 6 E 1 VPW nch L=4e-08 W=1.2e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 13 5 VPW nch L=4e-08 W=1.2e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.2e-07 
M7 25 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 25 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=1.2e-07 
M10 10 16 9 VPW nch L=4e-08 W=1.2e-07 
M11 26 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 26 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=1.2e-07 
M14 12 15 11 VPW nch L=4e-08 W=1.2e-07 
M15 27 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 27 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 QN 13 VSS VPW nch L=4e-08 W=1.55e-07 
M19 VSS 16 15 VPW nch L=4e-08 W=1.2e-07 
M20 16 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 VDD D 1 VNW pch L=4e-08 W=2.4e-07 
M22 4 E VDD VNW pch L=4e-08 W=2.2e-07 
M23 6 E 5 VNW pch L=4e-08 W=2.2e-07 
M24 1 4 6 VNW pch L=4e-08 W=2.2e-07 
M25 VDD 13 5 VNW pch L=4e-08 W=2.2e-07 
M26 7 SE VDD VNW pch L=4e-08 W=1.8e-07 
M27 8 SE 6 VNW pch L=4e-08 W=2.2e-07 
M28 22 7 8 VNW pch L=4e-08 W=1.55e-07 
M29 VDD SI 22 VNW pch L=4e-08 W=1.55e-07 
M30 9 8 VDD VNW pch L=4e-08 W=1.3e-07 
M31 10 15 9 VNW pch L=4e-08 W=1.2e-07 
M32 23 16 10 VNW pch L=4e-08 W=1.2e-07 
M33 VDD 11 23 VNW pch L=4e-08 W=1.2e-07 
M34 11 10 VDD VNW pch L=4e-08 W=1.55e-07 
M35 12 16 11 VNW pch L=4e-08 W=1.2e-07 
M36 24 15 12 VNW pch L=4e-08 W=1.2e-07 
M37 VDD 13 24 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 12 13 VNW pch L=4e-08 W=1.55e-07 
M39 QN 13 VDD VNW pch L=4e-08 W=2e-07 
M40 VDD 16 15 VNW pch L=4e-08 W=2.5e-07 
M41 16 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT ESDFFQN_X1M_A9TR QN VDD VNW VPW VSS CK D E SE SI
M0 VSS D 1 VPW nch L=4e-08 W=1.6e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.6e-07 
M2 6 E 1 VPW nch L=4e-08 W=1.6e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.6e-07 
M4 VSS 13 5 VPW nch L=4e-08 W=1.6e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.6e-07 
M7 25 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 25 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=1.6e-07 
M10 10 16 9 VPW nch L=4e-08 W=1.6e-07 
M11 26 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 26 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=1.6e-07 
M14 12 15 11 VPW nch L=4e-08 W=1.6e-07 
M15 27 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 27 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.75e-07 
M18 QN 13 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 16 15 VPW nch L=4e-08 W=1.2e-07 
M20 16 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 VDD D 1 VNW pch L=4e-08 W=3.4e-07 
M22 4 E VDD VNW pch L=4e-08 W=3.2e-07 
M23 6 E 5 VNW pch L=4e-08 W=3.2e-07 
M24 1 4 6 VNW pch L=4e-08 W=3.2e-07 
M25 VDD 13 5 VNW pch L=4e-08 W=3.2e-07 
M26 7 SE VDD VNW pch L=4e-08 W=1.8e-07 
M27 8 SE 6 VNW pch L=4e-08 W=3.2e-07 
M28 22 7 8 VNW pch L=4e-08 W=1.55e-07 
M29 VDD SI 22 VNW pch L=4e-08 W=1.55e-07 
M30 9 8 VDD VNW pch L=4e-08 W=1.7e-07 
M31 10 15 9 VNW pch L=4e-08 W=1.6e-07 
M32 23 16 10 VNW pch L=4e-08 W=1.2e-07 
M33 VDD 11 23 VNW pch L=4e-08 W=1.2e-07 
M34 11 10 VDD VNW pch L=4e-08 W=2.05e-07 
M35 12 16 11 VNW pch L=4e-08 W=1.6e-07 
M36 24 15 12 VNW pch L=4e-08 W=1.2e-07 
M37 VDD 13 24 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 12 13 VNW pch L=4e-08 W=2.45e-07 
M39 QN 13 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 16 15 VNW pch L=4e-08 W=2.5e-07 
M41 16 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT ESDFFQN_X2M_A9TR QN VDD VNW VPW VSS CK D E SE SI
M0 VSS D 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.8e-07 
M2 6 E 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS 13 5 VPW nch L=4e-08 W=1.8e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.8e-07 
M7 25 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 25 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=2.5e-07 
M10 10 16 9 VPW nch L=4e-08 W=2.5e-07 
M11 26 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 26 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=2.5e-07 
M14 12 15 11 VPW nch L=4e-08 W=2.5e-07 
M15 27 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 27 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=2.5e-07 
M18 QN 13 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 13 QN VPW nch L=4e-08 W=3.1e-07 
M20 VSS 16 15 VPW nch L=4e-08 W=1.3e-07 
M21 16 CK VSS VPW nch L=4e-08 W=1.3e-07 
M22 VDD D 1 VNW pch L=4e-08 W=4e-07 
M23 4 E VDD VNW pch L=4e-08 W=3.8e-07 
M24 6 E 5 VNW pch L=4e-08 W=3.8e-07 
M25 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M26 VDD 13 5 VNW pch L=4e-08 W=3.8e-07 
M27 7 SE VDD VNW pch L=4e-08 W=1.8e-07 
M28 8 SE 6 VNW pch L=4e-08 W=3.8e-07 
M29 22 7 8 VNW pch L=4e-08 W=1.55e-07 
M30 VDD SI 22 VNW pch L=4e-08 W=1.55e-07 
M31 9 8 VDD VNW pch L=4e-08 W=2.5e-07 
M32 10 15 9 VNW pch L=4e-08 W=2.5e-07 
M33 23 16 10 VNW pch L=4e-08 W=1.2e-07 
M34 VDD 11 23 VNW pch L=4e-08 W=1.2e-07 
M35 11 10 VDD VNW pch L=4e-08 W=3.25e-07 
M36 12 16 11 VNW pch L=4e-08 W=2.5e-07 
M37 24 15 12 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 13 24 VNW pch L=4e-08 W=1.2e-07 
M39 VDD 12 13 VNW pch L=4e-08 W=3.8e-07 
M40 QN 13 VDD VNW pch L=4e-08 W=3.8e-07 
M41 VDD 13 QN VNW pch L=4e-08 W=3.8e-07 
M42 VDD 16 15 VNW pch L=4e-08 W=2.7e-07 
M43 16 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT ESDFFQN_X3M_A9TR QN VDD VNW VPW VSS CK D E SE SI
M0 VSS D 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.8e-07 
M2 6 E 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS 13 5 VPW nch L=4e-08 W=1.8e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.8e-07 
M7 25 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 25 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=3.1e-07 
M10 10 16 9 VPW nch L=4e-08 W=3.1e-07 
M11 26 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 26 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=3.1e-07 
M14 12 15 11 VPW nch L=4e-08 W=3.1e-07 
M15 27 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 27 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=2.5e-07 
M18 QN 13 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 13 QN VPW nch L=4e-08 W=3.1e-07 
M20 QN 13 VSS VPW nch L=4e-08 W=3.1e-07 
M21 VSS 16 15 VPW nch L=4e-08 W=1.4e-07 
M22 16 CK VSS VPW nch L=4e-08 W=1.4e-07 
M23 VDD D 1 VNW pch L=4e-08 W=4e-07 
M24 4 E VDD VNW pch L=4e-08 W=3.8e-07 
M25 6 E 5 VNW pch L=4e-08 W=3.8e-07 
M26 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M27 VDD 13 5 VNW pch L=4e-08 W=3.8e-07 
M28 7 SE VDD VNW pch L=4e-08 W=1.8e-07 
M29 8 SE 6 VNW pch L=4e-08 W=3.8e-07 
M30 22 7 8 VNW pch L=4e-08 W=1.55e-07 
M31 VDD SI 22 VNW pch L=4e-08 W=1.55e-07 
M32 9 8 VDD VNW pch L=4e-08 W=3.1e-07 
M33 10 15 9 VNW pch L=4e-08 W=3.1e-07 
M34 23 16 10 VNW pch L=4e-08 W=1.2e-07 
M35 VDD 11 23 VNW pch L=4e-08 W=1.2e-07 
M36 11 10 VDD VNW pch L=4e-08 W=3.8e-07 
M37 12 16 11 VNW pch L=4e-08 W=3.1e-07 
M38 24 15 12 VNW pch L=4e-08 W=1.2e-07 
M39 VDD 13 24 VNW pch L=4e-08 W=1.2e-07 
M40 VDD 12 13 VNW pch L=4e-08 W=3.8e-07 
M41 QN 13 VDD VNW pch L=4e-08 W=3.8e-07 
M42 VDD 13 QN VNW pch L=4e-08 W=3.8e-07 
M43 QN 13 VDD VNW pch L=4e-08 W=3.8e-07 
M44 VDD 16 15 VNW pch L=4e-08 W=2.9e-07 
M45 16 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT ESDFFQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D E SE SI
M0 VSS D 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.2e-07 
M2 6 E 1 VPW nch L=4e-08 W=1.2e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 13 5 VPW nch L=4e-08 W=1.2e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.2e-07 
M7 25 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 25 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=1.2e-07 
M10 10 16 9 VPW nch L=4e-08 W=1.2e-07 
M11 26 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 26 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=1.2e-07 
M14 12 15 11 VPW nch L=4e-08 W=1.2e-07 
M15 27 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 27 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 Q 12 VSS VPW nch L=4e-08 W=1.55e-07 
M19 VSS 16 15 VPW nch L=4e-08 W=1.2e-07 
M20 16 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 VDD D 1 VNW pch L=4e-08 W=2.4e-07 
M22 4 E VDD VNW pch L=4e-08 W=2.2e-07 
M23 6 E 5 VNW pch L=4e-08 W=2.2e-07 
M24 1 4 6 VNW pch L=4e-08 W=2.2e-07 
M25 VDD 13 5 VNW pch L=4e-08 W=2.2e-07 
M26 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M27 8 SE 6 VNW pch L=4e-08 W=2.2e-07 
M28 22 7 8 VNW pch L=4e-08 W=1.55e-07 
M29 VDD SI 22 VNW pch L=4e-08 W=1.55e-07 
M30 9 8 VDD VNW pch L=4e-08 W=1.3e-07 
M31 10 15 9 VNW pch L=4e-08 W=1.2e-07 
M32 23 16 10 VNW pch L=4e-08 W=1.2e-07 
M33 VDD 11 23 VNW pch L=4e-08 W=1.2e-07 
M34 11 10 VDD VNW pch L=4e-08 W=1.8e-07 
M35 12 16 11 VNW pch L=4e-08 W=1.2e-07 
M36 24 15 12 VNW pch L=4e-08 W=1.2e-07 
M37 VDD 13 24 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 12 13 VNW pch L=4e-08 W=1.2e-07 
M39 Q 12 VDD VNW pch L=4e-08 W=2e-07 
M40 VDD 16 15 VNW pch L=4e-08 W=2.5e-07 
M41 16 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT ESDFFQ_X1M_A9TR Q VDD VNW VPW VSS CK D E SE SI
M0 VSS D 1 VPW nch L=4e-08 W=1.6e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.6e-07 
M2 6 E 1 VPW nch L=4e-08 W=1.6e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.6e-07 
M4 VSS 13 5 VPW nch L=4e-08 W=1.6e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.6e-07 
M7 25 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 25 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=1.6e-07 
M10 10 16 9 VPW nch L=4e-08 W=1.6e-07 
M11 26 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 26 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=1.6e-07 
M14 12 15 11 VPW nch L=4e-08 W=1.6e-07 
M15 27 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 27 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 16 15 VPW nch L=4e-08 W=1.2e-07 
M20 16 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 VDD D 1 VNW pch L=4e-08 W=3.4e-07 
M22 4 E VDD VNW pch L=4e-08 W=3.2e-07 
M23 6 E 5 VNW pch L=4e-08 W=3.2e-07 
M24 1 4 6 VNW pch L=4e-08 W=3.2e-07 
M25 VDD 13 5 VNW pch L=4e-08 W=3.2e-07 
M26 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M27 8 SE 6 VNW pch L=4e-08 W=3.2e-07 
M28 22 7 8 VNW pch L=4e-08 W=1.55e-07 
M29 VDD SI 22 VNW pch L=4e-08 W=1.55e-07 
M30 9 8 VDD VNW pch L=4e-08 W=1.75e-07 
M31 10 15 9 VNW pch L=4e-08 W=1.6e-07 
M32 23 16 10 VNW pch L=4e-08 W=1.2e-07 
M33 VDD 11 23 VNW pch L=4e-08 W=1.2e-07 
M34 11 10 VDD VNW pch L=4e-08 W=2.3e-07 
M35 12 16 11 VNW pch L=4e-08 W=1.6e-07 
M36 24 15 12 VNW pch L=4e-08 W=1.2e-07 
M37 VDD 13 24 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 12 13 VNW pch L=4e-08 W=1.2e-07 
M39 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 16 15 VNW pch L=4e-08 W=2.5e-07 
M41 16 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT ESDFFQ_X2M_A9TR Q VDD VNW VPW VSS CK D E SE SI
M0 VSS D 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.8e-07 
M2 6 E 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS 13 5 VPW nch L=4e-08 W=1.8e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.8e-07 
M7 25 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 25 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=2.5e-07 
M10 10 16 9 VPW nch L=4e-08 W=2.5e-07 
M11 26 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 26 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=2.5e-07 
M14 12 15 11 VPW nch L=4e-08 W=2.5e-07 
M15 27 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 27 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 12 Q VPW nch L=4e-08 W=3.1e-07 
M20 VSS 16 15 VPW nch L=4e-08 W=1.3e-07 
M21 16 CK VSS VPW nch L=4e-08 W=1.3e-07 
M22 VDD D 1 VNW pch L=4e-08 W=4e-07 
M23 4 E VDD VNW pch L=4e-08 W=3.8e-07 
M24 6 E 5 VNW pch L=4e-08 W=3.8e-07 
M25 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M26 VDD 13 5 VNW pch L=4e-08 W=3.8e-07 
M27 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M28 8 SE 6 VNW pch L=4e-08 W=3.8e-07 
M29 22 7 8 VNW pch L=4e-08 W=1.55e-07 
M30 VDD SI 22 VNW pch L=4e-08 W=1.55e-07 
M31 9 8 VDD VNW pch L=4e-08 W=2.7e-07 
M32 10 15 9 VNW pch L=4e-08 W=2.5e-07 
M33 23 16 10 VNW pch L=4e-08 W=1.2e-07 
M34 VDD 11 23 VNW pch L=4e-08 W=1.2e-07 
M35 11 10 VDD VNW pch L=4e-08 W=3.35e-07 
M36 12 16 11 VNW pch L=4e-08 W=2.5e-07 
M37 24 15 12 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 13 24 VNW pch L=4e-08 W=1.2e-07 
M39 VDD 12 13 VNW pch L=4e-08 W=1.2e-07 
M40 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M41 VDD 12 Q VNW pch L=4e-08 W=3.8e-07 
M42 VDD 16 15 VNW pch L=4e-08 W=2.7e-07 
M43 16 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT ESDFFQ_X3M_A9TR Q VDD VNW VPW VSS CK D E SE SI
M0 VSS D 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.8e-07 
M2 6 E 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS 13 5 VPW nch L=4e-08 W=1.8e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.8e-07 
M7 25 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 25 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=3.1e-07 
M10 10 16 9 VPW nch L=4e-08 W=3.1e-07 
M11 26 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 26 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=3.1e-07 
M14 12 15 11 VPW nch L=4e-08 W=3.1e-07 
M15 27 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 27 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 12 Q VPW nch L=4e-08 W=3.1e-07 
M20 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M21 VSS 16 15 VPW nch L=4e-08 W=1.4e-07 
M22 16 CK VSS VPW nch L=4e-08 W=1.4e-07 
M23 VDD D 1 VNW pch L=4e-08 W=4e-07 
M24 4 E VDD VNW pch L=4e-08 W=3.8e-07 
M25 6 E 5 VNW pch L=4e-08 W=3.8e-07 
M26 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M27 VDD 13 5 VNW pch L=4e-08 W=3.8e-07 
M28 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M29 8 SE 6 VNW pch L=4e-08 W=3.8e-07 
M30 22 7 8 VNW pch L=4e-08 W=1.55e-07 
M31 VDD SI 22 VNW pch L=4e-08 W=1.55e-07 
M32 9 8 VDD VNW pch L=4e-08 W=3.3e-07 
M33 10 15 9 VNW pch L=4e-08 W=3.1e-07 
M34 23 16 10 VNW pch L=4e-08 W=1.2e-07 
M35 VDD 11 23 VNW pch L=4e-08 W=1.2e-07 
M36 11 10 VDD VNW pch L=4e-08 W=3.8e-07 
M37 12 16 11 VNW pch L=4e-08 W=3.1e-07 
M38 24 15 12 VNW pch L=4e-08 W=1.2e-07 
M39 VDD 13 24 VNW pch L=4e-08 W=1.2e-07 
M40 VDD 12 13 VNW pch L=4e-08 W=1.2e-07 
M41 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M42 VDD 12 Q VNW pch L=4e-08 W=3.8e-07 
M43 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M44 VDD 16 15 VNW pch L=4e-08 W=2.9e-07 
M45 16 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS










.SUBCKT FILLCAP128_A9TR VDD VNW VPW VSS
M0 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M1 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M2 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M3 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M4 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M5 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M6 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M7 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M8 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M9 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M10 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M11 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M12 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M13 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M14 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M15 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M16 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M17 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M18 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M19 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M20 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M21 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M22 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M23 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M24 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M25 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M26 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M27 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M28 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M29 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M30 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M31 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M32 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M33 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M34 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M35 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M36 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M37 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M38 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M39 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M40 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M41 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M42 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M43 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M44 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M45 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M46 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M47 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M48 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M49 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M50 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M51 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M52 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M53 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M54 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M55 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M56 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M57 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M58 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M59 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M60 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M61 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M62 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M63 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
.ENDS


.SUBCKT FILLCAP16_A9TR VDD VNW VPW VSS
M0 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M1 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M2 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M3 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M4 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M5 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M6 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M7 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
.ENDS


.SUBCKT FILLCAP32_A9TR VDD VNW VPW VSS
M0 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M1 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M2 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M3 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M4 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M5 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M6 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M7 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M8 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M9 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M10 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M11 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M12 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M13 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M14 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M15 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
.ENDS


.SUBCKT FILLCAP4_A9TR VDD VNW VPW VSS
M0 VSS VDD VSS VPW nch L=3.5e-07 W=2.4e-07 
M1 VDD VSS VDD VNW pch L=3.5e-07 W=2.4e-07 
.ENDS


.SUBCKT FILLCAP64_A9TR VDD VNW VPW VSS
M0 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M1 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M2 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M3 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M4 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M5 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M6 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M7 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M8 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M9 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M10 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M11 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M12 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M13 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M14 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M15 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M16 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M17 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M18 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M19 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M20 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M21 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M22 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M23 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M24 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M25 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M26 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M27 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M28 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M29 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M30 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M31 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
.ENDS


.SUBCKT FILLCAP8_A9TR VDD VNW VPW VSS
M0 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M1 VSS VDD VSS VPW nch L=3.2e-07 W=2e-07 
M2 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
M3 VDD VSS VDD VNW pch L=3.2e-07 W=2e-07 
.ENDS


.SUBCKT FILLSGCAP128_A9TR VDD VNW VPW VSS
M0 VSS 4 VSS VPW nch L=3e-07 W=3.4e-07 
M1 VSS 6 VSS VPW nch L=3e-07 W=3.4e-07 
M2 VSS 8 VSS VPW nch L=3e-07 W=3.4e-07 
M3 VSS 10 VSS VPW nch L=3e-07 W=3.4e-07 
M4 VSS 12 VSS VPW nch L=3e-07 W=3.4e-07 
M5 VSS 14 VSS VPW nch L=3e-07 W=3.4e-07 
M6 VSS 16 VSS VPW nch L=3e-07 W=3.4e-07 
M7 VSS 18 VSS VPW nch L=3e-07 W=3.4e-07 
M8 VSS 20 VSS VPW nch L=3e-07 W=3.4e-07 
M9 VSS 22 VSS VPW nch L=3e-07 W=3.4e-07 
M10 VSS 24 VSS VPW nch L=3e-07 W=3.4e-07 
M11 VSS 26 VSS VPW nch L=3e-07 W=3.4e-07 
M12 VSS 28 VSS VPW nch L=3e-07 W=3.4e-07 
M13 VSS 30 VSS VPW nch L=3e-07 W=3.4e-07 
M14 VSS 32 VSS VPW nch L=3e-07 W=3.4e-07 
M15 VSS 34 VSS VPW nch L=3e-07 W=3.4e-07 
M16 VSS 36 VSS VPW nch L=3e-07 W=3.4e-07 
M17 VSS 38 VSS VPW nch L=3e-07 W=3.4e-07 
M18 VSS 40 VSS VPW nch L=3e-07 W=3.4e-07 
M19 VSS 42 VSS VPW nch L=3e-07 W=3.4e-07 
M20 VSS 44 VSS VPW nch L=3e-07 W=3.4e-07 
M21 VSS 46 VSS VPW nch L=3e-07 W=3.4e-07 
M22 VSS 48 VSS VPW nch L=3e-07 W=3.4e-07 
M23 VSS 50 VSS VPW nch L=3e-07 W=3.4e-07 
M24 VSS 52 VSS VPW nch L=3e-07 W=3.4e-07 
M25 VSS 54 VSS VPW nch L=3e-07 W=3.4e-07 
M26 VSS 56 VSS VPW nch L=3e-07 W=3.4e-07 
M27 VSS 58 VSS VPW nch L=3e-07 W=3.4e-07 
M28 VSS 60 VSS VPW nch L=3e-07 W=3.4e-07 
M29 VSS 62 VSS VPW nch L=3e-07 W=3.4e-07 
M30 VSS 64 VSS VPW nch L=3e-07 W=3.4e-07 
M31 VSS 66 VSS VPW nch L=3e-07 W=3.4e-07 
M32 VDD 4 VDD VNW pch L=3e-07 W=3.4e-07 
M33 VDD 6 VDD VNW pch L=3e-07 W=3.4e-07 
M34 VDD 8 VDD VNW pch L=3e-07 W=3.4e-07 
M35 VDD 10 VDD VNW pch L=3e-07 W=3.4e-07 
M36 VDD 12 VDD VNW pch L=3e-07 W=3.4e-07 
M37 VDD 14 VDD VNW pch L=3e-07 W=3.4e-07 
M38 VDD 16 VDD VNW pch L=3e-07 W=3.4e-07 
M39 VDD 18 VDD VNW pch L=3e-07 W=3.4e-07 
M40 VDD 20 VDD VNW pch L=3e-07 W=3.4e-07 
M41 VDD 22 VDD VNW pch L=3e-07 W=3.4e-07 
M42 VDD 24 VDD VNW pch L=3e-07 W=3.4e-07 
M43 VDD 26 VDD VNW pch L=3e-07 W=3.4e-07 
M44 VDD 28 VDD VNW pch L=3e-07 W=3.4e-07 
M45 VDD 30 VDD VNW pch L=3e-07 W=3.4e-07 
M46 VDD 32 VDD VNW pch L=3e-07 W=3.4e-07 
M47 VDD 34 VDD VNW pch L=3e-07 W=3.4e-07 
M48 VDD 36 VDD VNW pch L=3e-07 W=3.4e-07 
M49 VDD 38 VDD VNW pch L=3e-07 W=3.4e-07 
M50 VDD 40 VDD VNW pch L=3e-07 W=3.4e-07 
M51 VDD 42 VDD VNW pch L=3e-07 W=3.4e-07 
M52 VDD 44 VDD VNW pch L=3e-07 W=3.4e-07 
M53 VDD 46 VDD VNW pch L=3e-07 W=3.4e-07 
M54 VDD 48 VDD VNW pch L=3e-07 W=3.4e-07 
M55 VDD 50 VDD VNW pch L=3e-07 W=3.4e-07 
M56 VDD 52 VDD VNW pch L=3e-07 W=3.4e-07 
M57 VDD 54 VDD VNW pch L=3e-07 W=3.4e-07 
M58 VDD 56 VDD VNW pch L=3e-07 W=3.4e-07 
M59 VDD 58 VDD VNW pch L=3e-07 W=3.4e-07 
M60 VDD 60 VDD VNW pch L=3e-07 W=3.4e-07 
M61 VDD 62 VDD VNW pch L=3e-07 W=3.4e-07 
M62 VDD 64 VDD VNW pch L=3e-07 W=3.4e-07 
M63 VDD 66 VDD VNW pch L=3e-07 W=3.4e-07 
.ENDS


.SUBCKT FILLSGCAP16_A9TR VDD VNW VPW VSS
M0 VSS 4 VSS VPW nch L=3e-07 W=3.4e-07 
M1 VSS 6 VSS VPW nch L=3e-07 W=3.4e-07 
M2 VSS 8 VSS VPW nch L=3e-07 W=3.4e-07 
M3 VSS 10 VSS VPW nch L=3e-07 W=3.4e-07 
M4 VDD 4 VDD VNW pch L=3e-07 W=3.4e-07 
M5 VDD 6 VDD VNW pch L=3e-07 W=3.4e-07 
M6 VDD 8 VDD VNW pch L=3e-07 W=3.4e-07 
M7 VDD 10 VDD VNW pch L=3e-07 W=3.4e-07 
.ENDS


.SUBCKT FILLSGCAP32_A9TR VDD VNW VPW VSS
M0 VSS 4 VSS VPW nch L=3e-07 W=3.4e-07 
M1 VSS 6 VSS VPW nch L=3e-07 W=3.4e-07 
M2 VSS 8 VSS VPW nch L=3e-07 W=3.4e-07 
M3 VSS 10 VSS VPW nch L=3e-07 W=3.4e-07 
M4 VSS 12 VSS VPW nch L=3e-07 W=3.4e-07 
M5 VSS 14 VSS VPW nch L=3e-07 W=3.4e-07 
M6 VSS 16 VSS VPW nch L=3e-07 W=3.4e-07 
M7 VSS 18 VSS VPW nch L=3e-07 W=3.4e-07 
M8 VDD 4 VDD VNW pch L=3e-07 W=3.4e-07 
M9 VDD 6 VDD VNW pch L=3e-07 W=3.4e-07 
M10 VDD 8 VDD VNW pch L=3e-07 W=3.4e-07 
M11 VDD 10 VDD VNW pch L=3e-07 W=3.4e-07 
M12 VDD 12 VDD VNW pch L=3e-07 W=3.4e-07 
M13 VDD 14 VDD VNW pch L=3e-07 W=3.4e-07 
M14 VDD 16 VDD VNW pch L=3e-07 W=3.4e-07 
M15 VDD 18 VDD VNW pch L=3e-07 W=3.4e-07 
.ENDS


.SUBCKT FILLSGCAP4_A9TR VDD VNW VPW VSS
M0 VSS 4 VSS VPW nch L=3e-07 W=3.4e-07 
M1 VDD 4 VDD VNW pch L=3e-07 W=3.4e-07 
.ENDS


.SUBCKT FILLSGCAP64_A9TR VDD VNW VPW VSS
M0 VSS 4 VSS VPW nch L=3e-07 W=3.4e-07 
M1 VSS 6 VSS VPW nch L=3e-07 W=3.4e-07 
M2 VSS 8 VSS VPW nch L=3e-07 W=3.4e-07 
M3 VSS 10 VSS VPW nch L=3e-07 W=3.4e-07 
M4 VSS 12 VSS VPW nch L=3e-07 W=3.4e-07 
M5 VSS 14 VSS VPW nch L=3e-07 W=3.4e-07 
M6 VSS 16 VSS VPW nch L=3e-07 W=3.4e-07 
M7 VSS 18 VSS VPW nch L=3e-07 W=3.4e-07 
M8 VSS 20 VSS VPW nch L=3e-07 W=3.4e-07 
M9 VSS 22 VSS VPW nch L=3e-07 W=3.4e-07 
M10 VSS 24 VSS VPW nch L=3e-07 W=3.4e-07 
M11 VSS 26 VSS VPW nch L=3e-07 W=3.4e-07 
M12 VSS 28 VSS VPW nch L=3e-07 W=3.4e-07 
M13 VSS 30 VSS VPW nch L=3e-07 W=3.4e-07 
M14 VSS 32 VSS VPW nch L=3e-07 W=3.4e-07 
M15 VSS 34 VSS VPW nch L=3e-07 W=3.4e-07 
M16 VDD 4 VDD VNW pch L=3e-07 W=3.4e-07 
M17 VDD 6 VDD VNW pch L=3e-07 W=3.4e-07 
M18 VDD 8 VDD VNW pch L=3e-07 W=3.4e-07 
M19 VDD 10 VDD VNW pch L=3e-07 W=3.4e-07 
M20 VDD 12 VDD VNW pch L=3e-07 W=3.4e-07 
M21 VDD 14 VDD VNW pch L=3e-07 W=3.4e-07 
M22 VDD 16 VDD VNW pch L=3e-07 W=3.4e-07 
M23 VDD 18 VDD VNW pch L=3e-07 W=3.4e-07 
M24 VDD 20 VDD VNW pch L=3e-07 W=3.4e-07 
M25 VDD 22 VDD VNW pch L=3e-07 W=3.4e-07 
M26 VDD 24 VDD VNW pch L=3e-07 W=3.4e-07 
M27 VDD 26 VDD VNW pch L=3e-07 W=3.4e-07 
M28 VDD 28 VDD VNW pch L=3e-07 W=3.4e-07 
M29 VDD 30 VDD VNW pch L=3e-07 W=3.4e-07 
M30 VDD 32 VDD VNW pch L=3e-07 W=3.4e-07 
M31 VDD 34 VDD VNW pch L=3e-07 W=3.4e-07 
.ENDS


.SUBCKT FILLSGCAP8_A9TR VDD VNW VPW VSS
M0 VSS 4 VSS VPW nch L=3e-07 W=3.4e-07 
M1 VSS 6 VSS VPW nch L=3e-07 W=3.4e-07 
M2 VDD 4 VDD VNW pch L=3e-07 W=3.4e-07 
M3 VDD 6 VDD VNW pch L=3e-07 W=3.4e-07 
.ENDS



.SUBCKT FRICG_X0P5B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 CK 5 VPW nch L=4e-08 W=1.2e-07 
M2 VSS 4 8 VPW nch L=4e-08 W=1.2e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=1.2e-07 
M4 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M6 5 CK VDD VNW pch L=4e-08 W=1.4e-07 
M7 VDD 4 5 VNW pch L=4e-08 W=1.2e-07 
M8 ECK 5 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT FRICG_X0P6B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 CK 5 VPW nch L=4e-08 W=1.2e-07 
M2 VSS 4 8 VPW nch L=4e-08 W=1.2e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=1.35e-07 
M4 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M6 5 CK VDD VNW pch L=4e-08 W=1.4e-07 
M7 VDD 4 5 VNW pch L=4e-08 W=1.2e-07 
M8 ECK 5 VDD VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT FRICG_X0P7B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 CK 5 VPW nch L=4e-08 W=1.2e-07 
M2 VSS 4 8 VPW nch L=4e-08 W=1.2e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=1.6e-07 
M4 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M6 5 CK VDD VNW pch L=4e-08 W=1.4e-07 
M7 VDD 4 5 VNW pch L=4e-08 W=1.2e-07 
M8 ECK 5 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT FRICG_X0P8B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 CK 5 VPW nch L=4e-08 W=1.2e-07 
M2 VSS 4 8 VPW nch L=4e-08 W=1.2e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=1.9e-07 
M4 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M6 5 CK VDD VNW pch L=4e-08 W=1.4e-07 
M7 VDD 4 5 VNW pch L=4e-08 W=1.2e-07 
M8 ECK 5 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT FRICG_X11B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 CK 5 VPW nch L=4e-08 W=3.4e-07 
M2 VSS 4 8 VPW nch L=4e-08 W=3.4e-07 
M3 9 4 VSS VPW nch L=4e-08 W=3.4e-07 
M4 5 CK 9 VPW nch L=4e-08 W=3.4e-07 
M5 10 CK 5 VPW nch L=4e-08 W=3.4e-07 
M6 VSS 4 10 VPW nch L=4e-08 W=3.4e-07 
M7 VSS 5 ECK VPW nch L=4e-08 W=3.55e-07 
M8 ECK 5 VSS VPW nch L=4e-08 W=3.55e-07 
M9 VSS 5 ECK VPW nch L=4e-08 W=3.55e-07 
M10 ECK 5 VSS VPW nch L=4e-08 W=3.55e-07 
M11 VSS 5 ECK VPW nch L=4e-08 W=3.55e-07 
M12 ECK 5 VSS VPW nch L=4e-08 W=3.55e-07 
M13 VSS 5 ECK VPW nch L=4e-08 W=3.55e-07 
M14 4 1 VDD VNW pch L=4e-08 W=2.9e-07 
M15 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M16 5 CK VDD VNW pch L=4e-08 W=2.25e-07 
M17 VDD CK 5 VNW pch L=4e-08 W=2.25e-07 
M18 5 CK VDD VNW pch L=4e-08 W=2.25e-07 
M19 VDD CK 5 VNW pch L=4e-08 W=2.25e-07 
M20 5 CK VDD VNW pch L=4e-08 W=2.25e-07 
M21 VDD 4 5 VNW pch L=4e-08 W=1.2e-07 
M22 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M23 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M25 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M27 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M29 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M31 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT FRICG_X13B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 3 2 VPW nch L=4e-08 W=1.2e-07 
M1 9 3 VSS VPW nch L=4e-08 W=3e-07 
M2 5 CK 9 VPW nch L=4e-08 W=3e-07 
M3 10 CK 5 VPW nch L=4e-08 W=3e-07 
M4 VSS 3 10 VPW nch L=4e-08 W=3e-07 
M5 11 3 VSS VPW nch L=4e-08 W=3e-07 
M6 5 CK 11 VPW nch L=4e-08 W=3e-07 
M7 12 CK 5 VPW nch L=4e-08 W=3e-07 
M8 VSS 3 12 VPW nch L=4e-08 W=3e-07 
M9 VSS 5 ECK VPW nch L=4e-08 W=3.25e-07 
M10 ECK 5 VSS VPW nch L=4e-08 W=3.25e-07 
M11 VSS 5 ECK VPW nch L=4e-08 W=3.25e-07 
M12 ECK 5 VSS VPW nch L=4e-08 W=3.25e-07 
M13 VSS 5 ECK VPW nch L=4e-08 W=3.25e-07 
M14 ECK 5 VSS VPW nch L=4e-08 W=3.25e-07 
M15 VSS 5 ECK VPW nch L=4e-08 W=3.25e-07 
M16 ECK 5 VSS VPW nch L=4e-08 W=3.25e-07 
M17 VSS 5 ECK VPW nch L=4e-08 W=3.25e-07 
M18 3 2 VDD VNW pch L=4e-08 W=3.4e-07 
M19 VDD 3 3 VNW pch L=4e-08 W=1.55e-07 
M20 5 CK VDD VNW pch L=4e-08 W=2.3e-07 
M21 VDD CK 5 VNW pch L=4e-08 W=2.3e-07 
M22 5 CK VDD VNW pch L=4e-08 W=2.3e-07 
M23 VDD CK 5 VNW pch L=4e-08 W=2.3e-07 
M24 5 CK VDD VNW pch L=4e-08 W=2.3e-07 
M25 VDD CK 5 VNW pch L=4e-08 W=2.3e-07 
M26 5 3 VDD VNW pch L=4e-08 W=1.4e-07 
M27 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M28 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M30 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M32 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M33 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M34 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M36 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M38 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT FRICG_X16B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 3 2 VPW nch L=4e-08 W=1.2e-07 
M1 9 3 VSS VPW nch L=4e-08 W=3.5e-07 
M2 5 CK 9 VPW nch L=4e-08 W=3.5e-07 
M3 10 CK 5 VPW nch L=4e-08 W=3.5e-07 
M4 VSS 3 10 VPW nch L=4e-08 W=3.5e-07 
M5 11 3 VSS VPW nch L=4e-08 W=3.5e-07 
M6 5 CK 11 VPW nch L=4e-08 W=3.5e-07 
M7 12 CK 5 VPW nch L=4e-08 W=3.5e-07 
M8 VSS 3 12 VPW nch L=4e-08 W=3.5e-07 
M9 ECK 5 VSS VPW nch L=4e-08 W=3.6e-07 
M10 VSS 5 ECK VPW nch L=4e-08 W=3.6e-07 
M11 ECK 5 VSS VPW nch L=4e-08 W=3.6e-07 
M12 VSS 5 ECK VPW nch L=4e-08 W=3.6e-07 
M13 ECK 5 VSS VPW nch L=4e-08 W=3.6e-07 
M14 VSS 5 ECK VPW nch L=4e-08 W=3.6e-07 
M15 ECK 5 VSS VPW nch L=4e-08 W=3.6e-07 
M16 VSS 5 ECK VPW nch L=4e-08 W=3.6e-07 
M17 ECK 5 VSS VPW nch L=4e-08 W=3.6e-07 
M18 VSS 5 ECK VPW nch L=4e-08 W=3.6e-07 
M19 3 3 VDD VNW pch L=4e-08 W=1.55e-07 
M20 VDD 2 3 VNW pch L=4e-08 W=4e-07 
M21 5 CK VDD VNW pch L=4e-08 W=2.35e-07 
M22 VDD CK 5 VNW pch L=4e-08 W=2.35e-07 
M23 5 CK VDD VNW pch L=4e-08 W=2.35e-07 
M24 VDD CK 5 VNW pch L=4e-08 W=2.35e-07 
M25 5 CK VDD VNW pch L=4e-08 W=2.35e-07 
M26 VDD CK 5 VNW pch L=4e-08 W=2.35e-07 
M27 5 CK VDD VNW pch L=4e-08 W=2.35e-07 
M28 VDD 3 5 VNW pch L=4e-08 W=1.65e-07 
M29 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M31 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M33 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M35 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M37 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M39 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M41 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M42 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M43 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M44 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT FRICG_X1B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 4 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 CK 8 VPW nch L=4e-08 W=1.2e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=2.25e-07 
M4 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M6 5 4 VDD VNW pch L=4e-08 W=1.2e-07 
M7 VDD CK 5 VNW pch L=4e-08 W=1.4e-07 
M8 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT FRICG_X1P2B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 4 VSS VPW nch L=4e-08 W=1.45e-07 
M2 5 CK 8 VPW nch L=4e-08 W=1.45e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=2.7e-07 
M4 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M6 5 4 VDD VNW pch L=4e-08 W=1.2e-07 
M7 VDD CK 5 VNW pch L=4e-08 W=1.7e-07 
M8 ECK 5 VDD VNW pch L=4e-08 W=2.4e-07 
M9 VDD 5 ECK VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT FRICG_X1P4B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 4 VSS VPW nch L=4e-08 W=1.6e-07 
M2 5 CK 8 VPW nch L=4e-08 W=1.6e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=3.2e-07 
M4 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M6 5 4 VDD VNW pch L=4e-08 W=1.2e-07 
M7 VDD CK 5 VNW pch L=4e-08 W=1.9e-07 
M8 ECK 5 VDD VNW pch L=4e-08 W=2.85e-07 
M9 VDD 5 ECK VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT FRICG_X1P7B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 4 VSS VPW nch L=4e-08 W=1.8e-07 
M2 5 CK 8 VPW nch L=4e-08 W=1.8e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=3.8e-07 
M4 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M6 5 4 VDD VNW pch L=4e-08 W=1.2e-07 
M7 VDD CK 5 VNW pch L=4e-08 W=2.1e-07 
M8 ECK 5 VDD VNW pch L=4e-08 W=3.35e-07 
M9 VDD 5 ECK VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT FRICG_X2B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 4 VSS VPW nch L=4e-08 W=2.1e-07 
M2 5 CK 8 VPW nch L=4e-08 W=2.1e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=2.25e-07 
M4 VSS 5 ECK VPW nch L=4e-08 W=2.25e-07 
M5 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M6 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M7 5 4 VDD VNW pch L=4e-08 W=1.2e-07 
M8 VDD CK 5 VNW pch L=4e-08 W=2.4e-07 
M9 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT FRICG_X2P5B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 3 2 VPW nch L=4e-08 W=1.2e-07 
M1 9 3 VSS VPW nch L=4e-08 W=2.55e-07 
M2 5 CK 9 VPW nch L=4e-08 W=2.55e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=2.85e-07 
M4 VSS 5 ECK VPW nch L=4e-08 W=2.85e-07 
M5 3 2 VDD VNW pch L=4e-08 W=1.2e-07 
M6 VDD 3 3 VNW pch L=4e-08 W=1.55e-07 
M7 5 3 VDD VNW pch L=4e-08 W=1.2e-07 
M8 VDD CK 5 VNW pch L=4e-08 W=2.95e-07 
M9 ECK 5 VDD VNW pch L=4e-08 W=3.35e-07 
M10 VDD 5 ECK VNW pch L=4e-08 W=3.35e-07 
M11 ECK 5 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT FRICG_X3B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 3 2 VPW nch L=4e-08 W=1.2e-07 
M1 9 3 VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 CK 9 VPW nch L=4e-08 W=2.9e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=3.4e-07 
M4 VSS 5 ECK VPW nch L=4e-08 W=3.4e-07 
M5 3 2 VDD VNW pch L=4e-08 W=1.2e-07 
M6 VDD 3 3 VNW pch L=4e-08 W=1.55e-07 
M7 5 3 VDD VNW pch L=4e-08 W=1.2e-07 
M8 VDD CK 5 VNW pch L=4e-08 W=3.4e-07 
M9 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M11 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT FRICG_X3P5B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 4 VSS VPW nch L=4e-08 W=3.2e-07 
M2 5 CK 8 VPW nch L=4e-08 W=3.2e-07 
M3 ECK 5 VSS VPW nch L=4e-08 W=2e-07 
M4 VSS 5 ECK VPW nch L=4e-08 W=2e-07 
M5 ECK 5 VSS VPW nch L=4e-08 W=2e-07 
M6 VSS 5 ECK VPW nch L=4e-08 W=2e-07 
M7 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M8 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M9 5 4 VDD VNW pch L=4e-08 W=1.2e-07 
M10 VDD CK 5 VNW pch L=4e-08 W=3.65e-07 
M11 ECK 5 VDD VNW pch L=4e-08 W=3.5e-07 
M12 VDD 5 ECK VNW pch L=4e-08 W=3.5e-07 
M13 ECK 5 VDD VNW pch L=4e-08 W=3.5e-07 
M14 VDD 5 ECK VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT FRICG_X4B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 4 VSS VPW nch L=4e-08 W=2.05e-07 
M2 5 CK 8 VPW nch L=4e-08 W=2.05e-07 
M3 9 CK 5 VPW nch L=4e-08 W=2.05e-07 
M4 VSS 4 9 VPW nch L=4e-08 W=2.05e-07 
M5 VSS 5 ECK VPW nch L=4e-08 W=3e-07 
M6 ECK 5 VSS VPW nch L=4e-08 W=3e-07 
M7 VSS 5 ECK VPW nch L=4e-08 W=3e-07 
M8 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M9 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M10 5 CK VDD VNW pch L=4e-08 W=2.4e-07 
M11 VDD CK 5 VNW pch L=4e-08 W=2.4e-07 
M12 5 4 VDD VNW pch L=4e-08 W=1.2e-07 
M13 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M15 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT FRICG_X5B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 3 2 VPW nch L=4e-08 W=1.2e-07 
M1 9 3 VSS VPW nch L=4e-08 W=2.5e-07 
M2 5 CK 9 VPW nch L=4e-08 W=2.5e-07 
M3 10 CK 5 VPW nch L=4e-08 W=2.5e-07 
M4 VSS 3 10 VPW nch L=4e-08 W=2.5e-07 
M5 VSS 5 ECK VPW nch L=4e-08 W=2.25e-07 
M6 ECK 5 VSS VPW nch L=4e-08 W=2.25e-07 
M7 VSS 5 ECK VPW nch L=4e-08 W=2.25e-07 
M8 ECK 5 VSS VPW nch L=4e-08 W=2.25e-07 
M9 VSS 5 ECK VPW nch L=4e-08 W=2.25e-07 
M10 3 2 VDD VNW pch L=4e-08 W=1.4e-07 
M11 VDD 3 3 VNW pch L=4e-08 W=1.55e-07 
M12 5 CK VDD VNW pch L=4e-08 W=2e-07 
M13 VDD CK 5 VNW pch L=4e-08 W=2e-07 
M14 5 CK VDD VNW pch L=4e-08 W=2e-07 
M15 VDD 3 5 VNW pch L=4e-08 W=1.2e-07 
M16 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M17 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M19 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT FRICG_X6B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 3 2 VPW nch L=4e-08 W=1.2e-07 
M1 9 3 VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 CK 9 VPW nch L=4e-08 W=2.9e-07 
M3 10 CK 5 VPW nch L=4e-08 W=2.9e-07 
M4 VSS 3 10 VPW nch L=4e-08 W=2.9e-07 
M5 ECK 5 VSS VPW nch L=4e-08 W=3.35e-07 
M6 VSS 5 ECK VPW nch L=4e-08 W=3.35e-07 
M7 ECK 5 VSS VPW nch L=4e-08 W=3.35e-07 
M8 VSS 5 ECK VPW nch L=4e-08 W=3.35e-07 
M9 3 2 VDD VNW pch L=4e-08 W=1.65e-07 
M10 VDD 3 3 VNW pch L=4e-08 W=1.55e-07 
M11 5 CK VDD VNW pch L=4e-08 W=2.25e-07 
M12 VDD CK 5 VNW pch L=4e-08 W=2.25e-07 
M13 5 CK VDD VNW pch L=4e-08 W=2.25e-07 
M14 VDD 3 5 VNW pch L=4e-08 W=1.2e-07 
M15 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M17 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M19 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT FRICG_X7P5B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 CK 5 VPW nch L=4e-08 W=2.45e-07 
M2 VSS 4 8 VPW nch L=4e-08 W=2.45e-07 
M3 9 4 VSS VPW nch L=4e-08 W=2.45e-07 
M4 5 CK 9 VPW nch L=4e-08 W=2.45e-07 
M5 10 CK 5 VPW nch L=4e-08 W=2.45e-07 
M6 VSS 4 10 VPW nch L=4e-08 W=2.45e-07 
M7 ECK 5 VSS VPW nch L=4e-08 W=2.85e-07 
M8 VSS 5 ECK VPW nch L=4e-08 W=2.85e-07 
M9 ECK 5 VSS VPW nch L=4e-08 W=2.85e-07 
M10 VSS 5 ECK VPW nch L=4e-08 W=2.85e-07 
M11 ECK 5 VSS VPW nch L=4e-08 W=2.85e-07 
M12 VSS 5 ECK VPW nch L=4e-08 W=2.85e-07 
M13 4 1 VDD VNW pch L=4e-08 W=2.1e-07 
M14 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M15 5 CK VDD VNW pch L=4e-08 W=2.15e-07 
M16 VDD CK 5 VNW pch L=4e-08 W=2.15e-07 
M17 5 CK VDD VNW pch L=4e-08 W=2.15e-07 
M18 VDD CK 5 VNW pch L=4e-08 W=2.15e-07 
M19 5 4 VDD VNW pch L=4e-08 W=1.2e-07 
M20 ECK 5 VDD VNW pch L=4e-08 W=3.75e-07 
M21 VDD 5 ECK VNW pch L=4e-08 W=3.75e-07 
M22 ECK 5 VDD VNW pch L=4e-08 W=3.75e-07 
M23 VDD 5 ECK VNW pch L=4e-08 W=3.75e-07 
M24 ECK 5 VDD VNW pch L=4e-08 W=3.75e-07 
M25 VDD 5 ECK VNW pch L=4e-08 W=3.75e-07 
M26 ECK 5 VDD VNW pch L=4e-08 W=3.75e-07 
M27 VDD 5 ECK VNW pch L=4e-08 W=3.75e-07 
.ENDS


.SUBCKT FRICG_X9B_A9TR ECK VDD VNW VPW VSS CK
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 CK 5 VPW nch L=4e-08 W=2.75e-07 
M2 VSS 4 8 VPW nch L=4e-08 W=2.75e-07 
M3 9 4 VSS VPW nch L=4e-08 W=2.75e-07 
M4 5 CK 9 VPW nch L=4e-08 W=2.75e-07 
M5 10 CK 5 VPW nch L=4e-08 W=2.75e-07 
M6 VSS 4 10 VPW nch L=4e-08 W=2.75e-07 
M7 VSS 5 ECK VPW nch L=4e-08 W=2.9e-07 
M8 ECK 5 VSS VPW nch L=4e-08 W=2.9e-07 
M9 VSS 5 ECK VPW nch L=4e-08 W=2.9e-07 
M10 ECK 5 VSS VPW nch L=4e-08 W=2.9e-07 
M11 VSS 5 ECK VPW nch L=4e-08 W=2.9e-07 
M12 ECK 5 VSS VPW nch L=4e-08 W=2.9e-07 
M13 VSS 5 ECK VPW nch L=4e-08 W=2.9e-07 
M14 4 1 VDD VNW pch L=4e-08 W=2.4e-07 
M15 VDD 4 4 VNW pch L=4e-08 W=1.55e-07 
M16 5 CK VDD VNW pch L=4e-08 W=2.4e-07 
M17 VDD CK 5 VNW pch L=4e-08 W=2.4e-07 
M18 5 CK VDD VNW pch L=4e-08 W=2.4e-07 
M19 VDD CK 5 VNW pch L=4e-08 W=2.4e-07 
M20 5 4 VDD VNW pch L=4e-08 W=1.2e-07 
M21 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M22 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M24 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M26 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
M28 ECK 5 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 5 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X0P5B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT INV_X0P5M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=1.55e-07 
M1 Y A VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT INV_X0P6B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=1.35e-07 
M1 Y A VDD VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT INV_X0P6M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=1.85e-07 
M1 Y A VDD VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT INV_X0P7B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=1.6e-07 
M1 Y A VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT INV_X0P7M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.2e-07 
M1 Y A VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT INV_X0P8B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=1.9e-07 
M1 Y A VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT INV_X0P8M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.6e-07 
M1 Y A VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT INV_X11B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M5 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M6 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M7 Y A VDD VNW pch L=4e-08 W=4e-07 
M8 VDD A Y VNW pch L=4e-08 W=4e-07 
M9 Y A VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A Y VNW pch L=4e-08 W=4e-07 
M11 Y A VDD VNW pch L=4e-08 W=4e-07 
M12 VDD A Y VNW pch L=4e-08 W=4e-07 
M13 Y A VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A Y VNW pch L=4e-08 W=4e-07 
M15 Y A VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A Y VNW pch L=4e-08 W=4e-07 
M17 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X11M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.8e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.8e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.8e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.8e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.8e-07 
M5 VSS A Y VPW nch L=4e-08 W=3.8e-07 
M6 Y A VSS VPW nch L=4e-08 W=3.8e-07 
M7 VSS A Y VPW nch L=4e-08 W=3.8e-07 
M8 Y A VSS VPW nch L=4e-08 W=3.8e-07 
M9 Y A VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A Y VNW pch L=4e-08 W=4e-07 
M11 Y A VDD VNW pch L=4e-08 W=4e-07 
M12 VDD A Y VNW pch L=4e-08 W=4e-07 
M13 Y A VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A Y VNW pch L=4e-08 W=4e-07 
M15 Y A VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A Y VNW pch L=4e-08 W=4e-07 
M17 Y A VDD VNW pch L=4e-08 W=4e-07 
M18 VDD A Y VNW pch L=4e-08 W=4e-07 
M19 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X13B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.65e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.65e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.65e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.65e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.65e-07 
M5 VSS A Y VPW nch L=4e-08 W=3.65e-07 
M6 Y A VSS VPW nch L=4e-08 W=3.65e-07 
M7 VSS A Y VPW nch L=4e-08 W=3.65e-07 
M8 Y A VDD VNW pch L=4e-08 W=4e-07 
M9 VDD A Y VNW pch L=4e-08 W=4e-07 
M10 Y A VDD VNW pch L=4e-08 W=4e-07 
M11 VDD A Y VNW pch L=4e-08 W=4e-07 
M12 Y A VDD VNW pch L=4e-08 W=4e-07 
M13 VDD A Y VNW pch L=4e-08 W=4e-07 
M14 Y A VDD VNW pch L=4e-08 W=4e-07 
M15 VDD A Y VNW pch L=4e-08 W=4e-07 
M16 Y A VDD VNW pch L=4e-08 W=4e-07 
M17 VDD A Y VNW pch L=4e-08 W=4e-07 
M18 Y A VDD VNW pch L=4e-08 W=4e-07 
M19 VDD A Y VNW pch L=4e-08 W=4e-07 
M20 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X13M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.5e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.5e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.5e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.5e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.5e-07 
M5 VSS A Y VPW nch L=4e-08 W=3.5e-07 
M6 Y A VSS VPW nch L=4e-08 W=3.5e-07 
M7 VSS A Y VPW nch L=4e-08 W=3.5e-07 
M8 Y A VSS VPW nch L=4e-08 W=3.5e-07 
M9 VSS A Y VPW nch L=4e-08 W=3.5e-07 
M10 Y A VSS VPW nch L=4e-08 W=3.5e-07 
M11 VSS A Y VPW nch L=4e-08 W=3.5e-07 
M12 Y A VDD VNW pch L=4e-08 W=4e-07 
M13 VDD A Y VNW pch L=4e-08 W=4e-07 
M14 Y A VDD VNW pch L=4e-08 W=4e-07 
M15 VDD A Y VNW pch L=4e-08 W=4e-07 
M16 Y A VDD VNW pch L=4e-08 W=4e-07 
M17 VDD A Y VNW pch L=4e-08 W=4e-07 
M18 Y A VDD VNW pch L=4e-08 W=4e-07 
M19 VDD A Y VNW pch L=4e-08 W=4e-07 
M20 Y A VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A Y VNW pch L=4e-08 W=4e-07 
M22 Y A VDD VNW pch L=4e-08 W=4e-07 
M23 VDD A Y VNW pch L=4e-08 W=4e-07 
M24 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X16B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.6e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.6e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.6e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.6e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.6e-07 
M5 VSS A Y VPW nch L=4e-08 W=3.6e-07 
M6 Y A VSS VPW nch L=4e-08 W=3.6e-07 
M7 VSS A Y VPW nch L=4e-08 W=3.6e-07 
M8 Y A VSS VPW nch L=4e-08 W=3.6e-07 
M9 VSS A Y VPW nch L=4e-08 W=3.6e-07 
M10 Y A VDD VNW pch L=4e-08 W=4e-07 
M11 VDD A Y VNW pch L=4e-08 W=4e-07 
M12 Y A VDD VNW pch L=4e-08 W=4e-07 
M13 VDD A Y VNW pch L=4e-08 W=4e-07 
M14 Y A VDD VNW pch L=4e-08 W=4e-07 
M15 VDD A Y VNW pch L=4e-08 W=4e-07 
M16 Y A VDD VNW pch L=4e-08 W=4e-07 
M17 VDD A Y VNW pch L=4e-08 W=4e-07 
M18 Y A VDD VNW pch L=4e-08 W=4e-07 
M19 VDD A Y VNW pch L=4e-08 W=4e-07 
M20 Y A VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A Y VNW pch L=4e-08 W=4e-07 
M22 Y A VDD VNW pch L=4e-08 W=4e-07 
M23 VDD A Y VNW pch L=4e-08 W=4e-07 
M24 Y A VDD VNW pch L=4e-08 W=4e-07 
M25 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X16M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M5 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M6 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M7 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M8 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M9 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M10 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M11 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M12 Y A VSS VPW nch L=4e-08 W=3.55e-07 
M13 VSS A Y VPW nch L=4e-08 W=3.55e-07 
M14 Y A VDD VNW pch L=4e-08 W=4e-07 
M15 VDD A Y VNW pch L=4e-08 W=4e-07 
M16 Y A VDD VNW pch L=4e-08 W=4e-07 
M17 VDD A Y VNW pch L=4e-08 W=4e-07 
M18 Y A VDD VNW pch L=4e-08 W=4e-07 
M19 VDD A Y VNW pch L=4e-08 W=4e-07 
M20 Y A VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A Y VNW pch L=4e-08 W=4e-07 
M22 Y A VDD VNW pch L=4e-08 W=4e-07 
M23 VDD A Y VNW pch L=4e-08 W=4e-07 
M24 Y A VDD VNW pch L=4e-08 W=4e-07 
M25 VDD A Y VNW pch L=4e-08 W=4e-07 
M26 Y A VDD VNW pch L=4e-08 W=4e-07 
M27 VDD A Y VNW pch L=4e-08 W=4e-07 
M28 Y A VDD VNW pch L=4e-08 W=4e-07 
M29 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X1B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.25e-07 
M1 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X1M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.1e-07 
M1 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X1P2B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.7e-07 
M1 Y A VDD VNW pch L=4e-08 W=2.4e-07 
M2 VDD A Y VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT INV_X1P2M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.7e-07 
M1 Y A VDD VNW pch L=4e-08 W=2.4e-07 
M2 VDD A Y VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT INV_X1P4B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M1 Y A VDD VNW pch L=4e-08 W=2.85e-07 
M2 VDD A Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT INV_X1P4M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.2e-07 
M2 Y A VDD VNW pch L=4e-08 W=2.85e-07 
M3 VDD A Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT INV_X1P7B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.8e-07 
M1 Y A VDD VNW pch L=4e-08 W=3.35e-07 
M2 VDD A Y VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT INV_X1P7M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.6e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.6e-07 
M2 Y A VDD VNW pch L=4e-08 W=3.35e-07 
M3 VDD A Y VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT INV_X2B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.25e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.25e-07 
M2 Y A VDD VNW pch L=4e-08 W=4e-07 
M3 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X2M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.1e-07 
M2 Y A VDD VNW pch L=4e-08 W=4e-07 
M3 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X2P5B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M2 Y A VDD VNW pch L=4e-08 W=3.35e-07 
M3 VDD A Y VNW pch L=4e-08 W=3.35e-07 
M4 Y A VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT INV_X2P5M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.9e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.9e-07 
M2 Y A VDD VNW pch L=4e-08 W=3.35e-07 
M3 VDD A Y VNW pch L=4e-08 W=3.35e-07 
M4 Y A VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT INV_X3B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.4e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.4e-07 
M2 Y A VDD VNW pch L=4e-08 W=4e-07 
M3 VDD A Y VNW pch L=4e-08 W=4e-07 
M4 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X3M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.1e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.1e-07 
M3 Y A VDD VNW pch L=4e-08 W=4e-07 
M4 VDD A Y VNW pch L=4e-08 W=4e-07 
M5 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X3P5B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=4e-07 
M1 VSS A Y VPW nch L=4e-08 W=4e-07 
M2 Y A VDD VNW pch L=4e-08 W=3.5e-07 
M3 VDD A Y VNW pch L=4e-08 W=3.5e-07 
M4 Y A VDD VNW pch L=4e-08 W=3.5e-07 
M5 VDD A Y VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT INV_X3P5M_A9TR Y VDD VNW VPW VSS A
M0 VSS A Y VPW nch L=4e-08 W=3.6e-07 
M1 Y A VSS VPW nch L=4e-08 W=3.6e-07 
M2 VSS A Y VPW nch L=4e-08 W=3.6e-07 
M3 Y A VDD VNW pch L=4e-08 W=3.5e-07 
M4 VDD A Y VNW pch L=4e-08 W=3.5e-07 
M5 Y A VDD VNW pch L=4e-08 W=3.5e-07 
M6 VDD A Y VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT INV_X4B_A9TR Y VDD VNW VPW VSS A
M0 VSS A Y VPW nch L=4e-08 W=3e-07 
M1 Y A VSS VPW nch L=4e-08 W=3e-07 
M2 VSS A Y VPW nch L=4e-08 W=3e-07 
M3 Y A VDD VNW pch L=4e-08 W=4e-07 
M4 VDD A Y VNW pch L=4e-08 W=4e-07 
M5 Y A VDD VNW pch L=4e-08 W=4e-07 
M6 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X4M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.1e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.1e-07 
M4 Y A VDD VNW pch L=4e-08 W=4e-07 
M5 VDD A Y VNW pch L=4e-08 W=4e-07 
M6 Y A VDD VNW pch L=4e-08 W=4e-07 
M7 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X5B_A9TR Y VDD VNW VPW VSS A
M0 VSS A Y VPW nch L=4e-08 W=3.75e-07 
M1 Y A VSS VPW nch L=4e-08 W=3.75e-07 
M2 VSS A Y VPW nch L=4e-08 W=3.75e-07 
M3 Y A VDD VNW pch L=4e-08 W=4e-07 
M4 VDD A Y VNW pch L=4e-08 W=4e-07 
M5 Y A VDD VNW pch L=4e-08 W=4e-07 
M6 VDD A Y VNW pch L=4e-08 W=4e-07 
M7 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X5M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.9e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.9e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.9e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.9e-07 
M4 Y A VDD VNW pch L=4e-08 W=4e-07 
M5 VDD A Y VNW pch L=4e-08 W=4e-07 
M6 Y A VDD VNW pch L=4e-08 W=4e-07 
M7 VDD A Y VNW pch L=4e-08 W=4e-07 
M8 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X6B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=3.35e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.35e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.35e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.35e-07 
M4 Y A VDD VNW pch L=4e-08 W=4e-07 
M5 VDD A Y VNW pch L=4e-08 W=4e-07 
M6 Y A VDD VNW pch L=4e-08 W=4e-07 
M7 VDD A Y VNW pch L=4e-08 W=4e-07 
M8 Y A VDD VNW pch L=4e-08 W=4e-07 
M9 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X6M_A9TR Y VDD VNW VPW VSS A
M0 VSS A Y VPW nch L=4e-08 W=3.7e-07 
M1 Y A VSS VPW nch L=4e-08 W=3.7e-07 
M2 VSS A Y VPW nch L=4e-08 W=3.7e-07 
M3 Y A VSS VPW nch L=4e-08 W=3.7e-07 
M4 VSS A Y VPW nch L=4e-08 W=3.7e-07 
M5 Y A VDD VNW pch L=4e-08 W=4e-07 
M6 VDD A Y VNW pch L=4e-08 W=4e-07 
M7 Y A VDD VNW pch L=4e-08 W=4e-07 
M8 VDD A Y VNW pch L=4e-08 W=4e-07 
M9 Y A VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X7P5B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M3 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M4 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M5 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M6 Y A VDD VNW pch L=4e-08 W=3.75e-07 
M7 VDD A Y VNW pch L=4e-08 W=3.75e-07 
M8 Y A VDD VNW pch L=4e-08 W=3.75e-07 
M9 VDD A Y VNW pch L=4e-08 W=3.75e-07 
M10 Y A VDD VNW pch L=4e-08 W=3.75e-07 
M11 VDD A Y VNW pch L=4e-08 W=3.75e-07 
M12 Y A VDD VNW pch L=4e-08 W=3.75e-07 
M13 VDD A Y VNW pch L=4e-08 W=3.75e-07 
.ENDS


.SUBCKT INV_X7P5M_A9TR Y VDD VNW VPW VSS A
M0 VSS A Y VPW nch L=4e-08 W=3.3e-07 
M1 Y A VSS VPW nch L=4e-08 W=3.3e-07 
M2 VSS A Y VPW nch L=4e-08 W=3.3e-07 
M3 Y A VSS VPW nch L=4e-08 W=3.3e-07 
M4 VSS A Y VPW nch L=4e-08 W=3.3e-07 
M5 Y A VSS VPW nch L=4e-08 W=3.3e-07 
M6 VSS A Y VPW nch L=4e-08 W=3.3e-07 
M7 Y A VDD VNW pch L=4e-08 W=3.75e-07 
M8 VDD A Y VNW pch L=4e-08 W=3.75e-07 
M9 Y A VDD VNW pch L=4e-08 W=3.75e-07 
M10 VDD A Y VNW pch L=4e-08 W=3.75e-07 
M11 Y A VDD VNW pch L=4e-08 W=3.75e-07 
M12 VDD A Y VNW pch L=4e-08 W=3.75e-07 
M13 Y A VDD VNW pch L=4e-08 W=3.75e-07 
M14 VDD A Y VNW pch L=4e-08 W=3.75e-07 
.ENDS


.SUBCKT INV_X9B_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=2.9e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.9e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.9e-07 
M3 VSS A Y VPW nch L=4e-08 W=2.9e-07 
M4 Y A VSS VPW nch L=4e-08 W=2.9e-07 
M5 VSS A Y VPW nch L=4e-08 W=2.9e-07 
M6 Y A VSS VPW nch L=4e-08 W=2.9e-07 
M7 Y A VDD VNW pch L=4e-08 W=4e-07 
M8 VDD A Y VNW pch L=4e-08 W=4e-07 
M9 Y A VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A Y VNW pch L=4e-08 W=4e-07 
M11 Y A VDD VNW pch L=4e-08 W=4e-07 
M12 VDD A Y VNW pch L=4e-08 W=4e-07 
M13 Y A VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A Y VNW pch L=4e-08 W=4e-07 
M15 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT INV_X9M_A9TR Y VDD VNW VPW VSS A
M0 Y A VSS VPW nch L=4e-08 W=4e-07 
M1 VSS A Y VPW nch L=4e-08 W=4e-07 
M2 Y A VSS VPW nch L=4e-08 W=4e-07 
M3 VSS A Y VPW nch L=4e-08 W=4e-07 
M4 Y A VSS VPW nch L=4e-08 W=4e-07 
M5 VSS A Y VPW nch L=4e-08 W=4e-07 
M6 Y A VSS VPW nch L=4e-08 W=4e-07 
M7 Y A VDD VNW pch L=4e-08 W=4e-07 
M8 VDD A Y VNW pch L=4e-08 W=4e-07 
M9 Y A VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A Y VNW pch L=4e-08 W=4e-07 
M11 Y A VDD VNW pch L=4e-08 W=4e-07 
M12 VDD A Y VNW pch L=4e-08 W=4e-07 
M13 Y A VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A Y VNW pch L=4e-08 W=4e-07 
M15 Y A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATNQN_X0P5M_A9TR QN VDD VNW VPW VSS D GN
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.2e-07 
M3 11 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 QN 6 VSS VPW nch L=4e-08 W=1.55e-07 
M7 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M8 4 D VDD VNW pch L=4e-08 W=1.55e-07 
M9 5 GN 4 VNW pch L=4e-08 W=1.2e-07 
M10 10 1 5 VNW pch L=4e-08 W=1.2e-07 
M11 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M13 QN 6 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATNQN_X1M_A9TR QN VDD VNW VPW VSS D GN
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.6e-07 
M3 11 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.9e-07 
M6 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M8 4 D VDD VNW pch L=4e-08 W=2.15e-07 
M9 5 GN 4 VNW pch L=4e-08 W=1.6e-07 
M10 10 1 5 VNW pch L=4e-08 W=1.2e-07 
M11 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 5 6 VNW pch L=4e-08 W=2.25e-07 
M13 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNQN_X2M_A9TR QN VDD VNW VPW VSS D GN
M0 VSS GN 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.5e-07 
M3 11 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 7 11 VPW nch L=4e-08 W=1.2e-07 
M5 QN 7 VSS VPW nch L=4e-08 W=3.05e-07 
M6 VSS 7 QN VPW nch L=4e-08 W=3.05e-07 
M7 7 5 VSS VPW nch L=4e-08 W=3e-07 
M8 VDD GN 1 VNW pch L=4e-08 W=1.8e-07 
M9 4 D VDD VNW pch L=4e-08 W=3.45e-07 
M10 5 GN 4 VNW pch L=4e-08 W=2.5e-07 
M11 10 1 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 7 10 VNW pch L=4e-08 W=1.2e-07 
M13 QN 7 VDD VNW pch L=4e-08 W=3.75e-07 
M14 VDD 7 QN VNW pch L=4e-08 W=3.75e-07 
M15 7 5 VDD VNW pch L=4e-08 W=3.3e-07 
.ENDS


.SUBCKT LATNQN_X3M_A9TR QN VDD VNW VPW VSS D GN
M0 VSS GN 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.9e-07 
M3 11 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=3.1e-07 
M6 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M8 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VDD GN 1 VNW pch L=4e-08 W=1.9e-07 
M10 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M11 5 GN 4 VNW pch L=4e-08 W=2.9e-07 
M12 10 1 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 5 6 VNW pch L=4e-08 W=4e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 6 QN VNW pch L=4e-08 W=4e-07 
M17 QN 6 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATNQN_X4M_A9TR QN VDD VNW VPW VSS D GN
M0 VSS GN 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.9e-07 
M3 11 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=2.9e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=2.9e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 VDD GN 1 VNW pch L=4e-08 W=1.9e-07 
M12 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M13 5 GN 4 VNW pch L=4e-08 W=2.9e-07 
M14 10 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=3.4e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=3.4e-07 
M18 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M19 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
M20 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNQ_X0P5M_A9TR Q VDD VNW VPW VSS D GN
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.2e-07 
M3 11 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 Q 5 VSS VPW nch L=4e-08 W=1.55e-07 
M7 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M8 4 D VDD VNW pch L=4e-08 W=1.8e-07 
M9 5 GN 4 VNW pch L=4e-08 W=1.2e-07 
M10 10 1 5 VNW pch L=4e-08 W=1.2e-07 
M11 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M13 Q 5 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATNQ_X1M_A9TR Q VDD VNW VPW VSS D GN
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.6e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.6e-07 
M3 11 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M8 4 D VDD VNW pch L=4e-08 W=2.3e-07 
M9 5 GN 4 VNW pch L=4e-08 W=1.6e-07 
M10 10 1 5 VNW pch L=4e-08 W=1.2e-07 
M11 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M13 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNQ_X2M_A9TR Q VDD VNW VPW VSS D GN
M0 VSS GN 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.5e-07 
M3 11 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M8 VDD GN 1 VNW pch L=4e-08 W=1.7e-07 
M9 4 D VDD VNW pch L=4e-08 W=3.35e-07 
M10 5 GN 4 VNW pch L=4e-08 W=2.5e-07 
M11 10 1 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M14 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
M15 VDD 5 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNQ_X3M_A9TR Q VDD VNW VPW VSS D GN
M0 VSS GN 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.9e-07 
M3 11 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VDD GN 1 VNW pch L=4e-08 W=1.9e-07 
M10 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M11 5 GN 4 VNW pch L=4e-08 W=2.9e-07 
M12 10 1 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M15 Q 5 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 5 Q VNW pch L=4e-08 W=4e-07 
M17 Q 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATNRPQN_X0P5M_A9TR QN VDD VNW VPW VSS D GN R
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.2e-07 
M3 13 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS R 6 VPW nch L=4e-08 W=1.2e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=1.55e-07 
M8 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M9 4 D VDD VNW pch L=4e-08 W=1.55e-07 
M10 5 GN 4 VNW pch L=4e-08 W=1.2e-07 
M11 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M13 12 5 6 VNW pch L=4e-08 W=2.9e-07 
M14 VDD R 12 VNW pch L=4e-08 W=2.9e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATNRPQN_X1M_A9TR QN VDD VNW VPW VSS D GN R
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.6e-07 
M3 13 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=1.3e-07 
M6 VSS R 6 VPW nch L=4e-08 W=1.3e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M9 4 D VDD VNW pch L=4e-08 W=2.15e-07 
M10 5 GN 4 VNW pch L=4e-08 W=1.6e-07 
M11 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M13 12 5 6 VNW pch L=4e-08 W=3.1e-07 
M14 VDD R 12 VNW pch L=4e-08 W=3.1e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNRPQN_X2M_A9TR QN VDD VNW VPW VSS D GN R
M0 VSS GN 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.5e-07 
M3 13 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=1.6e-07 
M6 VSS R 6 VPW nch L=4e-08 W=1.6e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M9 VDD GN 1 VNW pch L=4e-08 W=1.8e-07 
M10 4 D VDD VNW pch L=4e-08 W=3.45e-07 
M11 5 GN 4 VNW pch L=4e-08 W=2.5e-07 
M12 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M14 12 5 6 VNW pch L=4e-08 W=4e-07 
M15 VDD R 12 VNW pch L=4e-08 W=4e-07 
M16 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M17 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNRPQN_X3M_A9TR QN VDD VNW VPW VSS D GN R
M0 VSS GN 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.9e-07 
M3 13 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=1.6e-07 
M6 VSS R 6 VPW nch L=4e-08 W=1.6e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VDD GN 1 VNW pch L=4e-08 W=1.9e-07 
M11 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M12 5 GN 4 VNW pch L=4e-08 W=2.9e-07 
M13 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M15 12 5 6 VNW pch L=4e-08 W=4e-07 
M16 VDD R 12 VNW pch L=4e-08 W=4e-07 
M17 QN 6 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 6 QN VNW pch L=4e-08 W=4e-07 
M19 QN 6 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATNRPQN_X4M_A9TR QN VDD VNW VPW VSS D GN R
M0 VSS GN 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.9e-07 
M3 14 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 6 R VSS VPW nch L=4e-08 W=1.5e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.5e-07 
M7 6 5 VSS VPW nch L=4e-08 W=1.5e-07 
M8 VSS R 6 VPW nch L=4e-08 W=1.5e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M13 VDD GN 1 VNW pch L=4e-08 W=1.9e-07 
M14 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M15 5 GN 4 VNW pch L=4e-08 W=2.9e-07 
M16 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M18 12 R VDD VNW pch L=4e-08 W=3.8e-07 
M19 6 5 12 VNW pch L=4e-08 W=3.8e-07 
M20 13 5 6 VNW pch L=4e-08 W=3.8e-07 
M21 VDD R 13 VNW pch L=4e-08 W=3.8e-07 
M22 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M23 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
M24 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNRQ_X0P5M_A9TR Q VDD VNW VPW VSS D GN RN
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 12 RN VSS VPW nch L=4e-08 W=1.4e-07 
M2 4 D 12 VPW nch L=4e-08 W=1.4e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.2e-07 
M4 13 GN 5 VPW nch L=4e-08 W=1.6e-07 
M5 14 6 13 VPW nch L=4e-08 W=1.6e-07 
M6 VSS RN 14 VPW nch L=4e-08 W=1.6e-07 
M7 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=1.55e-07 
M9 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M10 4 D VDD VNW pch L=4e-08 W=1.8e-07 
M11 5 GN 4 VNW pch L=4e-08 W=1.2e-07 
M12 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M14 5 RN VDD VNW pch L=4e-08 W=1.2e-07 
M15 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M16 Q 5 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATNRQ_X1M_A9TR Q VDD VNW VPW VSS D GN RN
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 12 RN VSS VPW nch L=4e-08 W=2e-07 
M2 4 D 12 VPW nch L=4e-08 W=2e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.6e-07 
M4 13 GN 5 VPW nch L=4e-08 W=1.6e-07 
M5 14 6 13 VPW nch L=4e-08 W=1.6e-07 
M6 VSS RN 14 VPW nch L=4e-08 W=1.6e-07 
M7 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M10 4 D VDD VNW pch L=4e-08 W=2.3e-07 
M11 5 GN 4 VNW pch L=4e-08 W=1.6e-07 
M12 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M14 5 RN VDD VNW pch L=4e-08 W=1.2e-07 
M15 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M16 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNRQ_X2M_A9TR Q VDD VNW VPW VSS D GN RN
M0 VSS GN 1 VPW nch L=4e-08 W=1.3e-07 
M1 12 RN VSS VPW nch L=4e-08 W=2.7e-07 
M2 4 D 12 VPW nch L=4e-08 W=2.7e-07 
M3 5 1 4 VPW nch L=4e-08 W=2.5e-07 
M4 13 GN 5 VPW nch L=4e-08 W=1.6e-07 
M5 14 6 13 VPW nch L=4e-08 W=1.6e-07 
M6 VSS RN 14 VPW nch L=4e-08 W=1.6e-07 
M7 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M10 VDD GN 1 VNW pch L=4e-08 W=1.7e-07 
M11 4 D VDD VNW pch L=4e-08 W=3.35e-07 
M12 5 GN 4 VNW pch L=4e-08 W=2.5e-07 
M13 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M15 5 RN VDD VNW pch L=4e-08 W=1.2e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M17 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
M18 VDD 5 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNRQ_X3M_A9TR Q VDD VNW VPW VSS D GN RN
M0 VSS GN 1 VPW nch L=4e-08 W=1.4e-07 
M1 12 RN VSS VPW nch L=4e-08 W=2.9e-07 
M2 4 D 12 VPW nch L=4e-08 W=2.9e-07 
M3 5 1 4 VPW nch L=4e-08 W=2.9e-07 
M4 13 GN 5 VPW nch L=4e-08 W=1.6e-07 
M5 14 6 13 VPW nch L=4e-08 W=1.6e-07 
M6 VSS RN 14 VPW nch L=4e-08 W=1.6e-07 
M7 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M10 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VDD GN 1 VNW pch L=4e-08 W=1.9e-07 
M12 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M13 5 GN 4 VNW pch L=4e-08 W=2.9e-07 
M14 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M16 5 RN VDD VNW pch L=4e-08 W=1.2e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M18 Q 5 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 5 Q VNW pch L=4e-08 W=4e-07 
M20 Q 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATNSPQ_X0P5M_A9TR Q VDD VNW VPW VSS D GN S
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.2e-07 
M3 14 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 5 S VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M7 Q 5 VSS VPW nch L=4e-08 W=1.55e-07 
M8 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M9 11 S VDD VNW pch L=4e-08 W=3e-07 
M10 4 D 11 VNW pch L=4e-08 W=3e-07 
M11 5 GN 4 VNW pch L=4e-08 W=1.6e-07 
M12 12 1 5 VNW pch L=4e-08 W=1.6e-07 
M13 13 6 12 VNW pch L=4e-08 W=1.6e-07 
M14 VDD S 13 VNW pch L=4e-08 W=1.6e-07 
M15 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M16 Q 5 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATNSPQ_X1M_A9TR Q VDD VNW VPW VSS D GN S
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.4e-07 
M3 14 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 5 S VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M7 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M9 11 S VDD VNW pch L=4e-08 W=3.3e-07 
M10 4 D 11 VNW pch L=4e-08 W=3.3e-07 
M11 5 GN 4 VNW pch L=4e-08 W=1.8e-07 
M12 12 1 5 VNW pch L=4e-08 W=1.6e-07 
M13 13 6 12 VNW pch L=4e-08 W=1.6e-07 
M14 VDD S 13 VNW pch L=4e-08 W=1.6e-07 
M15 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M16 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNSPQ_X2M_A9TR Q VDD VNW VPW VSS D GN S
M0 VSS GN 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2e-07 
M2 5 1 4 VPW nch L=4e-08 W=2e-07 
M3 14 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 5 S VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M7 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M9 VDD GN 1 VNW pch L=4e-08 W=1.7e-07 
M10 11 S VDD VNW pch L=4e-08 W=3.6e-07 
M11 4 D 11 VNW pch L=4e-08 W=3.6e-07 
M12 5 GN 4 VNW pch L=4e-08 W=3e-07 
M13 12 1 5 VNW pch L=4e-08 W=1.6e-07 
M14 13 6 12 VNW pch L=4e-08 W=1.6e-07 
M15 VDD S 13 VNW pch L=4e-08 W=1.6e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M17 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
M18 VDD 5 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNSPQ_X3M_A9TR Q VDD VNW VPW VSS D GN S
M0 VSS GN 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.3e-07 
M3 14 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 5 S VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M7 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M9 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VDD GN 1 VNW pch L=4e-08 W=1.9e-07 
M11 11 S VDD VNW pch L=4e-08 W=3.8e-07 
M12 4 D 11 VNW pch L=4e-08 W=3.8e-07 
M13 5 GN 4 VNW pch L=4e-08 W=2.9e-07 
M14 12 1 5 VNW pch L=4e-08 W=1.6e-07 
M15 13 6 12 VNW pch L=4e-08 W=1.6e-07 
M16 VDD S 13 VNW pch L=4e-08 W=1.6e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M18 Q 5 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 5 Q VNW pch L=4e-08 W=4e-07 
M20 Q 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATNSQN_X0P5M_A9TR QN VDD VNW VPW VSS D GN SN
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.2e-07 
M3 12 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 5 6 VPW nch L=4e-08 W=1.6e-07 
M6 VSS SN 13 VPW nch L=4e-08 W=1.6e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=1.55e-07 
M8 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M9 4 D VDD VNW pch L=4e-08 W=1.55e-07 
M10 5 GN 4 VNW pch L=4e-08 W=1.2e-07 
M11 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M13 6 5 VDD VNW pch L=4e-08 W=1.3e-07 
M14 VDD SN 6 VNW pch L=4e-08 W=1.3e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATNSQN_X1M_A9TR QN VDD VNW VPW VSS D GN SN
M0 VSS GN 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.6e-07 
M3 12 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 5 6 VPW nch L=4e-08 W=2.4e-07 
M6 VSS SN 13 VPW nch L=4e-08 W=2.4e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VDD GN 1 VNW pch L=4e-08 W=1.55e-07 
M9 4 D VDD VNW pch L=4e-08 W=2.15e-07 
M10 5 GN 4 VNW pch L=4e-08 W=1.6e-07 
M11 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M13 6 5 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD SN 6 VNW pch L=4e-08 W=4e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNSQN_X2M_A9TR QN VDD VNW VPW VSS D GN SN
M0 VSS GN 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.5e-07 
M3 12 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 SN VSS VPW nch L=4e-08 W=1.7e-07 
M6 6 5 13 VPW nch L=4e-08 W=1.7e-07 
M7 14 5 6 VPW nch L=4e-08 W=1.7e-07 
M8 VSS SN 14 VPW nch L=4e-08 W=1.7e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 VDD GN 1 VNW pch L=4e-08 W=1.8e-07 
M12 4 D VDD VNW pch L=4e-08 W=3.45e-07 
M13 5 GN 4 VNW pch L=4e-08 W=2.5e-07 
M14 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M16 6 SN VDD VNW pch L=4e-08 W=1.45e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.45e-07 
M18 6 5 VDD VNW pch L=4e-08 W=1.45e-07 
M19 VDD SN 6 VNW pch L=4e-08 W=1.45e-07 
M20 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATNSQN_X3M_A9TR QN VDD VNW VPW VSS D GN SN
M0 VSS GN 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.9e-07 
M3 12 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 SN VSS VPW nch L=4e-08 W=2e-07 
M6 6 5 13 VPW nch L=4e-08 W=2e-07 
M7 14 5 6 VPW nch L=4e-08 W=2e-07 
M8 VSS SN 14 VPW nch L=4e-08 W=2e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VDD GN 1 VNW pch L=4e-08 W=1.9e-07 
M13 4 D VDD VNW pch L=4e-08 W=3.45e-07 
M14 5 GN 4 VNW pch L=4e-08 W=2.9e-07 
M15 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M16 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M17 6 SN VDD VNW pch L=4e-08 W=1.7e-07 
M18 VDD 5 6 VNW pch L=4e-08 W=1.7e-07 
M19 6 5 VDD VNW pch L=4e-08 W=1.7e-07 
M20 VDD SN 6 VNW pch L=4e-08 W=1.7e-07 
M21 QN 6 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 6 QN VNW pch L=4e-08 W=4e-07 
M23 QN 6 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATNSQN_X4M_A9TR QN VDD VNW VPW VSS D GN SN
M0 VSS GN 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.9e-07 
M3 12 GN 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 SN VSS VPW nch L=4e-08 W=2.85e-07 
M6 6 5 13 VPW nch L=4e-08 W=2.85e-07 
M7 14 5 6 VPW nch L=4e-08 W=2.85e-07 
M8 VSS SN 14 VPW nch L=4e-08 W=2.85e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M13 VDD GN 1 VNW pch L=4e-08 W=1.9e-07 
M14 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M15 5 GN 4 VNW pch L=4e-08 W=2.9e-07 
M16 11 1 5 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M18 6 SN VDD VNW pch L=4e-08 W=2.45e-07 
M19 VDD 5 6 VNW pch L=4e-08 W=2.45e-07 
M20 6 5 VDD VNW pch L=4e-08 W=2.45e-07 
M21 VDD SN 6 VNW pch L=4e-08 W=2.45e-07 
M22 QN 6 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 6 QN VNW pch L=4e-08 W=4e-07 
M24 QN 6 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 6 QN VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATQN_X0P5M_A9TR QN VDD VNW VPW VSS D G
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.2e-07 
M3 11 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 QN 6 VSS VPW nch L=4e-08 W=1.55e-07 
M7 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M8 4 D VDD VNW pch L=4e-08 W=1.55e-07 
M9 5 1 4 VNW pch L=4e-08 W=1.2e-07 
M10 10 G 5 VNW pch L=4e-08 W=1.2e-07 
M11 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M13 QN 6 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATQN_X1M_A9TR QN VDD VNW VPW VSS D G
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.6e-07 
M3 11 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.9e-07 
M6 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M8 4 D VDD VNW pch L=4e-08 W=2.15e-07 
M9 5 1 4 VNW pch L=4e-08 W=1.6e-07 
M10 10 G 5 VNW pch L=4e-08 W=1.2e-07 
M11 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 5 6 VNW pch L=4e-08 W=2.25e-07 
M13 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATQN_X2M_A9TR QN VDD VNW VPW VSS D G
M0 VSS G 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.5e-07 
M3 11 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=3e-07 
M6 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M8 VDD G 1 VNW pch L=4e-08 W=1.8e-07 
M9 4 D VDD VNW pch L=4e-08 W=3.45e-07 
M10 5 1 4 VNW pch L=4e-08 W=2.5e-07 
M11 10 G 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 5 6 VNW pch L=4e-08 W=3.3e-07 
M14 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M15 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATQN_X3M_A9TR QN VDD VNW VPW VSS D G
M0 VSS G 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.9e-07 
M3 11 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=3.1e-07 
M6 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M8 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VDD G 1 VNW pch L=4e-08 W=1.9e-07 
M10 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M11 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M12 10 G 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 5 6 VNW pch L=4e-08 W=4e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 6 QN VNW pch L=4e-08 W=4e-07 
M17 QN 6 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATQN_X4M_A9TR QN VDD VNW VPW VSS D G
M0 VSS G 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.9e-07 
M3 11 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=2.9e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=2.9e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 VDD G 1 VNW pch L=4e-08 W=1.9e-07 
M12 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M13 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M14 10 G 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=3.4e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=3.4e-07 
M18 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M19 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
M20 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATQ_X0P5M_A9TR Q VDD VNW VPW VSS D G
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.2e-07 
M3 11 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 Q 5 VSS VPW nch L=4e-08 W=1.55e-07 
M7 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M8 4 D VDD VNW pch L=4e-08 W=1.8e-07 
M9 5 1 4 VNW pch L=4e-08 W=1.2e-07 
M10 10 G 5 VNW pch L=4e-08 W=1.2e-07 
M11 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M13 Q 5 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATQ_X1M_A9TR Q VDD VNW VPW VSS D G
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.6e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.6e-07 
M3 11 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M8 4 D VDD VNW pch L=4e-08 W=2.3e-07 
M9 5 1 4 VNW pch L=4e-08 W=1.6e-07 
M10 10 G 5 VNW pch L=4e-08 W=1.2e-07 
M11 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M13 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATQ_X2M_A9TR Q VDD VNW VPW VSS D G
M0 VSS G 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.5e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.5e-07 
M3 11 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M8 VDD G 1 VNW pch L=4e-08 W=1.7e-07 
M9 4 D VDD VNW pch L=4e-08 W=3.35e-07 
M10 5 1 4 VNW pch L=4e-08 W=2.5e-07 
M11 10 G 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M14 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
M15 VDD 5 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATQ_X3M_A9TR Q VDD VNW VPW VSS D G
M0 VSS G 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.9e-07 
M3 11 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 11 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VDD G 1 VNW pch L=4e-08 W=1.9e-07 
M10 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M11 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M12 10 G 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 10 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M15 Q 5 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 5 Q VNW pch L=4e-08 W=4e-07 
M17 Q 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATRPQN_X0P5M_A9TR QN VDD VNW VPW VSS D G R
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.2e-07 
M3 13 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS R 6 VPW nch L=4e-08 W=1.2e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=1.55e-07 
M8 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M9 4 D VDD VNW pch L=4e-08 W=1.55e-07 
M10 5 1 4 VNW pch L=4e-08 W=1.2e-07 
M11 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M13 12 5 6 VNW pch L=4e-08 W=2.9e-07 
M14 VDD R 12 VNW pch L=4e-08 W=2.9e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATRPQN_X1M_A9TR QN VDD VNW VPW VSS D G R
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.6e-07 
M3 13 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=1.3e-07 
M6 VSS R 6 VPW nch L=4e-08 W=1.3e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M9 4 D VDD VNW pch L=4e-08 W=2.15e-07 
M10 5 1 4 VNW pch L=4e-08 W=1.6e-07 
M11 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M13 12 5 6 VNW pch L=4e-08 W=3.1e-07 
M14 VDD R 12 VNW pch L=4e-08 W=3.1e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATRPQN_X2M_A9TR QN VDD VNW VPW VSS D G R
M0 VSS G 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.5e-07 
M3 13 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=1.6e-07 
M6 VSS R 6 VPW nch L=4e-08 W=1.6e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M9 VDD G 1 VNW pch L=4e-08 W=1.8e-07 
M10 4 D VDD VNW pch L=4e-08 W=3.45e-07 
M11 5 1 4 VNW pch L=4e-08 W=2.5e-07 
M12 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M14 12 5 6 VNW pch L=4e-08 W=4e-07 
M15 VDD R 12 VNW pch L=4e-08 W=4e-07 
M16 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M17 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATRPQN_X3M_A9TR QN VDD VNW VPW VSS D G R
M0 VSS G 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.9e-07 
M3 13 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 6 5 VSS VPW nch L=4e-08 W=1.6e-07 
M6 VSS R 6 VPW nch L=4e-08 W=1.6e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VDD G 1 VNW pch L=4e-08 W=1.9e-07 
M11 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M12 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M13 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M15 12 5 6 VNW pch L=4e-08 W=4e-07 
M16 VDD R 12 VNW pch L=4e-08 W=4e-07 
M17 QN 6 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 6 QN VNW pch L=4e-08 W=4e-07 
M19 QN 6 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATRPQN_X4M_A9TR QN VDD VNW VPW VSS D G R
M0 VSS G 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.9e-07 
M3 14 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 6 R VSS VPW nch L=4e-08 W=1.5e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.5e-07 
M7 6 5 VSS VPW nch L=4e-08 W=1.5e-07 
M8 VSS R 6 VPW nch L=4e-08 W=1.5e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M13 VDD G 1 VNW pch L=4e-08 W=1.9e-07 
M14 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M15 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M16 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M18 12 R VDD VNW pch L=4e-08 W=3.8e-07 
M19 6 5 12 VNW pch L=4e-08 W=3.8e-07 
M20 13 5 6 VNW pch L=4e-08 W=3.8e-07 
M21 VDD R 13 VNW pch L=4e-08 W=3.8e-07 
M22 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M23 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
M24 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATRQ_X0P5M_A9TR Q VDD VNW VPW VSS D G RN
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 12 RN VSS VPW nch L=4e-08 W=1.4e-07 
M2 4 D 12 VPW nch L=4e-08 W=1.4e-07 
M3 5 G 4 VPW nch L=4e-08 W=1.2e-07 
M4 13 1 5 VPW nch L=4e-08 W=1.6e-07 
M5 14 6 13 VPW nch L=4e-08 W=1.6e-07 
M6 VSS RN 14 VPW nch L=4e-08 W=1.6e-07 
M7 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=1.55e-07 
M9 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M10 4 D VDD VNW pch L=4e-08 W=1.8e-07 
M11 5 1 4 VNW pch L=4e-08 W=1.2e-07 
M12 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M14 5 RN VDD VNW pch L=4e-08 W=1.2e-07 
M15 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M16 Q 5 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATRQ_X1M_A9TR Q VDD VNW VPW VSS D G RN
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 12 RN VSS VPW nch L=4e-08 W=2e-07 
M2 4 D 12 VPW nch L=4e-08 W=2e-07 
M3 5 G 4 VPW nch L=4e-08 W=1.6e-07 
M4 13 1 5 VPW nch L=4e-08 W=1.6e-07 
M5 14 6 13 VPW nch L=4e-08 W=1.6e-07 
M6 VSS RN 14 VPW nch L=4e-08 W=1.6e-07 
M7 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M10 4 D VDD VNW pch L=4e-08 W=2.3e-07 
M11 5 1 4 VNW pch L=4e-08 W=1.6e-07 
M12 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M14 5 RN VDD VNW pch L=4e-08 W=1.2e-07 
M15 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M16 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATRQ_X2M_A9TR Q VDD VNW VPW VSS D G RN
M0 VSS G 1 VPW nch L=4e-08 W=1.3e-07 
M1 12 RN VSS VPW nch L=4e-08 W=2.7e-07 
M2 4 D 12 VPW nch L=4e-08 W=2.7e-07 
M3 5 G 4 VPW nch L=4e-08 W=2.5e-07 
M4 13 1 5 VPW nch L=4e-08 W=1.6e-07 
M5 14 6 13 VPW nch L=4e-08 W=1.6e-07 
M6 VSS RN 14 VPW nch L=4e-08 W=1.6e-07 
M7 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M10 VDD G 1 VNW pch L=4e-08 W=1.7e-07 
M11 4 D VDD VNW pch L=4e-08 W=3.35e-07 
M12 5 1 4 VNW pch L=4e-08 W=2.5e-07 
M13 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M15 5 RN VDD VNW pch L=4e-08 W=1.2e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M17 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
M18 VDD 5 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATRQ_X3M_A9TR Q VDD VNW VPW VSS D G RN
M0 VSS G 1 VPW nch L=4e-08 W=1.4e-07 
M1 12 RN VSS VPW nch L=4e-08 W=2.9e-07 
M2 4 D 12 VPW nch L=4e-08 W=2.9e-07 
M3 5 G 4 VPW nch L=4e-08 W=2.9e-07 
M4 13 1 5 VPW nch L=4e-08 W=1.6e-07 
M5 14 6 13 VPW nch L=4e-08 W=1.6e-07 
M6 VSS RN 14 VPW nch L=4e-08 W=1.6e-07 
M7 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M8 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M10 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VDD G 1 VNW pch L=4e-08 W=1.9e-07 
M12 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M13 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M14 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M16 5 RN VDD VNW pch L=4e-08 W=1.2e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M18 Q 5 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 5 Q VNW pch L=4e-08 W=4e-07 
M20 Q 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATSPQ_X0P5M_A9TR Q VDD VNW VPW VSS D G S
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.2e-07 
M3 14 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 5 S VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M7 Q 5 VSS VPW nch L=4e-08 W=1.55e-07 
M8 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M9 11 S VDD VNW pch L=4e-08 W=3e-07 
M10 4 D 11 VNW pch L=4e-08 W=3e-07 
M11 5 1 4 VNW pch L=4e-08 W=1.6e-07 
M12 12 G 5 VNW pch L=4e-08 W=1.6e-07 
M13 13 6 12 VNW pch L=4e-08 W=1.6e-07 
M14 VDD S 13 VNW pch L=4e-08 W=1.6e-07 
M15 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M16 Q 5 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATSPQ_X1M_A9TR Q VDD VNW VPW VSS D G S
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.4e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.4e-07 
M3 14 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 5 S VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M7 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M9 11 S VDD VNW pch L=4e-08 W=3.3e-07 
M10 4 D 11 VNW pch L=4e-08 W=3.3e-07 
M11 5 1 4 VNW pch L=4e-08 W=1.8e-07 
M12 12 G 5 VNW pch L=4e-08 W=1.6e-07 
M13 13 6 12 VNW pch L=4e-08 W=1.6e-07 
M14 VDD S 13 VNW pch L=4e-08 W=1.6e-07 
M15 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M16 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATSPQ_X2M_A9TR Q VDD VNW VPW VSS D G S
M0 VSS G 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2e-07 
M2 5 G 4 VPW nch L=4e-08 W=2e-07 
M3 14 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 5 S VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M7 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M9 VDD G 1 VNW pch L=4e-08 W=1.7e-07 
M10 11 S VDD VNW pch L=4e-08 W=3.6e-07 
M11 4 D 11 VNW pch L=4e-08 W=3.6e-07 
M12 5 1 4 VNW pch L=4e-08 W=3e-07 
M13 12 G 5 VNW pch L=4e-08 W=1.6e-07 
M14 13 6 12 VNW pch L=4e-08 W=1.6e-07 
M15 VDD S 13 VNW pch L=4e-08 W=1.6e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M17 Q 5 VDD VNW pch L=4e-08 W=3.8e-07 
M18 VDD 5 Q VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATSPQ_X3M_A9TR Q VDD VNW VPW VSS D G S
M0 VSS G 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.3e-07 
M3 14 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 5 S VSS VPW nch L=4e-08 W=1.2e-07 
M6 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M7 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS 5 Q VPW nch L=4e-08 W=3.1e-07 
M9 Q 5 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VDD G 1 VNW pch L=4e-08 W=1.9e-07 
M11 11 S VDD VNW pch L=4e-08 W=3.8e-07 
M12 4 D 11 VNW pch L=4e-08 W=3.8e-07 
M13 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M14 12 G 5 VNW pch L=4e-08 W=1.6e-07 
M15 13 6 12 VNW pch L=4e-08 W=1.6e-07 
M16 VDD S 13 VNW pch L=4e-08 W=1.6e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M18 Q 5 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 5 Q VNW pch L=4e-08 W=4e-07 
M20 Q 5 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATSQN_X0P5M_A9TR QN VDD VNW VPW VSS D G SN
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.2e-07 
M3 12 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 5 6 VPW nch L=4e-08 W=1.6e-07 
M6 VSS SN 13 VPW nch L=4e-08 W=1.6e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=1.55e-07 
M8 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M9 4 D VDD VNW pch L=4e-08 W=1.55e-07 
M10 5 1 4 VNW pch L=4e-08 W=1.2e-07 
M11 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M13 6 5 VDD VNW pch L=4e-08 W=1.3e-07 
M14 VDD SN 6 VNW pch L=4e-08 W=1.3e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT LATSQN_X1M_A9TR QN VDD VNW VPW VSS D G SN
M0 VSS G 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 D VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 G 4 VPW nch L=4e-08 W=1.6e-07 
M3 12 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 5 6 VPW nch L=4e-08 W=2.4e-07 
M6 VSS SN 13 VPW nch L=4e-08 W=2.4e-07 
M7 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VDD G 1 VNW pch L=4e-08 W=1.55e-07 
M9 4 D VDD VNW pch L=4e-08 W=2.15e-07 
M10 5 1 4 VNW pch L=4e-08 W=1.6e-07 
M11 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M12 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M13 6 5 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD SN 6 VNW pch L=4e-08 W=4e-07 
M15 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATSQN_X2M_A9TR QN VDD VNW VPW VSS D G SN
M0 VSS G 1 VPW nch L=4e-08 W=1.3e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.5e-07 
M3 12 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 SN VSS VPW nch L=4e-08 W=1.7e-07 
M6 6 5 13 VPW nch L=4e-08 W=1.7e-07 
M7 14 5 6 VPW nch L=4e-08 W=1.7e-07 
M8 VSS SN 14 VPW nch L=4e-08 W=1.7e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 VDD G 1 VNW pch L=4e-08 W=1.8e-07 
M12 4 D VDD VNW pch L=4e-08 W=3.45e-07 
M13 5 1 4 VNW pch L=4e-08 W=2.5e-07 
M14 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M16 6 SN VDD VNW pch L=4e-08 W=1.45e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.45e-07 
M18 6 5 VDD VNW pch L=4e-08 W=1.45e-07 
M19 VDD SN 6 VNW pch L=4e-08 W=1.45e-07 
M20 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT LATSQN_X3M_A9TR QN VDD VNW VPW VSS D G SN
M0 VSS G 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.9e-07 
M3 12 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 SN VSS VPW nch L=4e-08 W=2e-07 
M6 6 5 13 VPW nch L=4e-08 W=2e-07 
M7 14 5 6 VPW nch L=4e-08 W=2e-07 
M8 VSS SN 14 VPW nch L=4e-08 W=2e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VDD G 1 VNW pch L=4e-08 W=1.9e-07 
M13 4 D VDD VNW pch L=4e-08 W=3.45e-07 
M14 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M15 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M16 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M17 6 SN VDD VNW pch L=4e-08 W=1.7e-07 
M18 VDD 5 6 VNW pch L=4e-08 W=1.7e-07 
M19 6 5 VDD VNW pch L=4e-08 W=1.7e-07 
M20 VDD SN 6 VNW pch L=4e-08 W=1.7e-07 
M21 QN 6 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 6 QN VNW pch L=4e-08 W=4e-07 
M23 QN 6 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT LATSQN_X4M_A9TR QN VDD VNW VPW VSS D G SN
M0 VSS G 1 VPW nch L=4e-08 W=1.4e-07 
M1 4 D VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 G 4 VPW nch L=4e-08 W=2.9e-07 
M3 12 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M5 13 SN VSS VPW nch L=4e-08 W=2.85e-07 
M6 6 5 13 VPW nch L=4e-08 W=2.85e-07 
M7 14 5 6 VPW nch L=4e-08 W=2.85e-07 
M8 VSS SN 14 VPW nch L=4e-08 W=2.85e-07 
M9 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M11 QN 6 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 6 QN VPW nch L=4e-08 W=3.1e-07 
M13 VDD G 1 VNW pch L=4e-08 W=1.9e-07 
M14 4 D VDD VNW pch L=4e-08 W=3.8e-07 
M15 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M16 11 G 5 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 6 11 VNW pch L=4e-08 W=1.2e-07 
M18 6 SN VDD VNW pch L=4e-08 W=2.45e-07 
M19 VDD 5 6 VNW pch L=4e-08 W=2.45e-07 
M20 6 5 VDD VNW pch L=4e-08 W=2.45e-07 
M21 VDD SN 6 VNW pch L=4e-08 W=2.45e-07 
M22 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M23 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
M24 QN 6 VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD 6 QN VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT M2SDFFQN_X0P5M_A9TR QN VDD VNW VPW VSS CK D0 D1 S0 SE SI
M0 VSS D1 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.2e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.2e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.2e-07 
M4 VSS D0 5 VPW nch L=4e-08 W=1.2e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.2e-07 
M7 26 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=1.2e-07 
M10 10 16 9 VPW nch L=4e-08 W=1.2e-07 
M11 27 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 27 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=1.2e-07 
M14 12 15 11 VPW nch L=4e-08 W=1.2e-07 
M15 28 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 28 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 QN 13 VSS VPW nch L=4e-08 W=1.55e-07 
M19 VSS 16 15 VPW nch L=4e-08 W=1.2e-07 
M20 16 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 VDD D1 1 VNW pch L=4e-08 W=2.4e-07 
M22 4 S0 VDD VNW pch L=4e-08 W=2.2e-07 
M23 6 S0 5 VNW pch L=4e-08 W=2.2e-07 
M24 1 4 6 VNW pch L=4e-08 W=2.2e-07 
M25 VDD D0 5 VNW pch L=4e-08 W=2.4e-07 
M26 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M27 8 SE 6 VNW pch L=4e-08 W=2.2e-07 
M28 23 7 8 VNW pch L=4e-08 W=1.55e-07 
M29 VDD SI 23 VNW pch L=4e-08 W=1.55e-07 
M30 9 8 VDD VNW pch L=4e-08 W=1.3e-07 
M31 10 15 9 VNW pch L=4e-08 W=1.2e-07 
M32 24 16 10 VNW pch L=4e-08 W=1.2e-07 
M33 VDD 11 24 VNW pch L=4e-08 W=1.2e-07 
M34 11 10 VDD VNW pch L=4e-08 W=1.55e-07 
M35 12 16 11 VNW pch L=4e-08 W=1.2e-07 
M36 25 15 12 VNW pch L=4e-08 W=1.2e-07 
M37 VDD 13 25 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 12 13 VNW pch L=4e-08 W=1.55e-07 
M39 QN 13 VDD VNW pch L=4e-08 W=2e-07 
M40 VDD 16 15 VNW pch L=4e-08 W=2.5e-07 
M41 16 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT M2SDFFQN_X1M_A9TR QN VDD VNW VPW VSS CK D0 D1 S0 SE SI
M0 VSS D1 1 VPW nch L=4e-08 W=1.6e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.6e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.6e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.6e-07 
M4 VSS D0 5 VPW nch L=4e-08 W=1.6e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.6e-07 
M7 26 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=1.6e-07 
M10 10 16 9 VPW nch L=4e-08 W=1.6e-07 
M11 27 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 27 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=1.6e-07 
M14 12 15 11 VPW nch L=4e-08 W=1.6e-07 
M15 28 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 28 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.75e-07 
M18 QN 13 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 16 15 VPW nch L=4e-08 W=1.2e-07 
M20 16 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 VDD D1 1 VNW pch L=4e-08 W=3.4e-07 
M22 4 S0 VDD VNW pch L=4e-08 W=3.2e-07 
M23 6 S0 5 VNW pch L=4e-08 W=3.2e-07 
M24 1 4 6 VNW pch L=4e-08 W=3.2e-07 
M25 VDD D0 5 VNW pch L=4e-08 W=3.4e-07 
M26 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M27 8 SE 6 VNW pch L=4e-08 W=3.2e-07 
M28 23 7 8 VNW pch L=4e-08 W=1.55e-07 
M29 VDD SI 23 VNW pch L=4e-08 W=1.55e-07 
M30 9 8 VDD VNW pch L=4e-08 W=1.75e-07 
M31 10 15 9 VNW pch L=4e-08 W=1.6e-07 
M32 24 16 10 VNW pch L=4e-08 W=1.2e-07 
M33 VDD 11 24 VNW pch L=4e-08 W=1.2e-07 
M34 11 10 VDD VNW pch L=4e-08 W=2.05e-07 
M35 12 16 11 VNW pch L=4e-08 W=1.6e-07 
M36 25 15 12 VNW pch L=4e-08 W=1.2e-07 
M37 VDD 13 25 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 12 13 VNW pch L=4e-08 W=2.45e-07 
M39 QN 13 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 16 15 VNW pch L=4e-08 W=2.5e-07 
M41 16 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT M2SDFFQN_X2M_A9TR QN VDD VNW VPW VSS CK D0 D1 S0 SE SI
M0 VSS D1 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.8e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS D0 5 VPW nch L=4e-08 W=1.8e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.8e-07 
M7 26 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=2.5e-07 
M10 10 16 9 VPW nch L=4e-08 W=2.5e-07 
M11 27 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 27 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=2.5e-07 
M14 12 15 11 VPW nch L=4e-08 W=2.5e-07 
M15 28 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 28 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=2.5e-07 
M18 QN 13 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 13 QN VPW nch L=4e-08 W=3.1e-07 
M20 VSS 16 15 VPW nch L=4e-08 W=1.3e-07 
M21 16 CK VSS VPW nch L=4e-08 W=1.3e-07 
M22 VDD D1 1 VNW pch L=4e-08 W=4e-07 
M23 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M24 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M25 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M26 VDD D0 5 VNW pch L=4e-08 W=3.8e-07 
M27 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M28 8 SE 6 VNW pch L=4e-08 W=3.8e-07 
M29 23 7 8 VNW pch L=4e-08 W=1.55e-07 
M30 VDD SI 23 VNW pch L=4e-08 W=1.55e-07 
M31 9 8 VDD VNW pch L=4e-08 W=2.7e-07 
M32 10 15 9 VNW pch L=4e-08 W=2.5e-07 
M33 24 16 10 VNW pch L=4e-08 W=1.2e-07 
M34 VDD 11 24 VNW pch L=4e-08 W=1.2e-07 
M35 11 10 VDD VNW pch L=4e-08 W=3.25e-07 
M36 12 16 11 VNW pch L=4e-08 W=2.5e-07 
M37 25 15 12 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 13 25 VNW pch L=4e-08 W=1.2e-07 
M39 VDD 12 13 VNW pch L=4e-08 W=3.8e-07 
M40 QN 13 VDD VNW pch L=4e-08 W=3.8e-07 
M41 VDD 13 QN VNW pch L=4e-08 W=3.8e-07 
M42 VDD 16 15 VNW pch L=4e-08 W=2.7e-07 
M43 16 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT M2SDFFQN_X3M_A9TR QN VDD VNW VPW VSS CK D0 D1 S0 SE SI
M0 VSS D1 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.8e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS D0 5 VPW nch L=4e-08 W=1.8e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.8e-07 
M7 26 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=3.1e-07 
M10 10 16 9 VPW nch L=4e-08 W=3.1e-07 
M11 27 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 27 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=3.1e-07 
M14 12 15 11 VPW nch L=4e-08 W=3.1e-07 
M15 28 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 28 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=2.5e-07 
M18 QN 13 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 13 QN VPW nch L=4e-08 W=3.1e-07 
M20 QN 13 VSS VPW nch L=4e-08 W=3.1e-07 
M21 VSS 16 15 VPW nch L=4e-08 W=1.4e-07 
M22 16 CK VSS VPW nch L=4e-08 W=1.4e-07 
M23 VDD D1 1 VNW pch L=4e-08 W=4e-07 
M24 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M25 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M26 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M27 VDD D0 5 VNW pch L=4e-08 W=3.8e-07 
M28 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M29 8 SE 6 VNW pch L=4e-08 W=3.8e-07 
M30 23 7 8 VNW pch L=4e-08 W=1.55e-07 
M31 VDD SI 23 VNW pch L=4e-08 W=1.55e-07 
M32 9 8 VDD VNW pch L=4e-08 W=3.3e-07 
M33 10 15 9 VNW pch L=4e-08 W=3.1e-07 
M34 24 16 10 VNW pch L=4e-08 W=1.2e-07 
M35 VDD 11 24 VNW pch L=4e-08 W=1.2e-07 
M36 11 10 VDD VNW pch L=4e-08 W=3.8e-07 
M37 12 16 11 VNW pch L=4e-08 W=3.1e-07 
M38 25 15 12 VNW pch L=4e-08 W=1.2e-07 
M39 VDD 13 25 VNW pch L=4e-08 W=1.2e-07 
M40 VDD 12 13 VNW pch L=4e-08 W=3.8e-07 
M41 QN 13 VDD VNW pch L=4e-08 W=3.8e-07 
M42 VDD 13 QN VNW pch L=4e-08 W=3.8e-07 
M43 QN 13 VDD VNW pch L=4e-08 W=3.8e-07 
M44 VDD 16 15 VNW pch L=4e-08 W=2.9e-07 
M45 16 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT M2SDFFQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
M0 VSS D1 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.2e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.2e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.2e-07 
M4 VSS D0 5 VPW nch L=4e-08 W=1.2e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.2e-07 
M7 26 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=1.2e-07 
M10 10 16 9 VPW nch L=4e-08 W=1.2e-07 
M11 27 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 27 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=1.2e-07 
M14 12 15 11 VPW nch L=4e-08 W=1.2e-07 
M15 28 16 12 VPW nch L=4e-08 W=1.5e-07 
M16 VSS 13 28 VPW nch L=4e-08 W=1.5e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 Q 12 VSS VPW nch L=4e-08 W=1.55e-07 
M19 VSS 16 15 VPW nch L=4e-08 W=1.2e-07 
M20 16 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 VDD D1 1 VNW pch L=4e-08 W=2.4e-07 
M22 4 S0 VDD VNW pch L=4e-08 W=2.2e-07 
M23 6 S0 5 VNW pch L=4e-08 W=2.2e-07 
M24 1 4 6 VNW pch L=4e-08 W=2.2e-07 
M25 VDD D0 5 VNW pch L=4e-08 W=2.4e-07 
M26 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M27 8 SE 6 VNW pch L=4e-08 W=2.2e-07 
M28 23 7 8 VNW pch L=4e-08 W=1.55e-07 
M29 VDD SI 23 VNW pch L=4e-08 W=1.55e-07 
M30 9 8 VDD VNW pch L=4e-08 W=1.3e-07 
M31 10 15 9 VNW pch L=4e-08 W=1.2e-07 
M32 24 16 10 VNW pch L=4e-08 W=1.2e-07 
M33 VDD 11 24 VNW pch L=4e-08 W=1.2e-07 
M34 11 10 VDD VNW pch L=4e-08 W=1.8e-07 
M35 12 16 11 VNW pch L=4e-08 W=1.2e-07 
M36 25 15 12 VNW pch L=4e-08 W=1.5e-07 
M37 VDD 13 25 VNW pch L=4e-08 W=1.5e-07 
M38 VDD 12 13 VNW pch L=4e-08 W=1.2e-07 
M39 Q 12 VDD VNW pch L=4e-08 W=2e-07 
M40 VDD 16 15 VNW pch L=4e-08 W=2.5e-07 
M41 16 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT M2SDFFQ_X1M_A9TR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
M0 VSS D1 1 VPW nch L=4e-08 W=1.6e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.6e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.6e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.6e-07 
M4 VSS D0 5 VPW nch L=4e-08 W=1.6e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.6e-07 
M7 26 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=1.6e-07 
M10 10 16 9 VPW nch L=4e-08 W=1.6e-07 
M11 27 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 27 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=1.6e-07 
M14 12 15 11 VPW nch L=4e-08 W=1.6e-07 
M15 28 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 28 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 16 15 VPW nch L=4e-08 W=1.2e-07 
M20 16 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 VDD D1 1 VNW pch L=4e-08 W=3.4e-07 
M22 4 S0 VDD VNW pch L=4e-08 W=3.2e-07 
M23 6 S0 5 VNW pch L=4e-08 W=3.2e-07 
M24 1 4 6 VNW pch L=4e-08 W=3.2e-07 
M25 VDD D0 5 VNW pch L=4e-08 W=3.4e-07 
M26 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M27 8 SE 6 VNW pch L=4e-08 W=3.2e-07 
M28 23 7 8 VNW pch L=4e-08 W=1.55e-07 
M29 VDD SI 23 VNW pch L=4e-08 W=1.55e-07 
M30 9 8 VDD VNW pch L=4e-08 W=1.75e-07 
M31 10 15 9 VNW pch L=4e-08 W=1.6e-07 
M32 24 16 10 VNW pch L=4e-08 W=1.2e-07 
M33 VDD 11 24 VNW pch L=4e-08 W=1.2e-07 
M34 11 10 VDD VNW pch L=4e-08 W=2.3e-07 
M35 12 16 11 VNW pch L=4e-08 W=1.6e-07 
M36 25 15 12 VNW pch L=4e-08 W=1.2e-07 
M37 VDD 13 25 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 12 13 VNW pch L=4e-08 W=1.2e-07 
M39 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 16 15 VNW pch L=4e-08 W=2.5e-07 
M41 16 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT M2SDFFQ_X2M_A9TR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
M0 VSS D1 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.8e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS D0 5 VPW nch L=4e-08 W=1.8e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.8e-07 
M7 26 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=2.5e-07 
M10 10 16 9 VPW nch L=4e-08 W=2.5e-07 
M11 27 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 27 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=2.5e-07 
M14 12 15 11 VPW nch L=4e-08 W=2.5e-07 
M15 28 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 28 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 12 Q VPW nch L=4e-08 W=3.1e-07 
M20 VSS 16 15 VPW nch L=4e-08 W=1.3e-07 
M21 16 CK VSS VPW nch L=4e-08 W=1.3e-07 
M22 VDD D1 1 VNW pch L=4e-08 W=3.8e-07 
M23 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M24 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M25 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M26 VDD D0 5 VNW pch L=4e-08 W=3.8e-07 
M27 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M28 8 SE 6 VNW pch L=4e-08 W=3.8e-07 
M29 23 7 8 VNW pch L=4e-08 W=1.55e-07 
M30 VDD SI 23 VNW pch L=4e-08 W=1.55e-07 
M31 9 8 VDD VNW pch L=4e-08 W=2.7e-07 
M32 10 15 9 VNW pch L=4e-08 W=2.5e-07 
M33 24 16 10 VNW pch L=4e-08 W=1.2e-07 
M34 VDD 11 24 VNW pch L=4e-08 W=1.2e-07 
M35 11 10 VDD VNW pch L=4e-08 W=3.35e-07 
M36 12 16 11 VNW pch L=4e-08 W=2.5e-07 
M37 25 15 12 VNW pch L=4e-08 W=1.2e-07 
M38 VDD 13 25 VNW pch L=4e-08 W=1.2e-07 
M39 VDD 12 13 VNW pch L=4e-08 W=1.2e-07 
M40 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M41 VDD 12 Q VNW pch L=4e-08 W=3.8e-07 
M42 VDD 16 15 VNW pch L=4e-08 W=2.7e-07 
M43 16 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT M2SDFFQ_X3M_A9TR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
M0 VSS D1 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.8e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS D0 5 VPW nch L=4e-08 W=1.8e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.8e-07 
M7 26 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=3.1e-07 
M10 10 16 9 VPW nch L=4e-08 W=3.1e-07 
M11 27 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 27 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=3.1e-07 
M14 12 15 11 VPW nch L=4e-08 W=3.1e-07 
M15 28 16 12 VPW nch L=4e-08 W=1.2e-07 
M16 VSS 13 28 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M18 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 12 Q VPW nch L=4e-08 W=3.1e-07 
M20 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M21 VSS 16 15 VPW nch L=4e-08 W=1.4e-07 
M22 16 CK VSS VPW nch L=4e-08 W=1.4e-07 
M23 VDD D1 1 VNW pch L=4e-08 W=4e-07 
M24 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M25 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M26 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M27 VDD D0 5 VNW pch L=4e-08 W=3.8e-07 
M28 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M29 8 SE 6 VNW pch L=4e-08 W=3.8e-07 
M30 23 7 8 VNW pch L=4e-08 W=1.55e-07 
M31 VDD SI 23 VNW pch L=4e-08 W=1.55e-07 
M32 9 8 VDD VNW pch L=4e-08 W=3.3e-07 
M33 10 15 9 VNW pch L=4e-08 W=3.1e-07 
M34 24 16 10 VNW pch L=4e-08 W=1.2e-07 
M35 VDD 11 24 VNW pch L=4e-08 W=1.2e-07 
M36 11 10 VDD VNW pch L=4e-08 W=3.8e-07 
M37 12 16 11 VNW pch L=4e-08 W=3.1e-07 
M38 25 15 12 VNW pch L=4e-08 W=1.2e-07 
M39 VDD 13 25 VNW pch L=4e-08 W=1.2e-07 
M40 VDD 12 13 VNW pch L=4e-08 W=1.2e-07 
M41 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M42 VDD 12 Q VNW pch L=4e-08 W=3.8e-07 
M43 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M44 VDD 16 15 VNW pch L=4e-08 W=2.9e-07 
M45 16 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT M2SDFFQ_X4M_A9TR Q VDD VNW VPW VSS CK D0 D1 S0 SE SI
M0 VSS D1 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.8e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS D0 5 VPW nch L=4e-08 W=1.8e-07 
M5 7 SE VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 7 6 VPW nch L=4e-08 W=1.8e-07 
M7 26 SE 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M9 9 8 VSS VPW nch L=4e-08 W=3.1e-07 
M10 10 16 9 VPW nch L=4e-08 W=3.1e-07 
M11 27 15 10 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 11 27 VPW nch L=4e-08 W=1.2e-07 
M13 11 10 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 10 11 VPW nch L=4e-08 W=3.1e-07 
M15 12 15 11 VPW nch L=4e-08 W=3.1e-07 
M16 28 16 12 VPW nch L=4e-08 W=1.2e-07 
M17 VSS 13 28 VPW nch L=4e-08 W=1.2e-07 
M18 VSS 12 13 VPW nch L=4e-08 W=1.2e-07 
M19 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M20 VSS 12 Q VPW nch L=4e-08 W=3.1e-07 
M21 Q 12 VSS VPW nch L=4e-08 W=3.1e-07 
M22 VSS 12 Q VPW nch L=4e-08 W=3.1e-07 
M23 VSS 16 15 VPW nch L=4e-08 W=1.4e-07 
M24 16 CK VSS VPW nch L=4e-08 W=1.4e-07 
M25 VDD D1 1 VNW pch L=4e-08 W=4e-07 
M26 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M27 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M28 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M29 VDD D0 5 VNW pch L=4e-08 W=3.8e-07 
M30 7 SE VDD VNW pch L=4e-08 W=1.7e-07 
M31 8 SE 6 VNW pch L=4e-08 W=3.8e-07 
M32 23 7 8 VNW pch L=4e-08 W=1.55e-07 
M33 VDD SI 23 VNW pch L=4e-08 W=1.55e-07 
M34 9 8 VDD VNW pch L=4e-08 W=3.3e-07 
M35 10 15 9 VNW pch L=4e-08 W=3.1e-07 
M36 24 16 10 VNW pch L=4e-08 W=1.2e-07 
M37 VDD 11 24 VNW pch L=4e-08 W=1.2e-07 
M38 11 10 VDD VNW pch L=4e-08 W=3.8e-07 
M39 VDD 10 11 VNW pch L=4e-08 W=3.8e-07 
M40 12 16 11 VNW pch L=4e-08 W=3.1e-07 
M41 25 15 12 VNW pch L=4e-08 W=1.2e-07 
M42 VDD 13 25 VNW pch L=4e-08 W=1.2e-07 
M43 VDD 12 13 VNW pch L=4e-08 W=1.2e-07 
M44 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M45 VDD 12 Q VNW pch L=4e-08 W=3.8e-07 
M46 Q 12 VDD VNW pch L=4e-08 W=3.8e-07 
M47 VDD 12 Q VNW pch L=4e-08 W=3.8e-07 
M48 VDD 16 15 VNW pch L=4e-08 W=2.9e-07 
M49 16 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT MX2_X0P5B_A9TR Y VDD VNW VPW VSS A B S0
M0 10 B 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS S0 10 VPW nch L=4e-08 W=1.2e-07 
M2 11 1 VSS VPW nch L=4e-08 W=1.7e-07 
M3 Y 5 11 VPW nch L=4e-08 W=1.7e-07 
M4 12 A 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 12 VPW nch L=4e-08 W=1.2e-07 
M6 6 S0 VSS VPW nch L=4e-08 W=1.2e-07 
M7 1 B VDD VNW pch L=4e-08 W=1.4e-07 
M8 VDD S0 1 VNW pch L=4e-08 W=1.4e-07 
M9 Y 1 VDD VNW pch L=4e-08 W=2e-07 
M10 VDD 5 Y VNW pch L=4e-08 W=2e-07 
M11 5 A VDD VNW pch L=4e-08 W=1.4e-07 
M12 VDD 6 5 VNW pch L=4e-08 W=1.4e-07 
M13 6 S0 VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT MX2_X0P7B_A9TR Y VDD VNW VPW VSS A B S0
M0 10 B 1 VPW nch L=4e-08 W=1.35e-07 
M1 VSS S0 10 VPW nch L=4e-08 W=1.35e-07 
M2 11 1 VSS VPW nch L=4e-08 W=2.45e-07 
M3 Y 5 11 VPW nch L=4e-08 W=2.45e-07 
M4 12 A 5 VPW nch L=4e-08 W=1.35e-07 
M5 VSS 6 12 VPW nch L=4e-08 W=1.35e-07 
M6 6 S0 VSS VPW nch L=4e-08 W=1.35e-07 
M7 1 B VDD VNW pch L=4e-08 W=1.6e-07 
M8 VDD S0 1 VNW pch L=4e-08 W=1.6e-07 
M9 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
M10 VDD 5 Y VNW pch L=4e-08 W=2.85e-07 
M11 5 A VDD VNW pch L=4e-08 W=1.6e-07 
M12 VDD 6 5 VNW pch L=4e-08 W=1.6e-07 
M13 6 S0 VDD VNW pch L=4e-08 W=1.6e-07 
.ENDS


.SUBCKT MX2_X1B_A9TR Y VDD VNW VPW VSS A B S0
M0 10 B 1 VPW nch L=4e-08 W=1.7e-07 
M1 VSS S0 10 VPW nch L=4e-08 W=1.7e-07 
M2 11 1 VSS VPW nch L=4e-08 W=3.45e-07 
M3 Y 5 11 VPW nch L=4e-08 W=3.45e-07 
M4 12 A 5 VPW nch L=4e-08 W=1.7e-07 
M5 VSS 6 12 VPW nch L=4e-08 W=1.7e-07 
M6 6 S0 VSS VPW nch L=4e-08 W=1.7e-07 
M7 1 B VDD VNW pch L=4e-08 W=1.95e-07 
M8 VDD S0 1 VNW pch L=4e-08 W=1.95e-07 
M9 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD 5 Y VNW pch L=4e-08 W=4e-07 
M11 5 A VDD VNW pch L=4e-08 W=1.95e-07 
M12 VDD 6 5 VNW pch L=4e-08 W=1.95e-07 
M13 6 S0 VDD VNW pch L=4e-08 W=1.95e-07 
.ENDS


.SUBCKT MX2_X1P4B_A9TR Y VDD VNW VPW VSS A B S0
M0 11 B 1 VPW nch L=4e-08 W=2.25e-07 
M1 VSS S0 11 VPW nch L=4e-08 W=2.25e-07 
M2 VSS 1 4 VPW nch L=4e-08 W=2.45e-07 
M3 4 1 VSS VPW nch L=4e-08 W=2.45e-07 
M4 Y 6 4 VPW nch L=4e-08 W=2.45e-07 
M5 4 6 Y VPW nch L=4e-08 W=2.45e-07 
M6 12 A 6 VPW nch L=4e-08 W=2.25e-07 
M7 VSS 7 12 VPW nch L=4e-08 W=2.25e-07 
M8 7 S0 VSS VPW nch L=4e-08 W=2.25e-07 
M9 1 B VDD VNW pch L=4e-08 W=2.6e-07 
M10 VDD S0 1 VNW pch L=4e-08 W=2.6e-07 
M11 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
M12 VDD 1 Y VNW pch L=4e-08 W=2.85e-07 
M13 Y 6 VDD VNW pch L=4e-08 W=2.85e-07 
M14 VDD 6 Y VNW pch L=4e-08 W=2.85e-07 
M15 6 A VDD VNW pch L=4e-08 W=2.6e-07 
M16 VDD 7 6 VNW pch L=4e-08 W=2.6e-07 
M17 7 S0 VDD VNW pch L=4e-08 W=2.6e-07 
.ENDS


.SUBCKT MX2_X2B_A9TR Y VDD VNW VPW VSS A B S0
M0 11 B 1 VPW nch L=4e-08 W=2.9e-07 
M1 VSS S0 11 VPW nch L=4e-08 W=2.9e-07 
M2 VSS 1 4 VPW nch L=4e-08 W=3.45e-07 
M3 4 1 VSS VPW nch L=4e-08 W=3.45e-07 
M4 Y 6 4 VPW nch L=4e-08 W=3.45e-07 
M5 4 6 Y VPW nch L=4e-08 W=3.45e-07 
M6 12 A 6 VPW nch L=4e-08 W=2.9e-07 
M7 VSS 7 12 VPW nch L=4e-08 W=2.9e-07 
M8 7 S0 VSS VPW nch L=4e-08 W=2.9e-07 
M9 1 B VDD VNW pch L=4e-08 W=3.35e-07 
M10 VDD S0 1 VNW pch L=4e-08 W=3.35e-07 
M11 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M12 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M13 Y 6 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD 6 Y VNW pch L=4e-08 W=4e-07 
M15 6 A VDD VNW pch L=4e-08 W=3.35e-07 
M16 VDD 7 6 VNW pch L=4e-08 W=3.35e-07 
M17 7 S0 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT MX2_X3B_A9TR Y VDD VNW VPW VSS A B S0
M0 10 4 VSS VPW nch L=4e-08 W=2.3e-07 
M1 3 A 10 VPW nch L=4e-08 W=2.3e-07 
M2 11 A 3 VPW nch L=4e-08 W=2.3e-07 
M3 VSS 4 11 VPW nch L=4e-08 W=2.3e-07 
M4 4 S0 VSS VPW nch L=4e-08 W=2.3e-07 
M5 VSS S0 4 VPW nch L=4e-08 W=2.3e-07 
M6 12 S0 VSS VPW nch L=4e-08 W=2.3e-07 
M7 5 B 12 VPW nch L=4e-08 W=2.3e-07 
M8 13 B 5 VPW nch L=4e-08 W=2.3e-07 
M9 VSS S0 13 VPW nch L=4e-08 W=2.3e-07 
M10 14 5 VSS VPW nch L=4e-08 W=3.45e-07 
M11 Y 3 14 VPW nch L=4e-08 W=3.45e-07 
M12 15 3 Y VPW nch L=4e-08 W=3.45e-07 
M13 VSS 5 15 VPW nch L=4e-08 W=3.45e-07 
M14 16 5 VSS VPW nch L=4e-08 W=3.45e-07 
M15 Y 3 16 VPW nch L=4e-08 W=3.45e-07 
M16 3 4 VDD VNW pch L=4e-08 W=2.7e-07 
M17 VDD A 3 VNW pch L=4e-08 W=2.7e-07 
M18 3 A VDD VNW pch L=4e-08 W=2.7e-07 
M19 VDD 4 3 VNW pch L=4e-08 W=2.7e-07 
M20 4 S0 VDD VNW pch L=4e-08 W=2.7e-07 
M21 VDD S0 4 VNW pch L=4e-08 W=2.7e-07 
M22 5 S0 VDD VNW pch L=4e-08 W=2.7e-07 
M23 VDD B 5 VNW pch L=4e-08 W=2.7e-07 
M24 5 B VDD VNW pch L=4e-08 W=2.7e-07 
M25 VDD S0 5 VNW pch L=4e-08 W=2.7e-07 
M26 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M28 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 5 Y VNW pch L=4e-08 W=4e-07 
M30 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT MX2_X4B_A9TR Y VDD VNW VPW VSS A B S0
M0 10 4 VSS VPW nch L=4e-08 W=2.95e-07 
M1 3 A 10 VPW nch L=4e-08 W=2.95e-07 
M2 11 A 3 VPW nch L=4e-08 W=2.95e-07 
M3 VSS 4 11 VPW nch L=4e-08 W=2.95e-07 
M4 4 S0 VSS VPW nch L=4e-08 W=2.95e-07 
M5 VSS S0 4 VPW nch L=4e-08 W=2.95e-07 
M6 12 S0 VSS VPW nch L=4e-08 W=2.95e-07 
M7 5 B 12 VPW nch L=4e-08 W=2.95e-07 
M8 13 B 5 VPW nch L=4e-08 W=2.95e-07 
M9 VSS S0 13 VPW nch L=4e-08 W=2.95e-07 
M10 14 5 VSS VPW nch L=4e-08 W=3.45e-07 
M11 Y 3 14 VPW nch L=4e-08 W=3.45e-07 
M12 15 3 Y VPW nch L=4e-08 W=3.45e-07 
M13 VSS 5 15 VPW nch L=4e-08 W=3.45e-07 
M14 16 5 VSS VPW nch L=4e-08 W=3.45e-07 
M15 Y 3 16 VPW nch L=4e-08 W=3.45e-07 
M16 17 3 Y VPW nch L=4e-08 W=3.45e-07 
M17 VSS 5 17 VPW nch L=4e-08 W=3.45e-07 
M18 3 4 VDD VNW pch L=4e-08 W=3.4e-07 
M19 VDD A 3 VNW pch L=4e-08 W=3.4e-07 
M20 3 A VDD VNW pch L=4e-08 W=3.4e-07 
M21 VDD 4 3 VNW pch L=4e-08 W=3.4e-07 
M22 4 S0 VDD VNW pch L=4e-08 W=3.4e-07 
M23 VDD S0 4 VNW pch L=4e-08 W=3.4e-07 
M24 5 S0 VDD VNW pch L=4e-08 W=3.4e-07 
M25 VDD B 5 VNW pch L=4e-08 W=3.4e-07 
M26 5 B VDD VNW pch L=4e-08 W=3.4e-07 
M27 VDD S0 5 VNW pch L=4e-08 W=3.4e-07 
M28 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M30 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 5 Y VNW pch L=4e-08 W=4e-07 
M32 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M33 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M34 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 5 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT MX2_X6B_A9TR Y VDD VNW VPW VSS A B S0
M0 10 A 1 VPW nch L=4e-08 W=3e-07 
M1 VSS 4 10 VPW nch L=4e-08 W=3e-07 
M2 11 4 VSS VPW nch L=4e-08 W=3e-07 
M3 1 A 11 VPW nch L=4e-08 W=3e-07 
M4 12 A 1 VPW nch L=4e-08 W=3e-07 
M5 VSS 4 12 VPW nch L=4e-08 W=3e-07 
M6 4 S0 VSS VPW nch L=4e-08 W=3e-07 
M7 VSS S0 4 VPW nch L=4e-08 W=3e-07 
M8 4 S0 VSS VPW nch L=4e-08 W=3e-07 
M9 13 S0 VSS VPW nch L=4e-08 W=3e-07 
M10 5 B 13 VPW nch L=4e-08 W=3e-07 
M11 14 B 5 VPW nch L=4e-08 W=3e-07 
M12 VSS S0 14 VPW nch L=4e-08 W=3e-07 
M13 15 S0 VSS VPW nch L=4e-08 W=3e-07 
M14 5 B 15 VPW nch L=4e-08 W=3e-07 
M15 16 5 VSS VPW nch L=4e-08 W=3.45e-07 
M16 Y 1 16 VPW nch L=4e-08 W=3.45e-07 
M17 17 1 Y VPW nch L=4e-08 W=3.45e-07 
M18 VSS 5 17 VPW nch L=4e-08 W=3.45e-07 
M19 18 5 VSS VPW nch L=4e-08 W=3.45e-07 
M20 Y 1 18 VPW nch L=4e-08 W=3.45e-07 
M21 19 1 Y VPW nch L=4e-08 W=3.45e-07 
M22 VSS 5 19 VPW nch L=4e-08 W=3.45e-07 
M23 20 5 VSS VPW nch L=4e-08 W=3.45e-07 
M24 Y 1 20 VPW nch L=4e-08 W=3.45e-07 
M25 21 1 Y VPW nch L=4e-08 W=3.45e-07 
M26 VSS 5 21 VPW nch L=4e-08 W=3.45e-07 
M27 1 A VDD VNW pch L=4e-08 W=3.5e-07 
M28 VDD 4 1 VNW pch L=4e-08 W=3.5e-07 
M29 1 4 VDD VNW pch L=4e-08 W=3.5e-07 
M30 VDD A 1 VNW pch L=4e-08 W=3.5e-07 
M31 1 A VDD VNW pch L=4e-08 W=3.5e-07 
M32 VDD 4 1 VNW pch L=4e-08 W=3.5e-07 
M33 4 S0 VDD VNW pch L=4e-08 W=3.5e-07 
M34 VDD S0 4 VNW pch L=4e-08 W=3.5e-07 
M35 4 S0 VDD VNW pch L=4e-08 W=3.5e-07 
M36 5 S0 VDD VNW pch L=4e-08 W=3.5e-07 
M37 VDD B 5 VNW pch L=4e-08 W=3.5e-07 
M38 5 B VDD VNW pch L=4e-08 W=3.5e-07 
M39 VDD S0 5 VNW pch L=4e-08 W=3.5e-07 
M40 5 S0 VDD VNW pch L=4e-08 W=3.5e-07 
M41 VDD B 5 VNW pch L=4e-08 W=3.5e-07 
M42 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M43 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M44 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M45 VDD 5 Y VNW pch L=4e-08 W=4e-07 
M46 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M47 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M48 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M49 VDD 5 Y VNW pch L=4e-08 W=4e-07 
M50 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M51 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M52 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M53 VDD 5 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT MX2_X8B_A9TR Y VDD VNW VPW VSS A B S0
M0 10 4 VSS VPW nch L=4e-08 W=3e-07 
M1 3 A 10 VPW nch L=4e-08 W=3e-07 
M2 11 A 3 VPW nch L=4e-08 W=3e-07 
M3 VSS 4 11 VPW nch L=4e-08 W=3e-07 
M4 12 4 VSS VPW nch L=4e-08 W=3e-07 
M5 3 A 12 VPW nch L=4e-08 W=3e-07 
M6 13 A 3 VPW nch L=4e-08 W=3e-07 
M7 VSS 4 13 VPW nch L=4e-08 W=3e-07 
M8 4 S0 VSS VPW nch L=4e-08 W=3e-07 
M9 VSS S0 4 VPW nch L=4e-08 W=3e-07 
M10 4 S0 VSS VPW nch L=4e-08 W=3e-07 
M11 VSS S0 4 VPW nch L=4e-08 W=3e-07 
M12 14 S0 VSS VPW nch L=4e-08 W=3e-07 
M13 5 B 14 VPW nch L=4e-08 W=3e-07 
M14 15 B 5 VPW nch L=4e-08 W=3e-07 
M15 VSS S0 15 VPW nch L=4e-08 W=3e-07 
M16 16 S0 VSS VPW nch L=4e-08 W=3e-07 
M17 5 B 16 VPW nch L=4e-08 W=3e-07 
M18 17 B 5 VPW nch L=4e-08 W=3e-07 
M19 VSS S0 17 VPW nch L=4e-08 W=3e-07 
M20 18 5 VSS VPW nch L=4e-08 W=3.45e-07 
M21 Y 3 18 VPW nch L=4e-08 W=3.45e-07 
M22 19 3 Y VPW nch L=4e-08 W=3.45e-07 
M23 VSS 5 19 VPW nch L=4e-08 W=3.45e-07 
M24 20 5 VSS VPW nch L=4e-08 W=3.45e-07 
M25 Y 3 20 VPW nch L=4e-08 W=3.45e-07 
M26 21 3 Y VPW nch L=4e-08 W=3.45e-07 
M27 VSS 5 21 VPW nch L=4e-08 W=3.45e-07 
M28 22 5 VSS VPW nch L=4e-08 W=3.45e-07 
M29 Y 3 22 VPW nch L=4e-08 W=3.45e-07 
M30 23 3 Y VPW nch L=4e-08 W=3.45e-07 
M31 VSS 5 23 VPW nch L=4e-08 W=3.45e-07 
M32 24 5 VSS VPW nch L=4e-08 W=3.45e-07 
M33 Y 3 24 VPW nch L=4e-08 W=3.45e-07 
M34 25 3 Y VPW nch L=4e-08 W=3.45e-07 
M35 VSS 5 25 VPW nch L=4e-08 W=3.45e-07 
M36 3 4 VDD VNW pch L=4e-08 W=3.5e-07 
M37 VDD A 3 VNW pch L=4e-08 W=3.5e-07 
M38 3 A VDD VNW pch L=4e-08 W=3.5e-07 
M39 VDD 4 3 VNW pch L=4e-08 W=3.5e-07 
M40 3 4 VDD VNW pch L=4e-08 W=3.5e-07 
M41 VDD A 3 VNW pch L=4e-08 W=3.5e-07 
M42 3 A VDD VNW pch L=4e-08 W=3.5e-07 
M43 VDD 4 3 VNW pch L=4e-08 W=3.5e-07 
M44 4 S0 VDD VNW pch L=4e-08 W=3.5e-07 
M45 VDD S0 4 VNW pch L=4e-08 W=3.5e-07 
M46 4 S0 VDD VNW pch L=4e-08 W=3.5e-07 
M47 VDD S0 4 VNW pch L=4e-08 W=3.5e-07 
M48 5 S0 VDD VNW pch L=4e-08 W=3.5e-07 
M49 VDD B 5 VNW pch L=4e-08 W=3.5e-07 
M50 5 B VDD VNW pch L=4e-08 W=3.5e-07 
M51 VDD S0 5 VNW pch L=4e-08 W=3.5e-07 
M52 5 S0 VDD VNW pch L=4e-08 W=3.5e-07 
M53 VDD B 5 VNW pch L=4e-08 W=3.5e-07 
M54 5 B VDD VNW pch L=4e-08 W=3.5e-07 
M55 VDD S0 5 VNW pch L=4e-08 W=3.5e-07 
M56 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M57 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M58 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M59 VDD 5 Y VNW pch L=4e-08 W=4e-07 
M60 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M61 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M62 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M63 VDD 5 Y VNW pch L=4e-08 W=4e-07 
M64 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M65 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M66 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M67 VDD 5 Y VNW pch L=4e-08 W=4e-07 
M68 Y 5 VDD VNW pch L=4e-08 W=4e-07 
M69 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M70 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M71 VDD 5 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT MXGL2_X0P5B_A9TR Y VDD VNW VPW VSS A B S0
M0 11 B 1 VPW nch L=4e-08 W=1.35e-07 
M1 VSS S0 11 VPW nch L=4e-08 W=1.35e-07 
M2 VSS S0 4 VPW nch L=4e-08 W=1.35e-07 
M3 12 4 VSS VPW nch L=4e-08 W=1.35e-07 
M4 5 A 12 VPW nch L=4e-08 W=1.35e-07 
M5 13 5 Y VPW nch L=4e-08 W=2e-07 
M6 14 1 13 VPW nch L=4e-08 W=2e-07 
M7 VSS 7 14 VPW nch L=4e-08 W=2e-07 
M8 15 B VSS VPW nch L=4e-08 W=1.2e-07 
M9 7 A 15 VPW nch L=4e-08 W=1.2e-07 
M10 1 B VDD VNW pch L=4e-08 W=1.55e-07 
M11 VDD S0 1 VNW pch L=4e-08 W=1.55e-07 
M12 VDD S0 4 VNW pch L=4e-08 W=1.75e-07 
M13 5 4 VDD VNW pch L=4e-08 W=1.55e-07 
M14 VDD A 5 VNW pch L=4e-08 W=1.55e-07 
M15 VDD 5 Y VNW pch L=4e-08 W=1.75e-07 
M16 Y 1 VDD VNW pch L=4e-08 W=1.75e-07 
M17 VDD 7 Y VNW pch L=4e-08 W=1.75e-07 
M18 7 B VDD VNW pch L=4e-08 W=1.45e-07 
M19 VDD A 7 VNW pch L=4e-08 W=1.45e-07 
.ENDS


.SUBCKT MXGL2_X0P7B_A9TR Y VDD VNW VPW VSS A B S0
M0 11 B 1 VPW nch L=4e-08 W=1.6e-07 
M1 VSS S0 11 VPW nch L=4e-08 W=1.6e-07 
M2 VSS S0 4 VPW nch L=4e-08 W=1.5e-07 
M3 12 4 VSS VPW nch L=4e-08 W=1.6e-07 
M4 5 A 12 VPW nch L=4e-08 W=1.6e-07 
M5 13 5 Y VPW nch L=4e-08 W=2.8e-07 
M6 14 1 13 VPW nch L=4e-08 W=2.8e-07 
M7 VSS 7 14 VPW nch L=4e-08 W=2.8e-07 
M8 15 B VSS VPW nch L=4e-08 W=1.2e-07 
M9 7 A 15 VPW nch L=4e-08 W=1.2e-07 
M10 1 B VDD VNW pch L=4e-08 W=1.85e-07 
M11 VDD S0 1 VNW pch L=4e-08 W=1.85e-07 
M12 VDD S0 4 VNW pch L=4e-08 W=1.95e-07 
M13 5 4 VDD VNW pch L=4e-08 W=1.85e-07 
M14 VDD A 5 VNW pch L=4e-08 W=1.85e-07 
M15 VDD 5 Y VNW pch L=4e-08 W=2.4e-07 
M16 Y 1 VDD VNW pch L=4e-08 W=2.4e-07 
M17 VDD 7 Y VNW pch L=4e-08 W=2.4e-07 
M18 7 B VDD VNW pch L=4e-08 W=1.45e-07 
M19 VDD A 7 VNW pch L=4e-08 W=1.45e-07 
.ENDS


.SUBCKT MXGL2_X1B_A9TR Y VDD VNW VPW VSS A B S0
M0 11 B 1 VPW nch L=4e-08 W=1.9e-07 
M1 VSS S0 11 VPW nch L=4e-08 W=1.9e-07 
M2 VSS S0 4 VPW nch L=4e-08 W=1.65e-07 
M3 12 4 VSS VPW nch L=4e-08 W=1.9e-07 
M4 5 A 12 VPW nch L=4e-08 W=1.9e-07 
M5 13 5 Y VPW nch L=4e-08 W=4e-07 
M6 14 1 13 VPW nch L=4e-08 W=4e-07 
M7 VSS 7 14 VPW nch L=4e-08 W=4e-07 
M8 15 B VSS VPW nch L=4e-08 W=1.2e-07 
M9 7 A 15 VPW nch L=4e-08 W=1.2e-07 
M10 1 B VDD VNW pch L=4e-08 W=2.2e-07 
M11 VDD S0 1 VNW pch L=4e-08 W=2.2e-07 
M12 VDD S0 4 VNW pch L=4e-08 W=2.1e-07 
M13 5 4 VDD VNW pch L=4e-08 W=2.2e-07 
M14 VDD A 5 VNW pch L=4e-08 W=2.2e-07 
M15 VDD 5 Y VNW pch L=4e-08 W=3.45e-07 
M16 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M17 VDD 7 Y VNW pch L=4e-08 W=3.45e-07 
M18 7 B VDD VNW pch L=4e-08 W=1.45e-07 
M19 VDD A 7 VNW pch L=4e-08 W=1.45e-07 
.ENDS


.SUBCKT MXGL2_X1P4B_A9TR Y VDD VNW VPW VSS A B S0
M0 11 B 1 VPW nch L=4e-08 W=2.45e-07 
M1 VSS S0 11 VPW nch L=4e-08 W=2.45e-07 
M2 VSS S0 4 VPW nch L=4e-08 W=1.9e-07 
M3 12 4 VSS VPW nch L=4e-08 W=2.45e-07 
M4 5 A 12 VPW nch L=4e-08 W=2.45e-07 
M5 13 7 VSS VPW nch L=4e-08 W=2.8e-07 
M6 14 1 13 VPW nch L=4e-08 W=2.8e-07 
M7 Y 5 14 VPW nch L=4e-08 W=2.8e-07 
M8 15 5 Y VPW nch L=4e-08 W=2.8e-07 
M9 16 1 15 VPW nch L=4e-08 W=2.8e-07 
M10 VSS 7 16 VPW nch L=4e-08 W=2.8e-07 
M11 17 B VSS VPW nch L=4e-08 W=1.2e-07 
M12 7 A 17 VPW nch L=4e-08 W=1.2e-07 
M13 1 B VDD VNW pch L=4e-08 W=2.85e-07 
M14 VDD S0 1 VNW pch L=4e-08 W=2.85e-07 
M15 VDD S0 4 VNW pch L=4e-08 W=2.45e-07 
M16 5 4 VDD VNW pch L=4e-08 W=2.85e-07 
M17 VDD A 5 VNW pch L=4e-08 W=2.85e-07 
M18 Y 7 VDD VNW pch L=4e-08 W=2.4e-07 
M19 VDD 1 Y VNW pch L=4e-08 W=2.4e-07 
M20 Y 5 VDD VNW pch L=4e-08 W=2.4e-07 
M21 VDD 5 Y VNW pch L=4e-08 W=2.4e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=2.4e-07 
M23 VDD 7 Y VNW pch L=4e-08 W=2.4e-07 
M24 7 B VDD VNW pch L=4e-08 W=1.45e-07 
M25 VDD A 7 VNW pch L=4e-08 W=1.45e-07 
.ENDS


.SUBCKT MXGL2_X2B_A9TR Y VDD VNW VPW VSS A B S0
M0 11 B 1 VPW nch L=4e-08 W=3.15e-07 
M1 VSS S0 11 VPW nch L=4e-08 W=3.15e-07 
M2 VSS S0 4 VPW nch L=4e-08 W=2.2e-07 
M3 12 4 VSS VPW nch L=4e-08 W=3.15e-07 
M4 5 A 12 VPW nch L=4e-08 W=3.15e-07 
M5 13 7 VSS VPW nch L=4e-08 W=3.9e-07 
M6 14 1 13 VPW nch L=4e-08 W=3.9e-07 
M7 Y 5 14 VPW nch L=4e-08 W=3.9e-07 
M8 15 5 Y VPW nch L=4e-08 W=3.9e-07 
M9 16 1 15 VPW nch L=4e-08 W=3.9e-07 
M10 VSS 7 16 VPW nch L=4e-08 W=3.9e-07 
M11 17 B VSS VPW nch L=4e-08 W=1.55e-07 
M12 7 A 17 VPW nch L=4e-08 W=1.55e-07 
M13 1 B VDD VNW pch L=4e-08 W=3.65e-07 
M14 VDD S0 1 VNW pch L=4e-08 W=3.65e-07 
M15 VDD S0 4 VNW pch L=4e-08 W=2.85e-07 
M16 5 4 VDD VNW pch L=4e-08 W=3.65e-07 
M17 VDD A 5 VNW pch L=4e-08 W=3.65e-07 
M18 Y 7 VDD VNW pch L=4e-08 W=3.35e-07 
M19 VDD 1 Y VNW pch L=4e-08 W=3.35e-07 
M20 Y 5 VDD VNW pch L=4e-08 W=3.35e-07 
M21 VDD 5 Y VNW pch L=4e-08 W=3.35e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
M23 VDD 7 Y VNW pch L=4e-08 W=3.35e-07 
M24 7 B VDD VNW pch L=4e-08 W=1.8e-07 
M25 VDD A 7 VNW pch L=4e-08 W=1.8e-07 
.ENDS


.SUBCKT MXGL2_X3B_A9TR Y VDD VNW VPW VSS A B S0
M0 12 S0 VSS VPW nch L=4e-08 W=2.35e-07 
M1 3 B 12 VPW nch L=4e-08 W=2.35e-07 
M2 13 B 3 VPW nch L=4e-08 W=2.35e-07 
M3 VSS S0 13 VPW nch L=4e-08 W=2.35e-07 
M4 VSS S0 4 VPW nch L=4e-08 W=3.1e-07 
M5 14 4 VSS VPW nch L=4e-08 W=2.35e-07 
M6 5 A 14 VPW nch L=4e-08 W=2.35e-07 
M7 15 A 5 VPW nch L=4e-08 W=2.35e-07 
M8 VSS 4 15 VPW nch L=4e-08 W=2.35e-07 
M9 16 5 Y VPW nch L=4e-08 W=4e-07 
M10 7 3 16 VPW nch L=4e-08 W=4e-07 
M11 17 3 7 VPW nch L=4e-08 W=4e-07 
M12 Y 5 17 VPW nch L=4e-08 W=4e-07 
M13 18 5 Y VPW nch L=4e-08 W=4e-07 
M14 7 3 18 VPW nch L=4e-08 W=4e-07 
M15 VSS 8 7 VPW nch L=4e-08 W=4e-07 
M16 7 8 VSS VPW nch L=4e-08 W=4e-07 
M17 VSS 8 7 VPW nch L=4e-08 W=4e-07 
M18 19 B VSS VPW nch L=4e-08 W=2.35e-07 
M19 8 A 19 VPW nch L=4e-08 W=2.35e-07 
M20 3 S0 VDD VNW pch L=4e-08 W=2.75e-07 
M21 VDD B 3 VNW pch L=4e-08 W=2.75e-07 
M22 3 B VDD VNW pch L=4e-08 W=2.75e-07 
M23 VDD S0 3 VNW pch L=4e-08 W=2.75e-07 
M24 VDD S0 4 VNW pch L=4e-08 W=4e-07 
M25 5 4 VDD VNW pch L=4e-08 W=2.75e-07 
M26 VDD A 5 VNW pch L=4e-08 W=2.75e-07 
M27 5 A VDD VNW pch L=4e-08 W=2.75e-07 
M28 VDD 4 5 VNW pch L=4e-08 W=2.75e-07 
M29 VDD 5 Y VNW pch L=4e-08 W=3.45e-07 
M30 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M31 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M32 Y 5 VDD VNW pch L=4e-08 W=3.45e-07 
M33 VDD 5 Y VNW pch L=4e-08 W=3.45e-07 
M34 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M35 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M36 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M37 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M38 8 B VDD VNW pch L=4e-08 W=2.75e-07 
M39 VDD A 8 VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT MXGL2_X4B_A9TR Y VDD VNW VPW VSS A B S0
M0 12 S0 VSS VPW nch L=4e-08 W=3.1e-07 
M1 3 B 12 VPW nch L=4e-08 W=3.1e-07 
M2 13 B 3 VPW nch L=4e-08 W=3.1e-07 
M3 VSS S0 13 VPW nch L=4e-08 W=3.1e-07 
M4 4 S0 VSS VPW nch L=4e-08 W=1.9e-07 
M5 VSS S0 4 VPW nch L=4e-08 W=1.9e-07 
M6 14 4 VSS VPW nch L=4e-08 W=3.1e-07 
M7 5 A 14 VPW nch L=4e-08 W=3.1e-07 
M8 15 A 5 VPW nch L=4e-08 W=3.1e-07 
M9 VSS 4 15 VPW nch L=4e-08 W=3.1e-07 
M10 16 3 6 VPW nch L=4e-08 W=4e-07 
M11 Y 5 16 VPW nch L=4e-08 W=4e-07 
M12 17 5 Y VPW nch L=4e-08 W=4e-07 
M13 6 3 17 VPW nch L=4e-08 W=4e-07 
M14 18 3 6 VPW nch L=4e-08 W=4e-07 
M15 Y 5 18 VPW nch L=4e-08 W=4e-07 
M16 19 5 Y VPW nch L=4e-08 W=4e-07 
M17 6 3 19 VPW nch L=4e-08 W=4e-07 
M18 VSS 8 6 VPW nch L=4e-08 W=4e-07 
M19 6 8 VSS VPW nch L=4e-08 W=4e-07 
M20 VSS 8 6 VPW nch L=4e-08 W=4e-07 
M21 6 8 VSS VPW nch L=4e-08 W=4e-07 
M22 20 B VSS VPW nch L=4e-08 W=3.1e-07 
M23 8 A 20 VPW nch L=4e-08 W=3.1e-07 
M24 3 S0 VDD VNW pch L=4e-08 W=3.6e-07 
M25 VDD B 3 VNW pch L=4e-08 W=3.6e-07 
M26 3 B VDD VNW pch L=4e-08 W=3.6e-07 
M27 VDD S0 3 VNW pch L=4e-08 W=3.6e-07 
M28 4 S0 VDD VNW pch L=4e-08 W=2.45e-07 
M29 VDD S0 4 VNW pch L=4e-08 W=2.45e-07 
M30 5 4 VDD VNW pch L=4e-08 W=3.6e-07 
M31 VDD A 5 VNW pch L=4e-08 W=3.6e-07 
M32 5 A VDD VNW pch L=4e-08 W=3.6e-07 
M33 VDD 4 5 VNW pch L=4e-08 W=3.6e-07 
M34 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M35 Y 5 VDD VNW pch L=4e-08 W=3.45e-07 
M36 VDD 5 Y VNW pch L=4e-08 W=3.45e-07 
M37 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M38 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M39 Y 5 VDD VNW pch L=4e-08 W=3.45e-07 
M40 VDD 5 Y VNW pch L=4e-08 W=3.45e-07 
M41 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M42 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M43 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M44 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M45 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M46 8 B VDD VNW pch L=4e-08 W=3.6e-07 
M47 VDD A 8 VNW pch L=4e-08 W=3.6e-07 
.ENDS


.SUBCKT MXGL2_X6B_A9TR Y VDD VNW VPW VSS A B S0
M0 12 S0 VSS VPW nch L=4e-08 W=3.15e-07 
M1 3 B 12 VPW nch L=4e-08 W=3.15e-07 
M2 13 B 3 VPW nch L=4e-08 W=3.15e-07 
M3 VSS S0 13 VPW nch L=4e-08 W=3.15e-07 
M4 14 S0 VSS VPW nch L=4e-08 W=3.15e-07 
M5 3 B 14 VPW nch L=4e-08 W=3.15e-07 
M6 4 S0 VSS VPW nch L=4e-08 W=2.8e-07 
M7 VSS S0 4 VPW nch L=4e-08 W=2.8e-07 
M8 15 4 VSS VPW nch L=4e-08 W=3.15e-07 
M9 5 A 15 VPW nch L=4e-08 W=3.15e-07 
M10 16 A 5 VPW nch L=4e-08 W=3.15e-07 
M11 VSS 4 16 VPW nch L=4e-08 W=3.15e-07 
M12 17 4 VSS VPW nch L=4e-08 W=3.15e-07 
M13 5 A 17 VPW nch L=4e-08 W=3.15e-07 
M14 18 3 6 VPW nch L=4e-08 W=4e-07 
M15 Y 5 18 VPW nch L=4e-08 W=4e-07 
M16 19 5 Y VPW nch L=4e-08 W=4e-07 
M17 6 3 19 VPW nch L=4e-08 W=4e-07 
M18 20 3 6 VPW nch L=4e-08 W=4e-07 
M19 Y 5 20 VPW nch L=4e-08 W=4e-07 
M20 21 5 Y VPW nch L=4e-08 W=4e-07 
M21 6 3 21 VPW nch L=4e-08 W=4e-07 
M22 22 3 6 VPW nch L=4e-08 W=4e-07 
M23 Y 5 22 VPW nch L=4e-08 W=4e-07 
M24 23 5 Y VPW nch L=4e-08 W=4e-07 
M25 6 3 23 VPW nch L=4e-08 W=4e-07 
M26 VSS 8 6 VPW nch L=4e-08 W=4e-07 
M27 6 8 VSS VPW nch L=4e-08 W=4e-07 
M28 VSS 8 6 VPW nch L=4e-08 W=4e-07 
M29 6 8 VSS VPW nch L=4e-08 W=4e-07 
M30 VSS 8 6 VPW nch L=4e-08 W=4e-07 
M31 6 8 VSS VPW nch L=4e-08 W=4e-07 
M32 24 B VSS VPW nch L=4e-08 W=2.35e-07 
M33 8 A 24 VPW nch L=4e-08 W=2.35e-07 
M34 25 A 8 VPW nch L=4e-08 W=2.35e-07 
M35 VSS B 25 VPW nch L=4e-08 W=2.35e-07 
M36 3 S0 VDD VNW pch L=4e-08 W=3.65e-07 
M37 VDD B 3 VNW pch L=4e-08 W=3.65e-07 
M38 3 B VDD VNW pch L=4e-08 W=3.65e-07 
M39 VDD S0 3 VNW pch L=4e-08 W=3.65e-07 
M40 3 S0 VDD VNW pch L=4e-08 W=3.65e-07 
M41 VDD B 3 VNW pch L=4e-08 W=3.65e-07 
M42 4 S0 VDD VNW pch L=4e-08 W=3.6e-07 
M43 VDD S0 4 VNW pch L=4e-08 W=3.6e-07 
M44 5 4 VDD VNW pch L=4e-08 W=3.65e-07 
M45 VDD A 5 VNW pch L=4e-08 W=3.65e-07 
M46 5 A VDD VNW pch L=4e-08 W=3.65e-07 
M47 VDD 4 5 VNW pch L=4e-08 W=3.65e-07 
M48 5 4 VDD VNW pch L=4e-08 W=3.65e-07 
M49 VDD A 5 VNW pch L=4e-08 W=3.65e-07 
M50 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M51 VDD 5 Y VNW pch L=4e-08 W=3.45e-07 
M52 Y 5 VDD VNW pch L=4e-08 W=3.45e-07 
M53 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M54 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M55 VDD 5 Y VNW pch L=4e-08 W=3.45e-07 
M56 Y 5 VDD VNW pch L=4e-08 W=3.45e-07 
M57 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M58 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M59 VDD 5 Y VNW pch L=4e-08 W=3.45e-07 
M60 Y 5 VDD VNW pch L=4e-08 W=3.45e-07 
M61 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M62 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M63 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M64 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M65 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M66 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M67 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M68 8 B VDD VNW pch L=4e-08 W=2.75e-07 
M69 VDD A 8 VNW pch L=4e-08 W=2.75e-07 
M70 8 A VDD VNW pch L=4e-08 W=2.75e-07 
M71 VDD B 8 VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT MXIT2_X0P5M_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.2e-07 
M2 Y S0 1 VPW nch L=4e-08 W=1.2e-07 
M3 6 4 Y VPW nch L=4e-08 W=1.2e-07 
M4 VSS A 6 VPW nch L=4e-08 W=1.2e-07 
M5 VDD B 1 VNW pch L=4e-08 W=1.9e-07 
M6 4 S0 VDD VNW pch L=4e-08 W=1.9e-07 
M7 Y 4 1 VNW pch L=4e-08 W=1.9e-07 
M8 6 S0 Y VNW pch L=4e-08 W=1.9e-07 
M9 VDD A 6 VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT MXIT2_X0P7M_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=1.5e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.5e-07 
M2 Y S0 1 VPW nch L=4e-08 W=1.5e-07 
M3 6 4 Y VPW nch L=4e-08 W=1.5e-07 
M4 VSS A 6 VPW nch L=4e-08 W=1.5e-07 
M5 VDD B 1 VNW pch L=4e-08 W=2.25e-07 
M6 4 S0 VDD VNW pch L=4e-08 W=2.25e-07 
M7 Y 4 1 VNW pch L=4e-08 W=2.25e-07 
M8 6 S0 Y VNW pch L=4e-08 W=2.25e-07 
M9 VDD A 6 VNW pch L=4e-08 W=2.25e-07 
.ENDS


.SUBCKT MXIT2_X1M_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=2.6e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.6e-07 
M2 Y S0 1 VPW nch L=4e-08 W=2.6e-07 
M3 5 4 Y VPW nch L=4e-08 W=2.6e-07 
M4 VSS A 5 VPW nch L=4e-08 W=2.6e-07 
M5 VDD B 1 VNW pch L=4e-08 W=4e-07 
M6 4 S0 VDD VNW pch L=4e-08 W=4e-07 
M7 Y S0 5 VNW pch L=4e-08 W=4e-07 
M8 1 4 Y VNW pch L=4e-08 W=4e-07 
M9 VDD A 5 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT MXIT2_X1P4M_A9TR Y VDD VNW VPW VSS A B S0
M0 3 B VSS VPW nch L=4e-08 W=1.9e-07 
M1 VSS B 3 VPW nch L=4e-08 W=1.9e-07 
M2 4 S0 VSS VPW nch L=4e-08 W=1.9e-07 
M3 VSS S0 4 VPW nch L=4e-08 W=1.9e-07 
M4 Y S0 3 VPW nch L=4e-08 W=3.8e-07 
M5 5 4 Y VPW nch L=4e-08 W=3.8e-07 
M6 5 A VSS VPW nch L=4e-08 W=1.9e-07 
M7 VSS A 5 VPW nch L=4e-08 W=1.9e-07 
M8 3 B VDD VNW pch L=4e-08 W=3.3e-07 
M9 VDD B 3 VNW pch L=4e-08 W=3.3e-07 
M10 4 S0 VDD VNW pch L=4e-08 W=3.3e-07 
M11 VDD S0 4 VNW pch L=4e-08 W=3.3e-07 
M12 Y S0 5 VNW pch L=4e-08 W=4e-07 
M13 3 4 Y VNW pch L=4e-08 W=4e-07 
M14 5 A VDD VNW pch L=4e-08 W=3.3e-07 
M15 VDD A 5 VNW pch L=4e-08 W=3.3e-07 
.ENDS


.SUBCKT MXIT2_X2M_A9TR Y VDD VNW VPW VSS A B S0
M0 3 B VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.45e-07 
M2 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M3 VSS S0 4 VPW nch L=4e-08 W=2.45e-07 
M4 3 S0 Y VPW nch L=4e-08 W=2.45e-07 
M5 Y S0 3 VPW nch L=4e-08 W=2.45e-07 
M6 6 4 Y VPW nch L=4e-08 W=2.45e-07 
M7 Y 4 6 VPW nch L=4e-08 W=2.45e-07 
M8 6 A VSS VPW nch L=4e-08 W=2.45e-07 
M9 VSS A 6 VPW nch L=4e-08 W=2.45e-07 
M10 3 B VDD VNW pch L=4e-08 W=3.8e-07 
M11 VDD B 3 VNW pch L=4e-08 W=3.8e-07 
M12 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M13 VDD S0 4 VNW pch L=4e-08 W=3.8e-07 
M14 6 S0 Y VNW pch L=4e-08 W=3.8e-07 
M15 Y S0 6 VNW pch L=4e-08 W=3.8e-07 
M16 3 4 Y VNW pch L=4e-08 W=3.8e-07 
M17 Y 4 3 VNW pch L=4e-08 W=3.8e-07 
M18 6 A VDD VNW pch L=4e-08 W=3.8e-07 
M19 VDD A 6 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXIT2_X3M_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=2.45e-07 
M1 1 B VSS VPW nch L=4e-08 W=2.45e-07 
M2 VSS B 1 VPW nch L=4e-08 W=2.45e-07 
M3 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M4 VSS S0 4 VPW nch L=4e-08 W=2.45e-07 
M5 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M6 Y S0 1 VPW nch L=4e-08 W=2.45e-07 
M7 1 S0 Y VPW nch L=4e-08 W=2.45e-07 
M8 Y S0 1 VPW nch L=4e-08 W=2.45e-07 
M9 5 4 Y VPW nch L=4e-08 W=2.45e-07 
M10 Y 4 5 VPW nch L=4e-08 W=2.45e-07 
M11 5 4 Y VPW nch L=4e-08 W=2.45e-07 
M12 5 A VSS VPW nch L=4e-08 W=2.45e-07 
M13 VSS A 5 VPW nch L=4e-08 W=2.45e-07 
M14 5 A VSS VPW nch L=4e-08 W=2.45e-07 
M15 VDD B 1 VNW pch L=4e-08 W=3.8e-07 
M16 1 B VDD VNW pch L=4e-08 W=3.8e-07 
M17 VDD B 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M19 VDD S0 4 VNW pch L=4e-08 W=3.8e-07 
M20 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M21 Y S0 5 VNW pch L=4e-08 W=3.8e-07 
M22 5 S0 Y VNW pch L=4e-08 W=3.8e-07 
M23 Y S0 5 VNW pch L=4e-08 W=3.8e-07 
M24 1 4 Y VNW pch L=4e-08 W=3.8e-07 
M25 Y 4 1 VNW pch L=4e-08 W=3.8e-07 
M26 1 4 Y VNW pch L=4e-08 W=3.8e-07 
M27 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M28 VDD A 5 VNW pch L=4e-08 W=3.8e-07 
M29 5 A VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXIT2_X4M_A9TR Y VDD VNW VPW VSS A B S0
M0 3 B VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.45e-07 
M2 3 B VSS VPW nch L=4e-08 W=2.45e-07 
M3 VSS B 3 VPW nch L=4e-08 W=2.45e-07 
M4 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M5 VSS S0 4 VPW nch L=4e-08 W=2.45e-07 
M6 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M7 VSS S0 4 VPW nch L=4e-08 W=2.45e-07 
M8 3 S0 Y VPW nch L=4e-08 W=2.45e-07 
M9 Y S0 3 VPW nch L=4e-08 W=2.45e-07 
M10 3 S0 Y VPW nch L=4e-08 W=2.45e-07 
M11 Y S0 3 VPW nch L=4e-08 W=2.45e-07 
M12 6 4 Y VPW nch L=4e-08 W=2.45e-07 
M13 Y 4 6 VPW nch L=4e-08 W=2.45e-07 
M14 6 4 Y VPW nch L=4e-08 W=2.45e-07 
M15 Y 4 6 VPW nch L=4e-08 W=2.45e-07 
M16 6 A VSS VPW nch L=4e-08 W=2.45e-07 
M17 VSS A 6 VPW nch L=4e-08 W=2.45e-07 
M18 6 A VSS VPW nch L=4e-08 W=2.45e-07 
M19 VSS A 6 VPW nch L=4e-08 W=2.45e-07 
M20 3 B VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD B 3 VNW pch L=4e-08 W=3.8e-07 
M22 3 B VDD VNW pch L=4e-08 W=3.8e-07 
M23 VDD B 3 VNW pch L=4e-08 W=3.8e-07 
M24 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD S0 4 VNW pch L=4e-08 W=3.8e-07 
M26 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD S0 4 VNW pch L=4e-08 W=3.8e-07 
M28 6 S0 Y VNW pch L=4e-08 W=3.8e-07 
M29 Y S0 6 VNW pch L=4e-08 W=3.8e-07 
M30 6 S0 Y VNW pch L=4e-08 W=3.8e-07 
M31 Y S0 6 VNW pch L=4e-08 W=3.8e-07 
M32 3 4 Y VNW pch L=4e-08 W=3.8e-07 
M33 Y 4 3 VNW pch L=4e-08 W=3.8e-07 
M34 3 4 Y VNW pch L=4e-08 W=3.8e-07 
M35 Y 4 3 VNW pch L=4e-08 W=3.8e-07 
M36 6 A VDD VNW pch L=4e-08 W=3.8e-07 
M37 VDD A 6 VNW pch L=4e-08 W=3.8e-07 
M38 6 A VDD VNW pch L=4e-08 W=3.8e-07 
M39 VDD A 6 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXIT4_X0P5M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=1.55e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.2e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.55e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.55e-07 
M4 VSS C 5 VPW nch L=4e-08 W=1.55e-07 
M5 VSS 6 7 VPW nch L=4e-08 W=1.55e-07 
M6 8 S1 VSS VPW nch L=4e-08 W=1.55e-07 
M7 10 S1 7 VPW nch L=4e-08 W=1.55e-07 
M8 9 8 10 VPW nch L=4e-08 W=1.55e-07 
M9 Y 10 VSS VPW nch L=4e-08 W=1.55e-07 
M10 VSS 14 9 VPW nch L=4e-08 W=1.55e-07 
M11 12 A VSS VPW nch L=4e-08 W=1.55e-07 
M12 14 15 12 VPW nch L=4e-08 W=1.55e-07 
M13 13 S0 14 VPW nch L=4e-08 W=1.55e-07 
M14 VSS S0 15 VPW nch L=4e-08 W=1.2e-07 
M15 13 B VSS VPW nch L=4e-08 W=1.55e-07 
M16 VDD D 1 VNW pch L=4e-08 W=2.35e-07 
M17 4 S0 VDD VNW pch L=4e-08 W=1.9e-07 
M18 6 S0 5 VNW pch L=4e-08 W=2.35e-07 
M19 1 4 6 VNW pch L=4e-08 W=2.35e-07 
M20 VDD C 5 VNW pch L=4e-08 W=2.35e-07 
M21 VDD 6 7 VNW pch L=4e-08 W=1.8e-07 
M22 8 S1 VDD VNW pch L=4e-08 W=1.8e-07 
M23 10 S1 9 VNW pch L=4e-08 W=1.8e-07 
M24 7 8 10 VNW pch L=4e-08 W=1.8e-07 
M25 Y 10 VDD VNW pch L=4e-08 W=2e-07 
M26 VDD 14 9 VNW pch L=4e-08 W=1.8e-07 
M27 12 A VDD VNW pch L=4e-08 W=2.35e-07 
M28 14 15 13 VNW pch L=4e-08 W=2.35e-07 
M29 12 S0 14 VNW pch L=4e-08 W=2.35e-07 
M30 VDD S0 15 VNW pch L=4e-08 W=1.9e-07 
M31 13 B VDD VNW pch L=4e-08 W=2.35e-07 
.ENDS


.SUBCKT MXIT4_X0P7M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.2e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.8e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.8e-07 
M4 VSS C 5 VPW nch L=4e-08 W=1.8e-07 
M5 VSS 6 7 VPW nch L=4e-08 W=1.8e-07 
M6 8 S1 VSS VPW nch L=4e-08 W=1.8e-07 
M7 10 S1 7 VPW nch L=4e-08 W=1.8e-07 
M8 9 8 10 VPW nch L=4e-08 W=1.8e-07 
M9 Y 10 VSS VPW nch L=4e-08 W=2.2e-07 
M10 VSS 14 9 VPW nch L=4e-08 W=1.8e-07 
M11 12 A VSS VPW nch L=4e-08 W=1.8e-07 
M12 14 15 12 VPW nch L=4e-08 W=1.8e-07 
M13 13 S0 14 VPW nch L=4e-08 W=1.8e-07 
M14 VSS S0 15 VPW nch L=4e-08 W=1.2e-07 
M15 13 B VSS VPW nch L=4e-08 W=1.8e-07 
M16 VDD D 1 VNW pch L=4e-08 W=2.75e-07 
M17 4 S0 VDD VNW pch L=4e-08 W=1.9e-07 
M18 6 S0 5 VNW pch L=4e-08 W=2.75e-07 
M19 1 4 6 VNW pch L=4e-08 W=2.75e-07 
M20 VDD C 5 VNW pch L=4e-08 W=2.75e-07 
M21 VDD 6 7 VNW pch L=4e-08 W=2.05e-07 
M22 8 S1 VDD VNW pch L=4e-08 W=2.05e-07 
M23 10 S1 9 VNW pch L=4e-08 W=2.05e-07 
M24 7 8 10 VNW pch L=4e-08 W=2.05e-07 
M25 Y 10 VDD VNW pch L=4e-08 W=2.85e-07 
M26 VDD 14 9 VNW pch L=4e-08 W=2.05e-07 
M27 12 A VDD VNW pch L=4e-08 W=2.75e-07 
M28 14 15 13 VNW pch L=4e-08 W=2.75e-07 
M29 12 S0 14 VNW pch L=4e-08 W=2.75e-07 
M30 VDD S0 15 VNW pch L=4e-08 W=1.9e-07 
M31 13 B VDD VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT MXIT4_X1M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=2.1e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.2e-07 
M2 6 S0 1 VPW nch L=4e-08 W=2.1e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.1e-07 
M4 VSS C 5 VPW nch L=4e-08 W=2.1e-07 
M5 VSS 6 7 VPW nch L=4e-08 W=2.1e-07 
M6 8 S1 VSS VPW nch L=4e-08 W=2.1e-07 
M7 10 S1 7 VPW nch L=4e-08 W=2.1e-07 
M8 9 8 10 VPW nch L=4e-08 W=2.1e-07 
M9 Y 10 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 14 9 VPW nch L=4e-08 W=2.1e-07 
M11 12 A VSS VPW nch L=4e-08 W=2.1e-07 
M12 14 15 12 VPW nch L=4e-08 W=2.1e-07 
M13 13 S0 14 VPW nch L=4e-08 W=2.1e-07 
M14 VSS S0 15 VPW nch L=4e-08 W=1.2e-07 
M15 13 B VSS VPW nch L=4e-08 W=2.1e-07 
M16 VDD D 1 VNW pch L=4e-08 W=3.2e-07 
M17 4 S0 VDD VNW pch L=4e-08 W=1.9e-07 
M18 6 S0 5 VNW pch L=4e-08 W=3.2e-07 
M19 1 4 6 VNW pch L=4e-08 W=3.2e-07 
M20 VDD C 5 VNW pch L=4e-08 W=3.2e-07 
M21 VDD 6 7 VNW pch L=4e-08 W=2.4e-07 
M22 8 S1 VDD VNW pch L=4e-08 W=2.4e-07 
M23 10 S1 9 VNW pch L=4e-08 W=2.4e-07 
M24 7 8 10 VNW pch L=4e-08 W=2.4e-07 
M25 Y 10 VDD VNW pch L=4e-08 W=3.8e-07 
M26 VDD 14 9 VNW pch L=4e-08 W=2.4e-07 
M27 12 A VDD VNW pch L=4e-08 W=3.2e-07 
M28 14 15 13 VNW pch L=4e-08 W=3.2e-07 
M29 12 S0 14 VNW pch L=4e-08 W=3.2e-07 
M30 VDD S0 15 VNW pch L=4e-08 W=1.9e-07 
M31 13 B VDD VNW pch L=4e-08 W=3.2e-07 
.ENDS


.SUBCKT MXIT4_X1P4M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=2.4e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 6 S0 1 VPW nch L=4e-08 W=2.4e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.4e-07 
M4 VSS C 5 VPW nch L=4e-08 W=2.4e-07 
M5 VSS 6 7 VPW nch L=4e-08 W=2.85e-07 
M6 8 S1 VSS VPW nch L=4e-08 W=2.85e-07 
M7 10 S1 7 VPW nch L=4e-08 W=2.85e-07 
M8 9 8 10 VPW nch L=4e-08 W=2.85e-07 
M9 Y 10 VSS VPW nch L=4e-08 W=2.2e-07 
M10 VSS 10 Y VPW nch L=4e-08 W=2.2e-07 
M11 VSS 14 9 VPW nch L=4e-08 W=2.85e-07 
M12 12 A VSS VPW nch L=4e-08 W=2.4e-07 
M13 14 15 12 VPW nch L=4e-08 W=2.4e-07 
M14 13 S0 14 VPW nch L=4e-08 W=2.4e-07 
M15 VSS S0 15 VPW nch L=4e-08 W=2.4e-07 
M16 13 B VSS VPW nch L=4e-08 W=2.4e-07 
M17 VDD D 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M19 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M20 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M21 VDD C 5 VNW pch L=4e-08 W=3.8e-07 
M22 VDD 6 7 VNW pch L=4e-08 W=3.25e-07 
M23 8 S1 VDD VNW pch L=4e-08 W=3.25e-07 
M24 10 S1 9 VNW pch L=4e-08 W=3.25e-07 
M25 7 8 10 VNW pch L=4e-08 W=3.25e-07 
M26 Y 10 VDD VNW pch L=4e-08 W=2.85e-07 
M27 VDD 10 Y VNW pch L=4e-08 W=2.85e-07 
M28 VDD 14 9 VNW pch L=4e-08 W=3.25e-07 
M29 12 A VDD VNW pch L=4e-08 W=3.8e-07 
M30 14 15 13 VNW pch L=4e-08 W=3.8e-07 
M31 12 S0 14 VNW pch L=4e-08 W=3.8e-07 
M32 VDD S0 15 VNW pch L=4e-08 W=3.8e-07 
M33 13 B VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXIT4_X2M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=2.4e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 6 S0 1 VPW nch L=4e-08 W=2.4e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.4e-07 
M4 VSS C 5 VPW nch L=4e-08 W=2.4e-07 
M5 VSS 6 7 VPW nch L=4e-08 W=3.35e-07 
M6 8 S1 VSS VPW nch L=4e-08 W=3.35e-07 
M7 10 S1 7 VPW nch L=4e-08 W=3.35e-07 
M8 9 8 10 VPW nch L=4e-08 W=3.35e-07 
M9 Y 10 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 10 Y VPW nch L=4e-08 W=3.1e-07 
M11 VSS 14 9 VPW nch L=4e-08 W=3.35e-07 
M12 12 A VSS VPW nch L=4e-08 W=2.4e-07 
M13 14 15 12 VPW nch L=4e-08 W=2.4e-07 
M14 13 S0 14 VPW nch L=4e-08 W=2.4e-07 
M15 VSS S0 15 VPW nch L=4e-08 W=2.4e-07 
M16 13 B VSS VPW nch L=4e-08 W=2.4e-07 
M17 VDD D 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M19 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M20 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M21 VDD C 5 VNW pch L=4e-08 W=3.8e-07 
M22 VDD 6 7 VNW pch L=4e-08 W=3.8e-07 
M23 8 S1 VDD VNW pch L=4e-08 W=3.8e-07 
M24 10 S1 9 VNW pch L=4e-08 W=3.8e-07 
M25 7 8 10 VNW pch L=4e-08 W=3.8e-07 
M26 Y 10 VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD 10 Y VNW pch L=4e-08 W=3.8e-07 
M28 VDD 14 9 VNW pch L=4e-08 W=3.8e-07 
M29 12 A VDD VNW pch L=4e-08 W=3.8e-07 
M30 14 15 13 VNW pch L=4e-08 W=3.8e-07 
M31 12 S0 14 VNW pch L=4e-08 W=3.8e-07 
M32 VDD S0 15 VNW pch L=4e-08 W=3.8e-07 
M33 13 B VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXIT4_X3M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=2.4e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 6 S0 1 VPW nch L=4e-08 W=2.4e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.4e-07 
M4 VSS C 5 VPW nch L=4e-08 W=2.4e-07 
M5 VSS 6 7 VPW nch L=4e-08 W=3.35e-07 
M6 8 S1 VSS VPW nch L=4e-08 W=3.35e-07 
M7 10 S1 7 VPW nch L=4e-08 W=3.35e-07 
M8 9 8 10 VPW nch L=4e-08 W=3.35e-07 
M9 VSS 10 Y VPW nch L=4e-08 W=3.1e-07 
M10 Y 10 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 10 Y VPW nch L=4e-08 W=3.1e-07 
M12 VSS 14 9 VPW nch L=4e-08 W=3.35e-07 
M13 12 A VSS VPW nch L=4e-08 W=2.4e-07 
M14 14 15 12 VPW nch L=4e-08 W=2.4e-07 
M15 13 S0 14 VPW nch L=4e-08 W=2.4e-07 
M16 VSS S0 15 VPW nch L=4e-08 W=2.4e-07 
M17 13 B VSS VPW nch L=4e-08 W=2.4e-07 
M18 VDD D 1 VNW pch L=4e-08 W=3.8e-07 
M19 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M20 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M21 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M22 VDD C 5 VNW pch L=4e-08 W=3.8e-07 
M23 VDD 6 7 VNW pch L=4e-08 W=3.8e-07 
M24 8 S1 VDD VNW pch L=4e-08 W=3.8e-07 
M25 10 S1 9 VNW pch L=4e-08 W=3.8e-07 
M26 7 8 10 VNW pch L=4e-08 W=3.8e-07 
M27 VDD 10 Y VNW pch L=4e-08 W=3.8e-07 
M28 Y 10 VDD VNW pch L=4e-08 W=3.8e-07 
M29 VDD 10 Y VNW pch L=4e-08 W=3.8e-07 
M30 VDD 14 9 VNW pch L=4e-08 W=3.8e-07 
M31 12 A VDD VNW pch L=4e-08 W=3.8e-07 
M32 14 15 13 VNW pch L=4e-08 W=3.8e-07 
M33 12 S0 14 VNW pch L=4e-08 W=3.8e-07 
M34 VDD S0 15 VNW pch L=4e-08 W=3.8e-07 
M35 13 B VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXT2_X0P5B_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=1.45e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.45e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.45e-07 
M4 VSS 6 Y VPW nch L=4e-08 W=1.2e-07 
M5 5 A VSS VPW nch L=4e-08 W=1.45e-07 
M6 VDD B 1 VNW pch L=4e-08 W=2.25e-07 
M7 4 S0 VDD VNW pch L=4e-08 W=3.15e-07 
M8 6 S0 5 VNW pch L=4e-08 W=2.25e-07 
M9 1 4 6 VNW pch L=4e-08 W=2.25e-07 
M10 VDD 6 Y VNW pch L=4e-08 W=2.1e-07 
M11 5 A VDD VNW pch L=4e-08 W=2.25e-07 
.ENDS


.SUBCKT MXT2_X0P5M_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.2e-07 
M2 5 S0 1 VPW nch L=4e-08 W=1.2e-07 
M3 6 4 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS A 6 VPW nch L=4e-08 W=1.2e-07 
M5 Y 5 VSS VPW nch L=4e-08 W=1.75e-07 
M6 VDD B 1 VNW pch L=4e-08 W=1.9e-07 
M7 4 S0 VDD VNW pch L=4e-08 W=1.9e-07 
M8 5 4 1 VNW pch L=4e-08 W=1.9e-07 
M9 6 S0 5 VNW pch L=4e-08 W=1.9e-07 
M10 VDD A 6 VNW pch L=4e-08 W=1.9e-07 
M11 Y 5 VDD VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT MXT2_X0P7B_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=1.6e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.5e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.6e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.6e-07 
M4 VSS 6 Y VPW nch L=4e-08 W=1.6e-07 
M5 5 A VSS VPW nch L=4e-08 W=1.6e-07 
M6 VDD B 1 VNW pch L=4e-08 W=2.45e-07 
M7 4 S0 VDD VNW pch L=4e-08 W=3.25e-07 
M8 6 S0 5 VNW pch L=4e-08 W=2.45e-07 
M9 1 4 6 VNW pch L=4e-08 W=2.45e-07 
M10 VDD 6 Y VNW pch L=4e-08 W=2.85e-07 
M11 5 A VDD VNW pch L=4e-08 W=2.45e-07 
.ENDS


.SUBCKT MXT2_X0P7M_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=1.5e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 S0 1 VPW nch L=4e-08 W=1.5e-07 
M3 6 4 5 VPW nch L=4e-08 W=1.5e-07 
M4 VSS A 6 VPW nch L=4e-08 W=1.5e-07 
M5 Y 5 VSS VPW nch L=4e-08 W=2.45e-07 
M6 VDD B 1 VNW pch L=4e-08 W=2.25e-07 
M7 4 S0 VDD VNW pch L=4e-08 W=2.25e-07 
M8 5 4 1 VNW pch L=4e-08 W=2.25e-07 
M9 6 S0 5 VNW pch L=4e-08 W=2.25e-07 
M10 VDD A 6 VNW pch L=4e-08 W=2.25e-07 
M11 Y 5 VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT MXT2_X1B_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=1.85e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.65e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.85e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.85e-07 
M4 VSS 6 Y VPW nch L=4e-08 W=2.15e-07 
M5 5 A VSS VPW nch L=4e-08 W=1.85e-07 
M6 VDD B 1 VNW pch L=4e-08 W=2.85e-07 
M7 4 S0 VDD VNW pch L=4e-08 W=3.4e-07 
M8 6 S0 5 VNW pch L=4e-08 W=2.85e-07 
M9 1 4 6 VNW pch L=4e-08 W=2.85e-07 
M10 VDD 6 Y VNW pch L=4e-08 W=3.8e-07 
M11 5 A VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT MXT2_X1M_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=2.45e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M2 6 S0 1 VPW nch L=4e-08 W=2.45e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M4 VSS 6 Y VPW nch L=4e-08 W=3.5e-07 
M5 5 A VSS VPW nch L=4e-08 W=2.45e-07 
M6 VDD B 1 VNW pch L=4e-08 W=4e-07 
M7 4 S0 VDD VNW pch L=4e-08 W=4e-07 
M8 6 S0 5 VNW pch L=4e-08 W=4e-07 
M9 1 4 6 VNW pch L=4e-08 W=4e-07 
M10 VDD 6 Y VNW pch L=4e-08 W=3.8e-07 
M11 5 A VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXT2_X1P4B_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=2.4e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.95e-07 
M2 6 S0 1 VPW nch L=4e-08 W=2.4e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.4e-07 
M4 Y 6 VSS VPW nch L=4e-08 W=1.5e-07 
M5 VSS 6 Y VPW nch L=4e-08 W=1.5e-07 
M6 5 A VSS VPW nch L=4e-08 W=2.4e-07 
M7 VDD B 1 VNW pch L=4e-08 W=3.7e-07 
M8 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M9 6 S0 5 VNW pch L=4e-08 W=3.7e-07 
M10 1 4 6 VNW pch L=4e-08 W=3.7e-07 
M11 Y 6 VDD VNW pch L=4e-08 W=2.65e-07 
M12 VDD 6 Y VNW pch L=4e-08 W=2.65e-07 
M13 5 A VDD VNW pch L=4e-08 W=3.7e-07 
.ENDS


.SUBCKT MXT2_X1P4M_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=2.55e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.55e-07 
M2 6 S0 1 VPW nch L=4e-08 W=2.55e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.55e-07 
M4 Y 6 VSS VPW nch L=4e-08 W=2.6e-07 
M5 VSS 6 Y VPW nch L=4e-08 W=2.6e-07 
M6 5 A VSS VPW nch L=4e-08 W=2.55e-07 
M7 VDD B 1 VNW pch L=4e-08 W=4e-07 
M8 4 S0 VDD VNW pch L=4e-08 W=4e-07 
M9 6 S0 5 VNW pch L=4e-08 W=4e-07 
M10 1 4 6 VNW pch L=4e-08 W=4e-07 
M11 Y 6 VDD VNW pch L=4e-08 W=2.8e-07 
M12 VDD 6 Y VNW pch L=4e-08 W=2.8e-07 
M13 5 A VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT MXT2_X2B_A9TR Y VDD VNW VPW VSS A B S0
M0 3 B VSS VPW nch L=4e-08 W=1.45e-07 
M1 VSS B 3 VPW nch L=4e-08 W=1.45e-07 
M2 4 S0 VSS VPW nch L=4e-08 W=2.1e-07 
M3 VSS S0 4 VPW nch L=4e-08 W=2.1e-07 
M4 3 S0 5 VPW nch L=4e-08 W=1.45e-07 
M5 5 S0 3 VPW nch L=4e-08 W=1.45e-07 
M6 6 4 5 VPW nch L=4e-08 W=1.45e-07 
M7 5 4 6 VPW nch L=4e-08 W=1.45e-07 
M8 Y 5 VSS VPW nch L=4e-08 W=2.15e-07 
M9 VSS 5 Y VPW nch L=4e-08 W=2.15e-07 
M10 6 A VSS VPW nch L=4e-08 W=1.45e-07 
M11 VSS A 6 VPW nch L=4e-08 W=1.45e-07 
M12 3 B VDD VNW pch L=4e-08 W=2.25e-07 
M13 VDD B 3 VNW pch L=4e-08 W=2.25e-07 
M14 4 S0 VDD VNW pch L=4e-08 W=2.7e-07 
M15 VDD S0 4 VNW pch L=4e-08 W=2.7e-07 
M16 6 S0 5 VNW pch L=4e-08 W=2.25e-07 
M17 5 S0 6 VNW pch L=4e-08 W=2.25e-07 
M18 3 4 5 VNW pch L=4e-08 W=2.25e-07 
M19 5 4 3 VNW pch L=4e-08 W=2.25e-07 
M20 Y 5 VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M22 6 A VDD VNW pch L=4e-08 W=2.25e-07 
M23 VDD A 6 VNW pch L=4e-08 W=2.25e-07 
.ENDS


.SUBCKT MXT2_X2M_A9TR Y VDD VNW VPW VSS A B S0
M0 3 B VSS VPW nch L=4e-08 W=1.9e-07 
M1 VSS B 3 VPW nch L=4e-08 W=1.9e-07 
M2 4 S0 VSS VPW nch L=4e-08 W=1.9e-07 
M3 VSS S0 4 VPW nch L=4e-08 W=1.9e-07 
M4 6 S0 3 VPW nch L=4e-08 W=3.8e-07 
M5 5 4 6 VPW nch L=4e-08 W=3.8e-07 
M6 Y 6 VSS VPW nch L=4e-08 W=3.5e-07 
M7 VSS 6 Y VPW nch L=4e-08 W=3.5e-07 
M8 5 A VSS VPW nch L=4e-08 W=1.9e-07 
M9 VSS A 5 VPW nch L=4e-08 W=1.9e-07 
M10 3 B VDD VNW pch L=4e-08 W=3.3e-07 
M11 VDD B 3 VNW pch L=4e-08 W=3.3e-07 
M12 4 S0 VDD VNW pch L=4e-08 W=3.3e-07 
M13 VDD S0 4 VNW pch L=4e-08 W=3.3e-07 
M14 6 S0 5 VNW pch L=4e-08 W=4e-07 
M15 3 4 6 VNW pch L=4e-08 W=4e-07 
M16 Y 6 VDD VNW pch L=4e-08 W=3.8e-07 
M17 VDD 6 Y VNW pch L=4e-08 W=3.8e-07 
M18 5 A VDD VNW pch L=4e-08 W=3.3e-07 
M19 VDD A 5 VNW pch L=4e-08 W=3.3e-07 
.ENDS


.SUBCKT MXT2_X3B_A9TR Y VDD VNW VPW VSS A B S0
M0 3 B VSS VPW nch L=4e-08 W=2e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2e-07 
M2 4 S0 VSS VPW nch L=4e-08 W=2.4e-07 
M3 VSS S0 4 VPW nch L=4e-08 W=2.4e-07 
M4 3 S0 5 VPW nch L=4e-08 W=2e-07 
M5 5 S0 3 VPW nch L=4e-08 W=2e-07 
M6 6 4 5 VPW nch L=4e-08 W=2e-07 
M7 5 4 6 VPW nch L=4e-08 W=2e-07 
M8 VSS 5 Y VPW nch L=4e-08 W=2.15e-07 
M9 Y 5 VSS VPW nch L=4e-08 W=2.15e-07 
M10 VSS 5 Y VPW nch L=4e-08 W=2.15e-07 
M11 6 A VSS VPW nch L=4e-08 W=2e-07 
M12 VSS A 6 VPW nch L=4e-08 W=2e-07 
M13 3 B VDD VNW pch L=4e-08 W=3.1e-07 
M14 VDD B 3 VNW pch L=4e-08 W=3.1e-07 
M15 4 S0 VDD VNW pch L=4e-08 W=3.1e-07 
M16 VDD S0 4 VNW pch L=4e-08 W=3.1e-07 
M17 6 S0 5 VNW pch L=4e-08 W=3.1e-07 
M18 5 S0 6 VNW pch L=4e-08 W=3.1e-07 
M19 3 4 5 VNW pch L=4e-08 W=3.1e-07 
M20 5 4 3 VNW pch L=4e-08 W=3.1e-07 
M21 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M22 Y 5 VDD VNW pch L=4e-08 W=3.8e-07 
M23 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M24 6 A VDD VNW pch L=4e-08 W=3.1e-07 
M25 VDD A 6 VNW pch L=4e-08 W=3.1e-07 
.ENDS


.SUBCKT MXT2_X3M_A9TR Y VDD VNW VPW VSS A B S0
M0 3 B VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.45e-07 
M2 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M3 VSS S0 4 VPW nch L=4e-08 W=2.45e-07 
M4 3 S0 5 VPW nch L=4e-08 W=2.45e-07 
M5 5 S0 3 VPW nch L=4e-08 W=2.45e-07 
M6 6 4 5 VPW nch L=4e-08 W=2.45e-07 
M7 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M8 VSS 5 Y VPW nch L=4e-08 W=3.5e-07 
M9 Y 5 VSS VPW nch L=4e-08 W=3.5e-07 
M10 VSS 5 Y VPW nch L=4e-08 W=3.5e-07 
M11 6 A VSS VPW nch L=4e-08 W=2.45e-07 
M12 VSS A 6 VPW nch L=4e-08 W=2.45e-07 
M13 3 B VDD VNW pch L=4e-08 W=3.8e-07 
M14 VDD B 3 VNW pch L=4e-08 W=3.8e-07 
M15 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M16 VDD S0 4 VNW pch L=4e-08 W=3.8e-07 
M17 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M18 5 S0 6 VNW pch L=4e-08 W=3.8e-07 
M19 3 4 5 VNW pch L=4e-08 W=3.8e-07 
M20 5 4 3 VNW pch L=4e-08 W=3.8e-07 
M21 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M22 Y 5 VDD VNW pch L=4e-08 W=3.8e-07 
M23 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M24 6 A VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD A 6 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXT2_X4B_A9TR Y VDD VNW VPW VSS A B S0
M0 1 B VSS VPW nch L=4e-08 W=2.65e-07 
M1 VSS B 1 VPW nch L=4e-08 W=2.65e-07 
M2 4 S0 VSS VPW nch L=4e-08 W=2.75e-07 
M3 VSS S0 4 VPW nch L=4e-08 W=2.75e-07 
M4 1 S0 6 VPW nch L=4e-08 W=2.65e-07 
M5 6 S0 1 VPW nch L=4e-08 W=2.65e-07 
M6 5 4 6 VPW nch L=4e-08 W=2.65e-07 
M7 6 4 5 VPW nch L=4e-08 W=2.65e-07 
M8 Y 6 VSS VPW nch L=4e-08 W=2.85e-07 
M9 VSS 6 Y VPW nch L=4e-08 W=2.85e-07 
M10 Y 6 VSS VPW nch L=4e-08 W=2.85e-07 
M11 VSS A 5 VPW nch L=4e-08 W=2.65e-07 
M12 5 A VSS VPW nch L=4e-08 W=2.65e-07 
M13 VDD B 1 VNW pch L=4e-08 W=2.75e-07 
M14 1 B VDD VNW pch L=4e-08 W=2.75e-07 
M15 VDD B 1 VNW pch L=4e-08 W=2.75e-07 
M16 4 S0 VDD VNW pch L=4e-08 W=3.55e-07 
M17 VDD S0 4 VNW pch L=4e-08 W=3.55e-07 
M18 6 S0 5 VNW pch L=4e-08 W=2.75e-07 
M19 5 S0 6 VNW pch L=4e-08 W=2.75e-07 
M20 6 S0 5 VNW pch L=4e-08 W=2.75e-07 
M21 1 4 6 VNW pch L=4e-08 W=2.75e-07 
M22 6 4 1 VNW pch L=4e-08 W=2.75e-07 
M23 1 4 6 VNW pch L=4e-08 W=2.75e-07 
M24 Y 6 VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD 6 Y VNW pch L=4e-08 W=3.8e-07 
M26 Y 6 VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD 6 Y VNW pch L=4e-08 W=3.8e-07 
M28 5 A VDD VNW pch L=4e-08 W=2.75e-07 
M29 VDD A 5 VNW pch L=4e-08 W=2.75e-07 
M30 5 A VDD VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT MXT2_X4M_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 1 VPW nch L=4e-08 W=2.45e-07 
M1 1 B VSS VPW nch L=4e-08 W=2.45e-07 
M2 VSS B 1 VPW nch L=4e-08 W=2.45e-07 
M3 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M4 VSS S0 4 VPW nch L=4e-08 W=2.45e-07 
M5 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M6 6 S0 1 VPW nch L=4e-08 W=2.45e-07 
M7 1 S0 6 VPW nch L=4e-08 W=2.45e-07 
M8 6 S0 1 VPW nch L=4e-08 W=2.45e-07 
M9 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M10 6 4 5 VPW nch L=4e-08 W=2.45e-07 
M11 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M12 Y 6 VSS VPW nch L=4e-08 W=3.5e-07 
M13 VSS 6 Y VPW nch L=4e-08 W=3.5e-07 
M14 Y 6 VSS VPW nch L=4e-08 W=3.5e-07 
M15 VSS 6 Y VPW nch L=4e-08 W=3.5e-07 
M16 5 A VSS VPW nch L=4e-08 W=2.45e-07 
M17 VSS A 5 VPW nch L=4e-08 W=2.45e-07 
M18 5 A VSS VPW nch L=4e-08 W=2.45e-07 
M19 VDD B 1 VNW pch L=4e-08 W=3.8e-07 
M20 1 B VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD B 1 VNW pch L=4e-08 W=3.8e-07 
M22 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M23 VDD S0 4 VNW pch L=4e-08 W=3.8e-07 
M24 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M25 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M26 5 S0 6 VNW pch L=4e-08 W=3.8e-07 
M27 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M28 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M29 6 4 1 VNW pch L=4e-08 W=3.8e-07 
M30 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M31 Y 6 VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD 6 Y VNW pch L=4e-08 W=3.8e-07 
M33 Y 6 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 6 Y VNW pch L=4e-08 W=3.8e-07 
M35 5 A VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD A 5 VNW pch L=4e-08 W=3.8e-07 
M37 5 A VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXT2_X6B_A9TR Y VDD VNW VPW VSS A B S0
M0 VSS B 2 VPW nch L=4e-08 W=2.6e-07 
M1 2 B VSS VPW nch L=4e-08 W=2.6e-07 
M2 VSS B 2 VPW nch L=4e-08 W=2.6e-07 
M3 4 S0 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS S0 4 VPW nch L=4e-08 W=3.1e-07 
M5 4 S0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 5 S0 2 VPW nch L=4e-08 W=2.6e-07 
M7 2 S0 5 VPW nch L=4e-08 W=2.6e-07 
M8 5 S0 2 VPW nch L=4e-08 W=2.6e-07 
M9 6 4 5 VPW nch L=4e-08 W=2.6e-07 
M10 5 4 6 VPW nch L=4e-08 W=2.6e-07 
M11 6 4 5 VPW nch L=4e-08 W=2.6e-07 
M12 Y 5 VSS VPW nch L=4e-08 W=3.25e-07 
M13 VSS 5 Y VPW nch L=4e-08 W=3.25e-07 
M14 Y 5 VSS VPW nch L=4e-08 W=3.25e-07 
M15 VSS 5 Y VPW nch L=4e-08 W=3.25e-07 
M16 VSS A 6 VPW nch L=4e-08 W=2.6e-07 
M17 6 A VSS VPW nch L=4e-08 W=2.6e-07 
M18 VSS A 6 VPW nch L=4e-08 W=2.6e-07 
M19 2 B VDD VNW pch L=4e-08 W=3e-07 
M20 VDD B 2 VNW pch L=4e-08 W=3e-07 
M21 2 B VDD VNW pch L=4e-08 W=3e-07 
M22 VDD B 2 VNW pch L=4e-08 W=3e-07 
M23 4 S0 VDD VNW pch L=4e-08 W=3e-07 
M24 VDD S0 4 VNW pch L=4e-08 W=3e-07 
M25 4 S0 VDD VNW pch L=4e-08 W=3e-07 
M26 VDD S0 4 VNW pch L=4e-08 W=3e-07 
M27 6 S0 5 VNW pch L=4e-08 W=3e-07 
M28 5 S0 6 VNW pch L=4e-08 W=3e-07 
M29 6 S0 5 VNW pch L=4e-08 W=3e-07 
M30 5 S0 6 VNW pch L=4e-08 W=3e-07 
M31 2 4 5 VNW pch L=4e-08 W=3e-07 
M32 5 4 2 VNW pch L=4e-08 W=3e-07 
M33 2 4 5 VNW pch L=4e-08 W=3e-07 
M34 5 4 2 VNW pch L=4e-08 W=3e-07 
M35 Y 5 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M37 Y 5 VDD VNW pch L=4e-08 W=3.8e-07 
M38 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M39 Y 5 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M41 6 A VDD VNW pch L=4e-08 W=3e-07 
M42 VDD A 6 VNW pch L=4e-08 W=3e-07 
M43 6 A VDD VNW pch L=4e-08 W=3e-07 
M44 VDD A 6 VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT MXT2_X6M_A9TR Y VDD VNW VPW VSS A B S0
M0 3 B VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.45e-07 
M2 3 B VSS VPW nch L=4e-08 W=2.45e-07 
M3 VSS B 3 VPW nch L=4e-08 W=2.45e-07 
M4 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M5 VSS S0 4 VPW nch L=4e-08 W=2.45e-07 
M6 4 S0 VSS VPW nch L=4e-08 W=2.45e-07 
M7 VSS S0 4 VPW nch L=4e-08 W=2.45e-07 
M8 3 S0 5 VPW nch L=4e-08 W=2.45e-07 
M9 5 S0 3 VPW nch L=4e-08 W=2.45e-07 
M10 3 S0 5 VPW nch L=4e-08 W=2.45e-07 
M11 5 S0 3 VPW nch L=4e-08 W=2.45e-07 
M12 6 4 5 VPW nch L=4e-08 W=2.45e-07 
M13 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M14 6 4 5 VPW nch L=4e-08 W=2.45e-07 
M15 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M16 Y 5 VSS VPW nch L=4e-08 W=3.5e-07 
M17 VSS 5 Y VPW nch L=4e-08 W=3.5e-07 
M18 Y 5 VSS VPW nch L=4e-08 W=3.5e-07 
M19 VSS 5 Y VPW nch L=4e-08 W=3.5e-07 
M20 Y 5 VSS VPW nch L=4e-08 W=3.5e-07 
M21 VSS 5 Y VPW nch L=4e-08 W=3.5e-07 
M22 6 A VSS VPW nch L=4e-08 W=2.45e-07 
M23 VSS A 6 VPW nch L=4e-08 W=2.45e-07 
M24 6 A VSS VPW nch L=4e-08 W=2.45e-07 
M25 VSS A 6 VPW nch L=4e-08 W=2.45e-07 
M26 3 B VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD B 3 VNW pch L=4e-08 W=3.8e-07 
M28 3 B VDD VNW pch L=4e-08 W=3.8e-07 
M29 VDD B 3 VNW pch L=4e-08 W=3.8e-07 
M30 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD S0 4 VNW pch L=4e-08 W=3.8e-07 
M32 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD S0 4 VNW pch L=4e-08 W=3.8e-07 
M34 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M35 5 S0 6 VNW pch L=4e-08 W=3.8e-07 
M36 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M37 5 S0 6 VNW pch L=4e-08 W=3.8e-07 
M38 3 4 5 VNW pch L=4e-08 W=3.8e-07 
M39 5 4 3 VNW pch L=4e-08 W=3.8e-07 
M40 3 4 5 VNW pch L=4e-08 W=3.8e-07 
M41 5 4 3 VNW pch L=4e-08 W=3.8e-07 
M42 Y 5 VDD VNW pch L=4e-08 W=3.8e-07 
M43 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M44 Y 5 VDD VNW pch L=4e-08 W=3.8e-07 
M45 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M46 Y 5 VDD VNW pch L=4e-08 W=3.8e-07 
M47 VDD 5 Y VNW pch L=4e-08 W=3.8e-07 
M48 6 A VDD VNW pch L=4e-08 W=3.8e-07 
M49 VDD A 6 VNW pch L=4e-08 W=3.8e-07 
M50 6 A VDD VNW pch L=4e-08 W=3.8e-07 
M51 VDD A 6 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXT4_X0P5M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=1.5e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.5e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.5e-07 
M4 VSS C 5 VPW nch L=4e-08 W=1.5e-07 
M5 7 S1 VSS VPW nch L=4e-08 W=1.5e-07 
M6 9 S1 6 VPW nch L=4e-08 W=1.5e-07 
M7 8 7 9 VPW nch L=4e-08 W=1.5e-07 
M8 Y 9 VSS VPW nch L=4e-08 W=1.8e-07 
M9 11 A VSS VPW nch L=4e-08 W=1.5e-07 
M10 8 13 11 VPW nch L=4e-08 W=1.5e-07 
M11 12 S0 8 VPW nch L=4e-08 W=1.5e-07 
M12 VSS S0 13 VPW nch L=4e-08 W=2e-07 
M13 12 B VSS VPW nch L=4e-08 W=1.5e-07 
M14 VDD D 1 VNW pch L=4e-08 W=2.8e-07 
M15 4 S0 VDD VNW pch L=4e-08 W=2.65e-07 
M16 6 S0 5 VNW pch L=4e-08 W=2.8e-07 
M17 1 4 6 VNW pch L=4e-08 W=2.8e-07 
M18 VDD C 5 VNW pch L=4e-08 W=2.8e-07 
M19 7 S1 VDD VNW pch L=4e-08 W=2.8e-07 
M20 9 S1 8 VNW pch L=4e-08 W=2.8e-07 
M21 6 7 9 VNW pch L=4e-08 W=2.8e-07 
M22 Y 9 VDD VNW pch L=4e-08 W=2e-07 
M23 11 A VDD VNW pch L=4e-08 W=2.8e-07 
M24 8 13 12 VNW pch L=4e-08 W=2.8e-07 
M25 11 S0 8 VNW pch L=4e-08 W=2.8e-07 
M26 VDD S0 13 VNW pch L=4e-08 W=2.65e-07 
M27 12 B VDD VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT MXT4_X0P7M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=1.75e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2e-07 
M2 6 S0 1 VPW nch L=4e-08 W=1.75e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.75e-07 
M4 VSS C 5 VPW nch L=4e-08 W=1.75e-07 
M5 7 S1 VSS VPW nch L=4e-08 W=1.75e-07 
M6 9 S1 6 VPW nch L=4e-08 W=1.75e-07 
M7 8 7 9 VPW nch L=4e-08 W=1.75e-07 
M8 Y 9 VSS VPW nch L=4e-08 W=2.6e-07 
M9 11 A VSS VPW nch L=4e-08 W=1.75e-07 
M10 8 13 11 VPW nch L=4e-08 W=1.75e-07 
M11 12 S0 8 VPW nch L=4e-08 W=1.75e-07 
M12 VSS S0 13 VPW nch L=4e-08 W=2e-07 
M13 12 B VSS VPW nch L=4e-08 W=1.75e-07 
M14 VDD D 1 VNW pch L=4e-08 W=3.25e-07 
M15 4 S0 VDD VNW pch L=4e-08 W=2.65e-07 
M16 6 S0 5 VNW pch L=4e-08 W=3.25e-07 
M17 1 4 6 VNW pch L=4e-08 W=3.25e-07 
M18 VDD C 5 VNW pch L=4e-08 W=3.25e-07 
M19 7 S1 VDD VNW pch L=4e-08 W=3.25e-07 
M20 9 S1 8 VNW pch L=4e-08 W=3.25e-07 
M21 6 7 9 VNW pch L=4e-08 W=3.25e-07 
M22 Y 9 VDD VNW pch L=4e-08 W=2.85e-07 
M23 11 A VDD VNW pch L=4e-08 W=3.25e-07 
M24 8 13 12 VNW pch L=4e-08 W=3.25e-07 
M25 11 S0 8 VNW pch L=4e-08 W=3.25e-07 
M26 VDD S0 13 VNW pch L=4e-08 W=2.65e-07 
M27 12 B VDD VNW pch L=4e-08 W=3.25e-07 
.ENDS


.SUBCKT MXT4_X1M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=2.05e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.3e-07 
M2 6 S0 1 VPW nch L=4e-08 W=2.05e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.05e-07 
M4 VSS C 5 VPW nch L=4e-08 W=2.05e-07 
M5 7 S1 VSS VPW nch L=4e-08 W=2.05e-07 
M6 9 S1 6 VPW nch L=4e-08 W=2.05e-07 
M7 8 7 9 VPW nch L=4e-08 W=2.05e-07 
M8 Y 9 VSS VPW nch L=4e-08 W=3.1e-07 
M9 11 A VSS VPW nch L=4e-08 W=2.05e-07 
M10 8 13 11 VPW nch L=4e-08 W=2.05e-07 
M11 12 S0 8 VPW nch L=4e-08 W=2.05e-07 
M12 VSS S0 13 VPW nch L=4e-08 W=2.3e-07 
M13 12 B VSS VPW nch L=4e-08 W=2.05e-07 
M14 VDD D 1 VNW pch L=4e-08 W=3.8e-07 
M15 4 S0 VDD VNW pch L=4e-08 W=3.05e-07 
M16 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M17 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M18 VDD C 5 VNW pch L=4e-08 W=3.8e-07 
M19 7 S1 VDD VNW pch L=4e-08 W=3.8e-07 
M20 9 S1 8 VNW pch L=4e-08 W=3.8e-07 
M21 6 7 9 VNW pch L=4e-08 W=3.8e-07 
M22 Y 9 VDD VNW pch L=4e-08 W=3.8e-07 
M23 11 A VDD VNW pch L=4e-08 W=3.8e-07 
M24 8 13 12 VNW pch L=4e-08 W=3.8e-07 
M25 11 S0 8 VNW pch L=4e-08 W=3.8e-07 
M26 VDD S0 13 VNW pch L=4e-08 W=3.05e-07 
M27 12 B VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXT4_X1P4M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 VSS D 1 VPW nch L=4e-08 W=2.05e-07 
M1 4 S0 VSS VPW nch L=4e-08 W=2.3e-07 
M2 6 S0 1 VPW nch L=4e-08 W=2.05e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.05e-07 
M4 VSS C 5 VPW nch L=4e-08 W=2.05e-07 
M5 7 S1 VSS VPW nch L=4e-08 W=2.05e-07 
M6 9 S1 6 VPW nch L=4e-08 W=2.05e-07 
M7 8 7 9 VPW nch L=4e-08 W=2.05e-07 
M8 Y 9 VSS VPW nch L=4e-08 W=2.6e-07 
M9 VSS 9 Y VPW nch L=4e-08 W=2.6e-07 
M10 11 A VSS VPW nch L=4e-08 W=2.05e-07 
M11 8 13 11 VPW nch L=4e-08 W=2.05e-07 
M12 12 S0 8 VPW nch L=4e-08 W=2.05e-07 
M13 VSS S0 13 VPW nch L=4e-08 W=2.3e-07 
M14 12 B VSS VPW nch L=4e-08 W=2.05e-07 
M15 VDD D 1 VNW pch L=4e-08 W=3.8e-07 
M16 4 S0 VDD VNW pch L=4e-08 W=3.05e-07 
M17 6 S0 5 VNW pch L=4e-08 W=4e-07 
M18 1 4 6 VNW pch L=4e-08 W=4e-07 
M19 VDD C 5 VNW pch L=4e-08 W=3.8e-07 
M20 7 S1 VDD VNW pch L=4e-08 W=3.8e-07 
M21 9 S1 8 VNW pch L=4e-08 W=4e-07 
M22 6 7 9 VNW pch L=4e-08 W=4e-07 
M23 Y 9 VDD VNW pch L=4e-08 W=2.85e-07 
M24 VDD 9 Y VNW pch L=4e-08 W=2.85e-07 
M25 11 A VDD VNW pch L=4e-08 W=3.8e-07 
M26 8 13 12 VNW pch L=4e-08 W=4e-07 
M27 11 S0 8 VNW pch L=4e-08 W=4e-07 
M28 VDD S0 13 VNW pch L=4e-08 W=3.05e-07 
M29 12 B VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXT4_X2M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 3 D VSS VPW nch L=4e-08 W=2.05e-07 
M1 VSS D 3 VPW nch L=4e-08 W=2.05e-07 
M2 4 S0 VSS VPW nch L=4e-08 W=2.95e-07 
M3 3 S0 5 VPW nch L=4e-08 W=2.05e-07 
M4 5 S0 3 VPW nch L=4e-08 W=2.05e-07 
M5 6 4 5 VPW nch L=4e-08 W=2.05e-07 
M6 5 4 6 VPW nch L=4e-08 W=2.05e-07 
M7 6 C VSS VPW nch L=4e-08 W=2.05e-07 
M8 VSS C 6 VPW nch L=4e-08 W=2.05e-07 
M9 7 S1 VSS VPW nch L=4e-08 W=2.05e-07 
M10 VSS S1 7 VPW nch L=4e-08 W=2.05e-07 
M11 5 S1 8 VPW nch L=4e-08 W=2.05e-07 
M12 8 S1 5 VPW nch L=4e-08 W=2.05e-07 
M13 9 7 8 VPW nch L=4e-08 W=2.05e-07 
M14 8 7 9 VPW nch L=4e-08 W=2.05e-07 
M15 Y 8 VSS VPW nch L=4e-08 W=3.5e-07 
M16 VSS 8 Y VPW nch L=4e-08 W=3.5e-07 
M17 11 A VSS VPW nch L=4e-08 W=2.05e-07 
M18 VSS A 11 VPW nch L=4e-08 W=2.05e-07 
M19 11 13 9 VPW nch L=4e-08 W=2.05e-07 
M20 9 13 11 VPW nch L=4e-08 W=2.05e-07 
M21 12 S0 9 VPW nch L=4e-08 W=2.05e-07 
M22 9 S0 12 VPW nch L=4e-08 W=2.05e-07 
M23 VSS S0 13 VPW nch L=4e-08 W=2.95e-07 
M24 12 B VSS VPW nch L=4e-08 W=2.05e-07 
M25 VSS B 12 VPW nch L=4e-08 W=2.05e-07 
M26 3 D VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD D 3 VNW pch L=4e-08 W=3.8e-07 
M28 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M29 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M30 5 S0 6 VNW pch L=4e-08 W=3.8e-07 
M31 3 4 5 VNW pch L=4e-08 W=3.8e-07 
M32 5 4 3 VNW pch L=4e-08 W=3.8e-07 
M33 6 C VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD C 6 VNW pch L=4e-08 W=3.8e-07 
M35 7 S1 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD S1 7 VNW pch L=4e-08 W=3.8e-07 
M37 9 S1 8 VNW pch L=4e-08 W=3.8e-07 
M38 8 S1 9 VNW pch L=4e-08 W=3.8e-07 
M39 5 7 8 VNW pch L=4e-08 W=3.8e-07 
M40 8 7 5 VNW pch L=4e-08 W=3.8e-07 
M41 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M42 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
M43 11 A VDD VNW pch L=4e-08 W=3.8e-07 
M44 VDD A 11 VNW pch L=4e-08 W=3.8e-07 
M45 12 13 9 VNW pch L=4e-08 W=3.8e-07 
M46 9 13 12 VNW pch L=4e-08 W=3.8e-07 
M47 11 S0 9 VNW pch L=4e-08 W=3.8e-07 
M48 9 S0 11 VNW pch L=4e-08 W=3.8e-07 
M49 VDD S0 13 VNW pch L=4e-08 W=3.8e-07 
M50 12 B VDD VNW pch L=4e-08 W=3.8e-07 
M51 VDD B 12 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT MXT4_X3M_A9TR Y VDD VNW VPW VSS A B C D S0 S1
M0 3 D VSS VPW nch L=4e-08 W=2.05e-07 
M1 VSS D 3 VPW nch L=4e-08 W=2.05e-07 
M2 4 S0 VSS VPW nch L=4e-08 W=2.95e-07 
M3 3 S0 5 VPW nch L=4e-08 W=2.05e-07 
M4 5 S0 3 VPW nch L=4e-08 W=2.05e-07 
M5 6 4 5 VPW nch L=4e-08 W=2.05e-07 
M6 5 4 6 VPW nch L=4e-08 W=2.05e-07 
M7 6 C VSS VPW nch L=4e-08 W=2.05e-07 
M8 VSS C 6 VPW nch L=4e-08 W=2.05e-07 
M9 7 S1 VSS VPW nch L=4e-08 W=2.05e-07 
M10 VSS S1 7 VPW nch L=4e-08 W=2.05e-07 
M11 5 S1 8 VPW nch L=4e-08 W=2.05e-07 
M12 8 S1 5 VPW nch L=4e-08 W=2.05e-07 
M13 9 7 8 VPW nch L=4e-08 W=2.05e-07 
M14 8 7 9 VPW nch L=4e-08 W=2.05e-07 
M15 VSS 8 Y VPW nch L=4e-08 W=3.5e-07 
M16 Y 8 VSS VPW nch L=4e-08 W=3.5e-07 
M17 VSS 8 Y VPW nch L=4e-08 W=3.5e-07 
M18 11 A VSS VPW nch L=4e-08 W=2.05e-07 
M19 VSS A 11 VPW nch L=4e-08 W=2.05e-07 
M20 11 13 9 VPW nch L=4e-08 W=2.05e-07 
M21 9 13 11 VPW nch L=4e-08 W=2.05e-07 
M22 12 S0 9 VPW nch L=4e-08 W=2.05e-07 
M23 9 S0 12 VPW nch L=4e-08 W=2.05e-07 
M24 VSS S0 13 VPW nch L=4e-08 W=2.95e-07 
M25 12 B VSS VPW nch L=4e-08 W=2.05e-07 
M26 VSS B 12 VPW nch L=4e-08 W=2.05e-07 
M27 3 D VDD VNW pch L=4e-08 W=3.8e-07 
M28 VDD D 3 VNW pch L=4e-08 W=3.8e-07 
M29 4 S0 VDD VNW pch L=4e-08 W=3.8e-07 
M30 6 S0 5 VNW pch L=4e-08 W=3.8e-07 
M31 5 S0 6 VNW pch L=4e-08 W=3.8e-07 
M32 3 4 5 VNW pch L=4e-08 W=3.8e-07 
M33 5 4 3 VNW pch L=4e-08 W=3.8e-07 
M34 6 C VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD C 6 VNW pch L=4e-08 W=3.8e-07 
M36 7 S1 VDD VNW pch L=4e-08 W=3.8e-07 
M37 VDD S1 7 VNW pch L=4e-08 W=3.8e-07 
M38 9 S1 8 VNW pch L=4e-08 W=3.8e-07 
M39 8 S1 9 VNW pch L=4e-08 W=3.8e-07 
M40 5 7 8 VNW pch L=4e-08 W=3.8e-07 
M41 8 7 5 VNW pch L=4e-08 W=3.8e-07 
M42 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
M43 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M44 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
M45 11 A VDD VNW pch L=4e-08 W=3.8e-07 
M46 VDD A 11 VNW pch L=4e-08 W=3.8e-07 
M47 12 13 9 VNW pch L=4e-08 W=3.8e-07 
M48 9 13 12 VNW pch L=4e-08 W=3.8e-07 
M49 11 S0 9 VNW pch L=4e-08 W=3.8e-07 
M50 9 S0 11 VNW pch L=4e-08 W=3.8e-07 
M51 VDD S0 13 VNW pch L=4e-08 W=3.8e-07 
M52 12 B VDD VNW pch L=4e-08 W=3.8e-07 
M53 VDD B 12 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT NAND2B_X0P5M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 7 B VSS VPW nch L=4e-08 W=2e-07 
M2 Y 1 7 VPW nch L=4e-08 W=2e-07 
M3 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M4 Y B VDD VNW pch L=4e-08 W=1.7e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=1.7e-07 
.ENDS


.SUBCKT NAND2B_X0P7M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 7 B VSS VPW nch L=4e-08 W=2.85e-07 
M2 Y 1 7 VPW nch L=4e-08 W=2.85e-07 
M3 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M4 Y B VDD VNW pch L=4e-08 W=2.45e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=2.45e-07 
.ENDS


.SUBCKT NAND2B_X1M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 7 B VSS VPW nch L=4e-08 W=4e-07 
M2 Y 1 7 VPW nch L=4e-08 W=4e-07 
M3 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M4 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M5 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2B_X1P4M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.4e-07 
M1 7 B VSS VPW nch L=4e-08 W=2.85e-07 
M2 Y 1 7 VPW nch L=4e-08 W=2.85e-07 
M3 8 1 Y VPW nch L=4e-08 W=2.85e-07 
M4 VSS B 8 VPW nch L=4e-08 W=2.85e-07 
M5 VDD AN 1 VNW pch L=4e-08 W=1.8e-07 
M6 Y B VDD VNW pch L=4e-08 W=2.45e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=2.45e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=2.45e-07 
M9 VDD B Y VNW pch L=4e-08 W=2.45e-07 
.ENDS


.SUBCKT NAND2B_X2M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.85e-07 
M1 7 B VSS VPW nch L=4e-08 W=3.65e-07 
M2 Y 1 7 VPW nch L=4e-08 W=3.65e-07 
M3 8 1 Y VPW nch L=4e-08 W=4e-07 
M4 VSS B 8 VPW nch L=4e-08 W=4e-07 
M5 VDD AN 1 VNW pch L=4e-08 W=2.4e-07 
M6 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M9 VDD B Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2B_X3M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=2.75e-07 
M1 7 B VSS VPW nch L=4e-08 W=3.65e-07 
M2 Y 1 7 VPW nch L=4e-08 W=3.65e-07 
M3 8 1 Y VPW nch L=4e-08 W=4e-07 
M4 VSS B 8 VPW nch L=4e-08 W=4e-07 
M5 9 B VSS VPW nch L=4e-08 W=4e-07 
M6 Y 1 9 VPW nch L=4e-08 W=4e-07 
M7 VDD AN 1 VNW pch L=4e-08 W=3.5e-07 
M8 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M10 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M11 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M12 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M13 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2B_X4M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 2 VPW nch L=4e-08 W=3.7e-07 
M1 8 B VSS VPW nch L=4e-08 W=4e-07 
M2 Y 2 8 VPW nch L=4e-08 W=4e-07 
M3 9 2 Y VPW nch L=4e-08 W=4e-07 
M4 VSS B 9 VPW nch L=4e-08 W=4e-07 
M5 10 B VSS VPW nch L=4e-08 W=4e-07 
M6 Y 2 10 VPW nch L=4e-08 W=4e-07 
M7 11 2 Y VPW nch L=4e-08 W=4e-07 
M8 VSS B 11 VPW nch L=4e-08 W=4e-07 
M9 2 AN VDD VNW pch L=4e-08 W=2.35e-07 
M10 VDD AN 2 VNW pch L=4e-08 W=2.35e-07 
M11 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M12 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M13 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M14 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M15 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M16 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M17 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M18 VDD B Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2B_X6M_A9TR Y VDD VNW VPW VSS AN B
M0 3 AN VSS VPW nch L=4e-08 W=2.75e-07 
M1 VSS AN 3 VPW nch L=4e-08 W=2.75e-07 
M2 7 B VSS VPW nch L=4e-08 W=4e-07 
M3 Y 3 7 VPW nch L=4e-08 W=4e-07 
M4 8 3 Y VPW nch L=4e-08 W=4e-07 
M5 VSS B 8 VPW nch L=4e-08 W=4e-07 
M6 9 B VSS VPW nch L=4e-08 W=4e-07 
M7 Y 3 9 VPW nch L=4e-08 W=4e-07 
M8 10 3 Y VPW nch L=4e-08 W=4e-07 
M9 VSS B 10 VPW nch L=4e-08 W=4e-07 
M10 11 B VSS VPW nch L=4e-08 W=4e-07 
M11 Y 3 11 VPW nch L=4e-08 W=4e-07 
M12 12 3 Y VPW nch L=4e-08 W=4e-07 
M13 VSS B 12 VPW nch L=4e-08 W=4e-07 
M14 3 AN VDD VNW pch L=4e-08 W=3.5e-07 
M15 VDD AN 3 VNW pch L=4e-08 W=3.5e-07 
M16 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M17 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M18 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M19 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M20 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M21 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M22 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M23 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M24 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M25 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M26 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M27 VDD B Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2B_X8M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=2.45e-07 
M1 1 AN VSS VPW nch L=4e-08 W=2.45e-07 
M2 VSS AN 1 VPW nch L=4e-08 W=2.45e-07 
M3 7 B VSS VPW nch L=4e-08 W=4e-07 
M4 Y 1 7 VPW nch L=4e-08 W=4e-07 
M5 8 1 Y VPW nch L=4e-08 W=4e-07 
M6 VSS B 8 VPW nch L=4e-08 W=4e-07 
M7 9 B VSS VPW nch L=4e-08 W=4e-07 
M8 Y 1 9 VPW nch L=4e-08 W=4e-07 
M9 10 1 Y VPW nch L=4e-08 W=4e-07 
M10 VSS B 10 VPW nch L=4e-08 W=4e-07 
M11 11 B VSS VPW nch L=4e-08 W=4e-07 
M12 Y 1 11 VPW nch L=4e-08 W=4e-07 
M13 12 1 Y VPW nch L=4e-08 W=4e-07 
M14 VSS B 12 VPW nch L=4e-08 W=4e-07 
M15 13 B VSS VPW nch L=4e-08 W=4e-07 
M16 Y 1 13 VPW nch L=4e-08 W=4e-07 
M17 14 1 Y VPW nch L=4e-08 W=4e-07 
M18 VSS B 14 VPW nch L=4e-08 W=4e-07 
M19 VDD AN 1 VNW pch L=4e-08 W=3.15e-07 
M20 1 AN VDD VNW pch L=4e-08 W=3.15e-07 
M21 VDD AN 1 VNW pch L=4e-08 W=3.15e-07 
M22 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M23 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M24 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M25 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M26 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M27 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M28 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M29 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M30 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M31 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M32 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M33 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M34 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M35 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M36 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M37 VDD B Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2XB_X0P5M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.2e-07 
M1 7 1 VSS VPW nch L=4e-08 W=2e-07 
M2 Y A 7 VPW nch L=4e-08 W=2e-07 
M3 VDD BN 1 VNW pch L=4e-08 W=1.55e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=1.7e-07 
M5 VDD A Y VNW pch L=4e-08 W=1.7e-07 
.ENDS


.SUBCKT NAND2XB_X0P7M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.2e-07 
M1 7 1 VSS VPW nch L=4e-08 W=2.85e-07 
M2 Y A 7 VPW nch L=4e-08 W=2.85e-07 
M3 VDD BN 1 VNW pch L=4e-08 W=1.55e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=2.45e-07 
M5 VDD A Y VNW pch L=4e-08 W=2.45e-07 
.ENDS


.SUBCKT NAND2XB_X1M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.2e-07 
M1 7 1 VSS VPW nch L=4e-08 W=4e-07 
M2 Y A 7 VPW nch L=4e-08 W=4e-07 
M3 VDD BN 1 VNW pch L=4e-08 W=1.55e-07 
M4 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M5 VDD A Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2XB_X1P4M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.4e-07 
M1 7 1 VSS VPW nch L=4e-08 W=2.85e-07 
M2 Y A 7 VPW nch L=4e-08 W=2.85e-07 
M3 8 A Y VPW nch L=4e-08 W=2.85e-07 
M4 VSS 1 8 VPW nch L=4e-08 W=2.85e-07 
M5 VDD BN 1 VNW pch L=4e-08 W=1.8e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=2.45e-07 
M7 VDD A Y VNW pch L=4e-08 W=2.45e-07 
M8 Y A VDD VNW pch L=4e-08 W=2.45e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=2.45e-07 
.ENDS


.SUBCKT NAND2XB_X2M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.85e-07 
M1 7 1 VSS VPW nch L=4e-08 W=4e-07 
M2 Y A 7 VPW nch L=4e-08 W=4e-07 
M3 8 A Y VPW nch L=4e-08 W=4e-07 
M4 VSS 1 8 VPW nch L=4e-08 W=4e-07 
M5 VDD BN 1 VNW pch L=4e-08 W=2.4e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M7 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M8 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2XB_X3M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=2.75e-07 
M1 7 1 VSS VPW nch L=4e-08 W=4e-07 
M2 Y A 7 VPW nch L=4e-08 W=4e-07 
M3 8 A Y VPW nch L=4e-08 W=4e-07 
M4 VSS 1 8 VPW nch L=4e-08 W=4e-07 
M5 9 1 VSS VPW nch L=4e-08 W=4e-07 
M6 Y A 9 VPW nch L=4e-08 W=4e-07 
M7 VDD BN 1 VNW pch L=4e-08 W=3.5e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M9 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M10 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M11 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M12 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M13 VDD A Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2XB_X4M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 2 VPW nch L=4e-08 W=3.7e-07 
M1 8 2 VSS VPW nch L=4e-08 W=4e-07 
M2 Y A 8 VPW nch L=4e-08 W=4e-07 
M3 9 A Y VPW nch L=4e-08 W=4e-07 
M4 VSS 2 9 VPW nch L=4e-08 W=4e-07 
M5 10 2 VSS VPW nch L=4e-08 W=4e-07 
M6 Y A 10 VPW nch L=4e-08 W=4e-07 
M7 11 A Y VPW nch L=4e-08 W=4e-07 
M8 VSS 2 11 VPW nch L=4e-08 W=4e-07 
M9 2 BN VDD VNW pch L=4e-08 W=2.35e-07 
M10 VDD BN 2 VNW pch L=4e-08 W=2.35e-07 
M11 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M12 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M13 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M14 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M15 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M16 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M17 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M18 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2XB_X6M_A9TR Y VDD VNW VPW VSS A BN
M0 3 BN VSS VPW nch L=4e-08 W=2.75e-07 
M1 VSS BN 3 VPW nch L=4e-08 W=2.75e-07 
M2 7 3 VSS VPW nch L=4e-08 W=4e-07 
M3 Y A 7 VPW nch L=4e-08 W=4e-07 
M4 8 A Y VPW nch L=4e-08 W=4e-07 
M5 VSS 3 8 VPW nch L=4e-08 W=4e-07 
M6 9 3 VSS VPW nch L=4e-08 W=4e-07 
M7 Y A 9 VPW nch L=4e-08 W=4e-07 
M8 10 A Y VPW nch L=4e-08 W=4e-07 
M9 VSS 3 10 VPW nch L=4e-08 W=4e-07 
M10 11 3 VSS VPW nch L=4e-08 W=4e-07 
M11 Y A 11 VPW nch L=4e-08 W=4e-07 
M12 12 A Y VPW nch L=4e-08 W=4e-07 
M13 VSS 3 12 VPW nch L=4e-08 W=4e-07 
M14 3 BN VDD VNW pch L=4e-08 W=3.5e-07 
M15 VDD BN 3 VNW pch L=4e-08 W=3.5e-07 
M16 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M17 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M18 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M19 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M20 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M21 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M22 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M23 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M24 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M25 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M26 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M27 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2XB_X8M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=2.45e-07 
M1 1 BN VSS VPW nch L=4e-08 W=2.45e-07 
M2 VSS BN 1 VPW nch L=4e-08 W=2.45e-07 
M3 7 1 VSS VPW nch L=4e-08 W=4e-07 
M4 Y A 7 VPW nch L=4e-08 W=4e-07 
M5 8 A Y VPW nch L=4e-08 W=4e-07 
M6 VSS 1 8 VPW nch L=4e-08 W=4e-07 
M7 9 1 VSS VPW nch L=4e-08 W=4e-07 
M8 Y A 9 VPW nch L=4e-08 W=4e-07 
M9 10 A Y VPW nch L=4e-08 W=4e-07 
M10 VSS 1 10 VPW nch L=4e-08 W=4e-07 
M11 11 1 VSS VPW nch L=4e-08 W=4e-07 
M12 Y A 11 VPW nch L=4e-08 W=4e-07 
M13 12 A Y VPW nch L=4e-08 W=4e-07 
M14 VSS 1 12 VPW nch L=4e-08 W=4e-07 
M15 13 1 VSS VPW nch L=4e-08 W=4e-07 
M16 Y A 13 VPW nch L=4e-08 W=4e-07 
M17 14 A Y VPW nch L=4e-08 W=4e-07 
M18 VSS 1 14 VPW nch L=4e-08 W=4e-07 
M19 VDD BN 1 VNW pch L=4e-08 W=3.15e-07 
M20 1 BN VDD VNW pch L=4e-08 W=3.15e-07 
M21 VDD BN 1 VNW pch L=4e-08 W=3.15e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M23 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M24 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M25 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M26 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M27 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M28 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M29 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M30 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M31 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M32 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M33 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M34 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M35 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M36 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M37 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2_X0P5A_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=2e-07 
M1 Y A 6 VPW nch L=4e-08 W=2e-07 
M2 Y B VDD VNW pch L=4e-08 W=1.95e-07 
M3 VDD A Y VNW pch L=4e-08 W=1.95e-07 
.ENDS


.SUBCKT NAND2_X0P5B_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=1.7e-07 
M1 Y A 6 VPW nch L=4e-08 W=1.7e-07 
M2 Y B VDD VNW pch L=4e-08 W=2e-07 
M3 VDD A Y VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT NAND2_X0P5M_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=2e-07 
M1 Y A 6 VPW nch L=4e-08 W=2e-07 
M2 Y B VDD VNW pch L=4e-08 W=1.7e-07 
M3 VDD A Y VNW pch L=4e-08 W=1.7e-07 
.ENDS


.SUBCKT NAND2_X0P7A_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=2.8e-07 
M1 Y A 6 VPW nch L=4e-08 W=2.8e-07 
M2 Y B VDD VNW pch L=4e-08 W=2.75e-07 
M3 VDD A Y VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT NAND2_X0P7B_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=2.45e-07 
M1 Y A 6 VPW nch L=4e-08 W=2.45e-07 
M2 Y B VDD VNW pch L=4e-08 W=2.85e-07 
M3 VDD A Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NAND2_X0P7M_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=2.85e-07 
M1 Y A 6 VPW nch L=4e-08 W=2.85e-07 
M2 Y B VDD VNW pch L=4e-08 W=2.45e-07 
M3 VDD A Y VNW pch L=4e-08 W=2.45e-07 
.ENDS


.SUBCKT NAND2_X1A_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.9e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.9e-07 
M2 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M3 VDD A Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND2_X1B_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.45e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.45e-07 
M2 Y B VDD VNW pch L=4e-08 W=4e-07 
M3 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NAND2_X1M_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=4e-07 
M1 Y A 6 VPW nch L=4e-08 W=4e-07 
M2 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M3 VDD A Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2_X1P4A_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=2.8e-07 
M1 Y A 6 VPW nch L=4e-08 W=2.8e-07 
M2 7 A Y VPW nch L=4e-08 W=2.8e-07 
M3 VSS B 7 VPW nch L=4e-08 W=2.8e-07 
M4 Y B VDD VNW pch L=4e-08 W=2.75e-07 
M5 VDD A Y VNW pch L=4e-08 W=2.75e-07 
M6 Y A VDD VNW pch L=4e-08 W=2.75e-07 
M7 VDD B Y VNW pch L=4e-08 W=2.75e-07 
.ENDS


.SUBCKT NAND2_X1P4B_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=2.45e-07 
M1 Y A 6 VPW nch L=4e-08 W=2.45e-07 
M2 7 A Y VPW nch L=4e-08 W=2.45e-07 
M3 VSS B 7 VPW nch L=4e-08 W=2.45e-07 
M4 Y B VDD VNW pch L=4e-08 W=2.85e-07 
M5 VDD A Y VNW pch L=4e-08 W=2.85e-07 
M6 Y A VDD VNW pch L=4e-08 W=2.85e-07 
M7 VDD B Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NAND2_X1P4M_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=2.85e-07 
M1 Y A 6 VPW nch L=4e-08 W=2.85e-07 
M2 7 A Y VPW nch L=4e-08 W=2.85e-07 
M3 VSS B 7 VPW nch L=4e-08 W=2.85e-07 
M4 Y B VDD VNW pch L=4e-08 W=2.45e-07 
M5 VDD A Y VNW pch L=4e-08 W=2.45e-07 
M6 Y A VDD VNW pch L=4e-08 W=2.45e-07 
M7 VDD B Y VNW pch L=4e-08 W=2.45e-07 
.ENDS


.SUBCKT NAND2_X2A_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.9e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.9e-07 
M2 7 A Y VPW nch L=4e-08 W=3.9e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.9e-07 
M4 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M5 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M6 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M7 VDD B Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND2_X2B_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.45e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.45e-07 
M2 7 A Y VPW nch L=4e-08 W=3.45e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.45e-07 
M4 Y B VDD VNW pch L=4e-08 W=4e-07 
M5 VDD A Y VNW pch L=4e-08 W=4e-07 
M6 Y A VDD VNW pch L=4e-08 W=4e-07 
M7 VDD B Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NAND2_X2M_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=4e-07 
M1 Y A 6 VPW nch L=4e-08 W=4e-07 
M2 7 A Y VPW nch L=4e-08 W=4e-07 
M3 VSS B 7 VPW nch L=4e-08 W=4e-07 
M4 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M5 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M6 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M7 VDD B Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2_X3A_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.9e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.9e-07 
M2 7 A Y VPW nch L=4e-08 W=3.9e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.9e-07 
M4 8 B VSS VPW nch L=4e-08 W=3.9e-07 
M5 Y A 8 VPW nch L=4e-08 W=3.9e-07 
M6 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M7 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M8 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M9 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M10 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M11 VDD A Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND2_X3B_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.45e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.45e-07 
M2 7 A Y VPW nch L=4e-08 W=3.45e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.45e-07 
M4 8 B VSS VPW nch L=4e-08 W=3.45e-07 
M5 Y A 8 VPW nch L=4e-08 W=3.45e-07 
M6 Y B VDD VNW pch L=4e-08 W=4e-07 
M7 VDD A Y VNW pch L=4e-08 W=4e-07 
M8 Y A VDD VNW pch L=4e-08 W=4e-07 
M9 VDD B Y VNW pch L=4e-08 W=4e-07 
M10 Y B VDD VNW pch L=4e-08 W=4e-07 
M11 VDD A Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NAND2_X3M_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=4e-07 
M1 Y A 6 VPW nch L=4e-08 W=4e-07 
M2 7 A Y VPW nch L=4e-08 W=4e-07 
M3 VSS B 7 VPW nch L=4e-08 W=4e-07 
M4 8 B VSS VPW nch L=4e-08 W=4e-07 
M5 Y A 8 VPW nch L=4e-08 W=4e-07 
M6 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M7 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M8 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M9 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M10 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M11 VDD A Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2_X4A_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.9e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.9e-07 
M2 7 A Y VPW nch L=4e-08 W=3.9e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.9e-07 
M4 8 B VSS VPW nch L=4e-08 W=3.9e-07 
M5 Y A 8 VPW nch L=4e-08 W=3.9e-07 
M6 9 A Y VPW nch L=4e-08 W=3.9e-07 
M7 VSS B 9 VPW nch L=4e-08 W=3.9e-07 
M8 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M9 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M10 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M11 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M12 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M13 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M14 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M15 VDD B Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND2_X4B_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.45e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.45e-07 
M2 7 A Y VPW nch L=4e-08 W=3.45e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.45e-07 
M4 8 B VSS VPW nch L=4e-08 W=3.45e-07 
M5 Y A 8 VPW nch L=4e-08 W=3.45e-07 
M6 9 A Y VPW nch L=4e-08 W=3.45e-07 
M7 VSS B 9 VPW nch L=4e-08 W=3.45e-07 
M8 Y B VDD VNW pch L=4e-08 W=4e-07 
M9 VDD A Y VNW pch L=4e-08 W=4e-07 
M10 Y A VDD VNW pch L=4e-08 W=4e-07 
M11 VDD B Y VNW pch L=4e-08 W=4e-07 
M12 Y B VDD VNW pch L=4e-08 W=4e-07 
M13 VDD A Y VNW pch L=4e-08 W=4e-07 
M14 Y A VDD VNW pch L=4e-08 W=4e-07 
M15 VDD B Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NAND2_X4M_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=4e-07 
M1 Y A 6 VPW nch L=4e-08 W=4e-07 
M2 7 A Y VPW nch L=4e-08 W=4e-07 
M3 VSS B 7 VPW nch L=4e-08 W=4e-07 
M4 8 B VSS VPW nch L=4e-08 W=4e-07 
M5 Y A 8 VPW nch L=4e-08 W=4e-07 
M6 9 A Y VPW nch L=4e-08 W=4e-07 
M7 VSS B 9 VPW nch L=4e-08 W=4e-07 
M8 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M9 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M10 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M11 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M12 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M13 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M14 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M15 VDD B Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2_X6A_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.9e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.9e-07 
M2 7 A Y VPW nch L=4e-08 W=3.9e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.9e-07 
M4 8 B VSS VPW nch L=4e-08 W=3.9e-07 
M5 Y A 8 VPW nch L=4e-08 W=3.9e-07 
M6 9 A Y VPW nch L=4e-08 W=3.9e-07 
M7 VSS B 9 VPW nch L=4e-08 W=3.9e-07 
M8 10 B VSS VPW nch L=4e-08 W=3.9e-07 
M9 Y A 10 VPW nch L=4e-08 W=3.9e-07 
M10 11 A Y VPW nch L=4e-08 W=3.9e-07 
M11 VSS B 11 VPW nch L=4e-08 W=3.9e-07 
M12 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M13 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M14 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M15 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M16 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M17 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M18 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M19 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M20 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M21 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M22 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M23 VDD B Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND2_X6B_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.45e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.45e-07 
M2 7 A Y VPW nch L=4e-08 W=3.45e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.45e-07 
M4 8 B VSS VPW nch L=4e-08 W=3.45e-07 
M5 Y A 8 VPW nch L=4e-08 W=3.45e-07 
M6 9 A Y VPW nch L=4e-08 W=3.45e-07 
M7 VSS B 9 VPW nch L=4e-08 W=3.45e-07 
M8 10 B VSS VPW nch L=4e-08 W=3.45e-07 
M9 Y A 10 VPW nch L=4e-08 W=3.45e-07 
M10 11 A Y VPW nch L=4e-08 W=3.45e-07 
M11 VSS B 11 VPW nch L=4e-08 W=3.45e-07 
M12 Y B VDD VNW pch L=4e-08 W=4e-07 
M13 VDD A Y VNW pch L=4e-08 W=4e-07 
M14 Y A VDD VNW pch L=4e-08 W=4e-07 
M15 VDD B Y VNW pch L=4e-08 W=4e-07 
M16 Y B VDD VNW pch L=4e-08 W=4e-07 
M17 VDD A Y VNW pch L=4e-08 W=4e-07 
M18 Y A VDD VNW pch L=4e-08 W=4e-07 
M19 VDD B Y VNW pch L=4e-08 W=4e-07 
M20 Y B VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A Y VNW pch L=4e-08 W=4e-07 
M22 Y A VDD VNW pch L=4e-08 W=4e-07 
M23 VDD B Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NAND2_X6M_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=4e-07 
M1 Y A 6 VPW nch L=4e-08 W=4e-07 
M2 7 A Y VPW nch L=4e-08 W=4e-07 
M3 VSS B 7 VPW nch L=4e-08 W=4e-07 
M4 8 B VSS VPW nch L=4e-08 W=4e-07 
M5 Y A 8 VPW nch L=4e-08 W=4e-07 
M6 9 A Y VPW nch L=4e-08 W=4e-07 
M7 VSS B 9 VPW nch L=4e-08 W=4e-07 
M8 10 B VSS VPW nch L=4e-08 W=4e-07 
M9 Y A 10 VPW nch L=4e-08 W=4e-07 
M10 11 A Y VPW nch L=4e-08 W=4e-07 
M11 VSS B 11 VPW nch L=4e-08 W=4e-07 
M12 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M13 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M14 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M15 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M16 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M17 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M18 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M19 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M20 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M21 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M22 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M23 VDD B Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND2_X8A_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.9e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.9e-07 
M2 7 A Y VPW nch L=4e-08 W=3.9e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.9e-07 
M4 8 B VSS VPW nch L=4e-08 W=3.9e-07 
M5 Y A 8 VPW nch L=4e-08 W=3.9e-07 
M6 9 A Y VPW nch L=4e-08 W=3.9e-07 
M7 VSS B 9 VPW nch L=4e-08 W=3.9e-07 
M8 10 B VSS VPW nch L=4e-08 W=3.9e-07 
M9 Y A 10 VPW nch L=4e-08 W=3.9e-07 
M10 11 A Y VPW nch L=4e-08 W=3.9e-07 
M11 VSS B 11 VPW nch L=4e-08 W=3.9e-07 
M12 12 B VSS VPW nch L=4e-08 W=3.9e-07 
M13 Y A 12 VPW nch L=4e-08 W=3.9e-07 
M14 13 A Y VPW nch L=4e-08 W=3.9e-07 
M15 VSS B 13 VPW nch L=4e-08 W=3.9e-07 
M16 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M17 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M18 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M19 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M20 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M21 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M22 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M23 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M24 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M25 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M26 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M27 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M28 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M29 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M30 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M31 VDD B Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND2_X8B_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=3.45e-07 
M1 Y A 6 VPW nch L=4e-08 W=3.45e-07 
M2 7 A Y VPW nch L=4e-08 W=3.45e-07 
M3 VSS B 7 VPW nch L=4e-08 W=3.45e-07 
M4 8 B VSS VPW nch L=4e-08 W=3.45e-07 
M5 Y A 8 VPW nch L=4e-08 W=3.45e-07 
M6 9 A Y VPW nch L=4e-08 W=3.45e-07 
M7 VSS B 9 VPW nch L=4e-08 W=3.45e-07 
M8 10 B VSS VPW nch L=4e-08 W=3.45e-07 
M9 Y A 10 VPW nch L=4e-08 W=3.45e-07 
M10 11 A Y VPW nch L=4e-08 W=3.45e-07 
M11 VSS B 11 VPW nch L=4e-08 W=3.45e-07 
M12 12 B VSS VPW nch L=4e-08 W=3.45e-07 
M13 Y A 12 VPW nch L=4e-08 W=3.45e-07 
M14 13 A Y VPW nch L=4e-08 W=3.45e-07 
M15 VSS B 13 VPW nch L=4e-08 W=3.45e-07 
M16 Y B VDD VNW pch L=4e-08 W=4e-07 
M17 VDD A Y VNW pch L=4e-08 W=4e-07 
M18 Y A VDD VNW pch L=4e-08 W=4e-07 
M19 VDD B Y VNW pch L=4e-08 W=4e-07 
M20 Y B VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A Y VNW pch L=4e-08 W=4e-07 
M22 Y A VDD VNW pch L=4e-08 W=4e-07 
M23 VDD B Y VNW pch L=4e-08 W=4e-07 
M24 Y B VDD VNW pch L=4e-08 W=4e-07 
M25 VDD A Y VNW pch L=4e-08 W=4e-07 
M26 Y A VDD VNW pch L=4e-08 W=4e-07 
M27 VDD B Y VNW pch L=4e-08 W=4e-07 
M28 Y B VDD VNW pch L=4e-08 W=4e-07 
M29 VDD A Y VNW pch L=4e-08 W=4e-07 
M30 Y A VDD VNW pch L=4e-08 W=4e-07 
M31 VDD B Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NAND2_X8M_A9TR Y VDD VNW VPW VSS A B
M0 6 B VSS VPW nch L=4e-08 W=4e-07 
M1 Y A 6 VPW nch L=4e-08 W=4e-07 
M2 7 A Y VPW nch L=4e-08 W=4e-07 
M3 VSS B 7 VPW nch L=4e-08 W=4e-07 
M4 8 B VSS VPW nch L=4e-08 W=4e-07 
M5 Y A 8 VPW nch L=4e-08 W=4e-07 
M6 9 A Y VPW nch L=4e-08 W=4e-07 
M7 VSS B 9 VPW nch L=4e-08 W=4e-07 
M8 10 B VSS VPW nch L=4e-08 W=4e-07 
M9 Y A 10 VPW nch L=4e-08 W=4e-07 
M10 11 A Y VPW nch L=4e-08 W=4e-07 
M11 VSS B 11 VPW nch L=4e-08 W=4e-07 
M12 12 B VSS VPW nch L=4e-08 W=4e-07 
M13 Y A 12 VPW nch L=4e-08 W=4e-07 
M14 13 A Y VPW nch L=4e-08 W=4e-07 
M15 VSS B 13 VPW nch L=4e-08 W=4e-07 
M16 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M17 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M18 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M19 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M20 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M21 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M22 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M23 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M24 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M25 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M26 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M27 VDD B Y VNW pch L=4e-08 W=3.45e-07 
M28 Y B VDD VNW pch L=4e-08 W=3.45e-07 
M29 VDD A Y VNW pch L=4e-08 W=3.45e-07 
M30 Y A VDD VNW pch L=4e-08 W=3.45e-07 
M31 VDD B Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND3BB_X0P5M_A9TR Y VDD VNW VPW VSS AN BN C
M0 2 AN VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=1.2e-07 
M2 9 C VSS VPW nch L=4e-08 W=2e-07 
M3 Y 2 9 VPW nch L=4e-08 W=2e-07 
M4 8 AN 2 VNW pch L=4e-08 W=2.1e-07 
M5 VDD BN 8 VNW pch L=4e-08 W=2.1e-07 
M6 Y C VDD VNW pch L=4e-08 W=1.7e-07 
M7 VDD 2 Y VNW pch L=4e-08 W=1.7e-07 
.ENDS


.SUBCKT NAND3BB_X0P7M_A9TR Y VDD VNW VPW VSS AN BN C
M0 2 AN VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=1.2e-07 
M2 9 C VSS VPW nch L=4e-08 W=2.85e-07 
M3 Y 2 9 VPW nch L=4e-08 W=2.85e-07 
M4 8 AN 2 VNW pch L=4e-08 W=2.6e-07 
M5 VDD BN 8 VNW pch L=4e-08 W=2.6e-07 
M6 Y C VDD VNW pch L=4e-08 W=2.45e-07 
M7 VDD 2 Y VNW pch L=4e-08 W=2.45e-07 
.ENDS


.SUBCKT NAND3BB_X1M_A9TR Y VDD VNW VPW VSS AN BN C
M0 2 AN VSS VPW nch L=4e-08 W=1.3e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=1.3e-07 
M2 9 C VSS VPW nch L=4e-08 W=3.9e-07 
M3 Y 2 9 VPW nch L=4e-08 W=3.9e-07 
M4 8 AN 2 VNW pch L=4e-08 W=3.25e-07 
M5 VDD BN 8 VNW pch L=4e-08 W=3.25e-07 
M6 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M7 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND3BB_X1P4M_A9TR Y VDD VNW VPW VSS AN BN C
M0 2 AN VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=1.6e-07 
M2 9 C VSS VPW nch L=4e-08 W=2.85e-07 
M3 Y 2 9 VPW nch L=4e-08 W=2.85e-07 
M4 10 2 Y VPW nch L=4e-08 W=2.85e-07 
M5 VSS C 10 VPW nch L=4e-08 W=2.85e-07 
M6 8 AN 2 VNW pch L=4e-08 W=4e-07 
M7 VDD BN 8 VNW pch L=4e-08 W=4e-07 
M8 Y C VDD VNW pch L=4e-08 W=2.45e-07 
M9 VDD 2 Y VNW pch L=4e-08 W=2.45e-07 
M10 Y 2 VDD VNW pch L=4e-08 W=2.45e-07 
M11 VDD C Y VNW pch L=4e-08 W=2.45e-07 
.ENDS


.SUBCKT NAND3BB_X2M_A9TR Y VDD VNW VPW VSS AN BN C
M0 3 BN VSS VPW nch L=4e-08 W=2.55e-07 
M1 VSS AN 3 VPW nch L=4e-08 W=2.55e-07 
M2 11 C VSS VPW nch L=4e-08 W=4e-07 
M3 Y 3 11 VPW nch L=4e-08 W=4e-07 
M4 12 3 Y VPW nch L=4e-08 W=4e-07 
M5 VSS C 12 VPW nch L=4e-08 W=4e-07 
M6 8 BN VDD VNW pch L=4e-08 W=3.15e-07 
M7 3 AN 8 VNW pch L=4e-08 W=3.15e-07 
M8 9 AN 3 VNW pch L=4e-08 W=3.15e-07 
M9 VDD BN 9 VNW pch L=4e-08 W=3.15e-07 
M10 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M11 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M12 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M13 VDD C Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND3BB_X3M_A9TR Y VDD VNW VPW VSS AN BN C
M0 3 BN VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS AN 3 VPW nch L=4e-08 W=3.2e-07 
M2 11 C VSS VPW nch L=4e-08 W=4e-07 
M3 Y 3 11 VPW nch L=4e-08 W=4e-07 
M4 12 3 Y VPW nch L=4e-08 W=4e-07 
M5 VSS C 12 VPW nch L=4e-08 W=4e-07 
M6 13 C VSS VPW nch L=4e-08 W=4e-07 
M7 Y 3 13 VPW nch L=4e-08 W=4e-07 
M8 8 BN VDD VNW pch L=4e-08 W=4e-07 
M9 3 AN 8 VNW pch L=4e-08 W=4e-07 
M10 9 AN 3 VNW pch L=4e-08 W=4e-07 
M11 VDD BN 9 VNW pch L=4e-08 W=4e-07 
M12 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M13 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M15 VDD C Y VNW pch L=4e-08 W=3.45e-07 
M16 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M17 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND3BB_X4M_A9TR Y VDD VNW VPW VSS AN BN C
M0 2 AN VSS VPW nch L=4e-08 W=2.4e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=2.4e-07 
M2 2 BN VSS VPW nch L=4e-08 W=2.4e-07 
M3 VSS AN 2 VPW nch L=4e-08 W=2.4e-07 
M4 12 C VSS VPW nch L=4e-08 W=4e-07 
M5 Y 2 12 VPW nch L=4e-08 W=4e-07 
M6 13 2 Y VPW nch L=4e-08 W=4e-07 
M7 VSS C 13 VPW nch L=4e-08 W=4e-07 
M8 14 C VSS VPW nch L=4e-08 W=4e-07 
M9 Y 2 14 VPW nch L=4e-08 W=4e-07 
M10 15 2 Y VPW nch L=4e-08 W=4e-07 
M11 VSS C 15 VPW nch L=4e-08 W=4e-07 
M12 8 AN 2 VNW pch L=4e-08 W=4e-07 
M13 VDD BN 8 VNW pch L=4e-08 W=4e-07 
M14 9 BN VDD VNW pch L=4e-08 W=4e-07 
M15 2 AN 9 VNW pch L=4e-08 W=4e-07 
M16 10 AN 2 VNW pch L=4e-08 W=4e-07 
M17 VDD BN 10 VNW pch L=4e-08 W=4e-07 
M18 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M19 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M20 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M21 VDD C Y VNW pch L=4e-08 W=3.45e-07 
M22 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M23 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M24 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M25 VDD C Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND3BB_X6M_A9TR Y VDD VNW VPW VSS AN BN C
M0 2 BN VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS AN 2 VPW nch L=4e-08 W=3.2e-07 
M2 2 AN VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS BN 2 VPW nch L=4e-08 W=3.2e-07 
M4 14 C VSS VPW nch L=4e-08 W=4e-07 
M5 Y 2 14 VPW nch L=4e-08 W=4e-07 
M6 15 2 Y VPW nch L=4e-08 W=4e-07 
M7 VSS C 15 VPW nch L=4e-08 W=4e-07 
M8 16 C VSS VPW nch L=4e-08 W=4e-07 
M9 Y 2 16 VPW nch L=4e-08 W=4e-07 
M10 17 2 Y VPW nch L=4e-08 W=4e-07 
M11 VSS C 17 VPW nch L=4e-08 W=4e-07 
M12 18 C VSS VPW nch L=4e-08 W=4e-07 
M13 Y 2 18 VPW nch L=4e-08 W=4e-07 
M14 19 2 Y VPW nch L=4e-08 W=4e-07 
M15 VSS C 19 VPW nch L=4e-08 W=4e-07 
M16 8 BN VDD VNW pch L=4e-08 W=4e-07 
M17 2 AN 8 VNW pch L=4e-08 W=4e-07 
M18 9 AN 2 VNW pch L=4e-08 W=4e-07 
M19 VDD BN 9 VNW pch L=4e-08 W=4e-07 
M20 10 BN VDD VNW pch L=4e-08 W=4e-07 
M21 2 AN 10 VNW pch L=4e-08 W=4e-07 
M22 11 AN 2 VNW pch L=4e-08 W=4e-07 
M23 VDD BN 11 VNW pch L=4e-08 W=4e-07 
M24 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M25 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M26 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M27 VDD C Y VNW pch L=4e-08 W=3.45e-07 
M28 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M29 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M30 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M31 VDD C Y VNW pch L=4e-08 W=3.45e-07 
M32 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M33 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M34 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M35 VDD C Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND3BB_X8M_A9TR Y VDD VNW VPW VSS AN BN C
M0 2 AN VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=3.2e-07 
M2 2 BN VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS AN 2 VPW nch L=4e-08 W=3.2e-07 
M4 2 AN VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS BN 2 VPW nch L=4e-08 W=3.2e-07 
M6 16 C VSS VPW nch L=4e-08 W=4e-07 
M7 Y 2 16 VPW nch L=4e-08 W=4e-07 
M8 17 2 Y VPW nch L=4e-08 W=4e-07 
M9 VSS C 17 VPW nch L=4e-08 W=4e-07 
M10 18 C VSS VPW nch L=4e-08 W=4e-07 
M11 Y 2 18 VPW nch L=4e-08 W=4e-07 
M12 19 2 Y VPW nch L=4e-08 W=4e-07 
M13 VSS C 19 VPW nch L=4e-08 W=4e-07 
M14 20 C VSS VPW nch L=4e-08 W=4e-07 
M15 Y 2 20 VPW nch L=4e-08 W=4e-07 
M16 21 2 Y VPW nch L=4e-08 W=4e-07 
M17 VSS C 21 VPW nch L=4e-08 W=4e-07 
M18 22 C VSS VPW nch L=4e-08 W=4e-07 
M19 Y 2 22 VPW nch L=4e-08 W=4e-07 
M20 23 2 Y VPW nch L=4e-08 W=4e-07 
M21 VSS C 23 VPW nch L=4e-08 W=4e-07 
M22 8 BN VDD VNW pch L=4e-08 W=4e-07 
M23 2 AN 8 VNW pch L=4e-08 W=4e-07 
M24 9 AN 2 VNW pch L=4e-08 W=4e-07 
M25 VDD BN 9 VNW pch L=4e-08 W=4e-07 
M26 10 BN VDD VNW pch L=4e-08 W=4e-07 
M27 2 AN 10 VNW pch L=4e-08 W=4e-07 
M28 11 AN 2 VNW pch L=4e-08 W=4e-07 
M29 VDD BN 11 VNW pch L=4e-08 W=4e-07 
M30 12 BN VDD VNW pch L=4e-08 W=4e-07 
M31 2 AN 12 VNW pch L=4e-08 W=4e-07 
M32 13 AN 2 VNW pch L=4e-08 W=4e-07 
M33 VDD BN 13 VNW pch L=4e-08 W=4e-07 
M34 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M35 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M36 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M37 VDD C Y VNW pch L=4e-08 W=3.45e-07 
M38 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M39 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M40 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M41 VDD C Y VNW pch L=4e-08 W=3.45e-07 
M42 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M43 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M44 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M45 VDD C Y VNW pch L=4e-08 W=3.45e-07 
M46 Y C VDD VNW pch L=4e-08 W=3.45e-07 
M47 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M48 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M49 VDD C Y VNW pch L=4e-08 W=3.45e-07 
.ENDS


.SUBCKT NAND3B_X0P5M_A9TR Y VDD VNW VPW VSS AN B C
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 C VSS VPW nch L=4e-08 W=2e-07 
M2 9 B 8 VPW nch L=4e-08 W=2e-07 
M3 Y 1 9 VPW nch L=4e-08 W=2e-07 
M4 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M5 Y C VDD VNW pch L=4e-08 W=1.35e-07 
M6 VDD B Y VNW pch L=4e-08 W=1.35e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=1.35e-07 
.ENDS


.SUBCKT NAND3B_X0P7M_A9TR Y VDD VNW VPW VSS AN B C
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 C VSS VPW nch L=4e-08 W=2.85e-07 
M2 9 B 8 VPW nch L=4e-08 W=2.85e-07 
M3 Y 1 9 VPW nch L=4e-08 W=2.85e-07 
M4 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M5 Y C VDD VNW pch L=4e-08 W=1.9e-07 
M6 VDD B Y VNW pch L=4e-08 W=1.9e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT NAND3B_X1M_A9TR Y VDD VNW VPW VSS AN B C
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 C VSS VPW nch L=4e-08 W=3.9e-07 
M2 9 B 8 VPW nch L=4e-08 W=3.9e-07 
M3 Y 1 9 VPW nch L=4e-08 W=3.9e-07 
M4 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M5 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M6 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3B_X1P4M_A9TR Y VDD VNW VPW VSS AN B C
M0 VSS AN 1 VPW nch L=4e-08 W=1.3e-07 
M1 VSS C 4 VPW nch L=4e-08 W=2.85e-07 
M2 4 C VSS VPW nch L=4e-08 W=2.85e-07 
M3 9 B 4 VPW nch L=4e-08 W=2.85e-07 
M4 Y 1 9 VPW nch L=4e-08 W=2.85e-07 
M5 10 1 Y VPW nch L=4e-08 W=2.85e-07 
M6 4 B 10 VPW nch L=4e-08 W=2.85e-07 
M7 VDD AN 1 VNW pch L=4e-08 W=1.65e-07 
M8 Y C VDD VNW pch L=4e-08 W=1.9e-07 
M9 VDD C Y VNW pch L=4e-08 W=1.9e-07 
M10 Y B VDD VNW pch L=4e-08 W=1.9e-07 
M11 VDD 1 Y VNW pch L=4e-08 W=1.9e-07 
M12 Y 1 VDD VNW pch L=4e-08 W=1.9e-07 
M13 VDD B Y VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT NAND3B_X2M_A9TR Y VDD VNW VPW VSS AN B C
M0 VSS AN 1 VPW nch L=4e-08 W=1.7e-07 
M1 VSS C 4 VPW nch L=4e-08 W=4e-07 
M2 4 C VSS VPW nch L=4e-08 W=4e-07 
M3 9 B 4 VPW nch L=4e-08 W=4e-07 
M4 Y 1 9 VPW nch L=4e-08 W=4e-07 
M5 10 1 Y VPW nch L=4e-08 W=4e-07 
M6 4 B 10 VPW nch L=4e-08 W=4e-07 
M7 VDD AN 1 VNW pch L=4e-08 W=2.2e-07 
M8 Y C VDD VNW pch L=4e-08 W=2.6e-07 
M9 VDD C Y VNW pch L=4e-08 W=2.6e-07 
M10 Y B VDD VNW pch L=4e-08 W=2.6e-07 
M11 VDD 1 Y VNW pch L=4e-08 W=2.6e-07 
M12 Y 1 VDD VNW pch L=4e-08 W=2.6e-07 
M13 VDD B Y VNW pch L=4e-08 W=2.6e-07 
.ENDS


.SUBCKT NAND3B_X3M_A9TR Y VDD VNW VPW VSS AN B C
M0 VSS AN 1 VPW nch L=4e-08 W=2.5e-07 
M1 4 C VSS VPW nch L=4e-08 W=4e-07 
M2 VSS C 4 VPW nch L=4e-08 W=4e-07 
M3 4 C VSS VPW nch L=4e-08 W=4e-07 
M4 9 B 4 VPW nch L=4e-08 W=4e-07 
M5 Y 1 9 VPW nch L=4e-08 W=4e-07 
M6 10 1 Y VPW nch L=4e-08 W=4e-07 
M7 4 B 10 VPW nch L=4e-08 W=4e-07 
M8 11 B 4 VPW nch L=4e-08 W=4e-07 
M9 Y 1 11 VPW nch L=4e-08 W=4e-07 
M10 VDD AN 1 VNW pch L=4e-08 W=3.2e-07 
M11 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M12 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M13 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M14 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M15 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
M16 VDD 1 Y VNW pch L=4e-08 W=2.65e-07 
M17 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M18 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M19 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3B_X4M_A9TR Y VDD VNW VPW VSS AN B C
M0 VSS AN 1 VPW nch L=4e-08 W=3.1e-07 
M1 VSS C 4 VPW nch L=4e-08 W=4e-07 
M2 4 C VSS VPW nch L=4e-08 W=4e-07 
M3 VSS C 4 VPW nch L=4e-08 W=4e-07 
M4 4 C VSS VPW nch L=4e-08 W=4e-07 
M5 9 B 4 VPW nch L=4e-08 W=4e-07 
M6 Y 1 9 VPW nch L=4e-08 W=4e-07 
M7 10 1 Y VPW nch L=4e-08 W=4e-07 
M8 4 B 10 VPW nch L=4e-08 W=4e-07 
M9 11 B 4 VPW nch L=4e-08 W=4e-07 
M10 Y 1 11 VPW nch L=4e-08 W=4e-07 
M11 12 1 Y VPW nch L=4e-08 W=4e-07 
M12 4 B 12 VPW nch L=4e-08 W=4e-07 
M13 VDD AN 1 VNW pch L=4e-08 W=4e-07 
M14 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M15 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M16 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M17 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M18 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M19 VDD 1 Y VNW pch L=4e-08 W=2.65e-07 
M20 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
M21 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M22 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M23 VDD 1 Y VNW pch L=4e-08 W=2.65e-07 
M24 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
M25 VDD B Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3B_X6M_A9TR Y VDD VNW VPW VSS AN B C
M0 3 AN VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS AN 3 VPW nch L=4e-08 W=2.45e-07 
M2 VSS C 4 VPW nch L=4e-08 W=4e-07 
M3 4 C VSS VPW nch L=4e-08 W=4e-07 
M4 VSS C 4 VPW nch L=4e-08 W=4e-07 
M5 4 C VSS VPW nch L=4e-08 W=4e-07 
M6 VSS C 4 VPW nch L=4e-08 W=4e-07 
M7 4 C VSS VPW nch L=4e-08 W=4e-07 
M8 9 B 4 VPW nch L=4e-08 W=4e-07 
M9 Y 3 9 VPW nch L=4e-08 W=4e-07 
M10 10 3 Y VPW nch L=4e-08 W=4e-07 
M11 4 B 10 VPW nch L=4e-08 W=4e-07 
M12 11 B 4 VPW nch L=4e-08 W=4e-07 
M13 Y 3 11 VPW nch L=4e-08 W=4e-07 
M14 12 3 Y VPW nch L=4e-08 W=4e-07 
M15 4 B 12 VPW nch L=4e-08 W=4e-07 
M16 13 B 4 VPW nch L=4e-08 W=4e-07 
M17 Y 3 13 VPW nch L=4e-08 W=4e-07 
M18 14 3 Y VPW nch L=4e-08 W=4e-07 
M19 4 B 14 VPW nch L=4e-08 W=4e-07 
M20 3 AN VDD VNW pch L=4e-08 W=3.15e-07 
M21 VDD AN 3 VNW pch L=4e-08 W=3.15e-07 
M22 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M23 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M24 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M25 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M26 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M27 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M28 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M29 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M30 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M31 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M32 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M33 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M34 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M35 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M36 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M37 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M38 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M39 VDD B Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3XXB_X0P5M_A9TR Y VDD VNW VPW VSS A B CN
M0 VSS CN 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 1 VSS VPW nch L=4e-08 W=2e-07 
M2 9 B 8 VPW nch L=4e-08 W=2e-07 
M3 Y A 9 VPW nch L=4e-08 W=2e-07 
M4 VDD CN 1 VNW pch L=4e-08 W=1.55e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=1.35e-07 
M6 VDD B Y VNW pch L=4e-08 W=1.35e-07 
M7 Y A VDD VNW pch L=4e-08 W=1.35e-07 
.ENDS


.SUBCKT NAND3XXB_X0P7M_A9TR Y VDD VNW VPW VSS A B CN
M0 VSS CN 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 1 VSS VPW nch L=4e-08 W=2.85e-07 
M2 9 B 8 VPW nch L=4e-08 W=2.85e-07 
M3 Y A 9 VPW nch L=4e-08 W=2.85e-07 
M4 VDD CN 1 VNW pch L=4e-08 W=1.55e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=1.9e-07 
M6 VDD B Y VNW pch L=4e-08 W=1.9e-07 
M7 Y A VDD VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT NAND3XXB_X1M_A9TR Y VDD VNW VPW VSS A B CN
M0 VSS CN 1 VPW nch L=4e-08 W=1.2e-07 
M1 8 1 VSS VPW nch L=4e-08 W=4e-07 
M2 9 B 8 VPW nch L=4e-08 W=4e-07 
M3 Y A 9 VPW nch L=4e-08 W=4e-07 
M4 VDD CN 1 VNW pch L=4e-08 W=1.55e-07 
M5 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
M6 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M7 Y A VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3XXB_X1P4M_A9TR Y VDD VNW VPW VSS A B CN
M0 VSS CN 1 VPW nch L=4e-08 W=1.3e-07 
M1 VSS 1 4 VPW nch L=4e-08 W=2.85e-07 
M2 4 1 VSS VPW nch L=4e-08 W=2.85e-07 
M3 9 B 4 VPW nch L=4e-08 W=2.85e-07 
M4 Y A 9 VPW nch L=4e-08 W=2.85e-07 
M5 10 A Y VPW nch L=4e-08 W=2.85e-07 
M6 4 B 10 VPW nch L=4e-08 W=2.85e-07 
M7 VDD CN 1 VNW pch L=4e-08 W=1.65e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=1.9e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=1.9e-07 
M10 Y B VDD VNW pch L=4e-08 W=1.9e-07 
M11 VDD A Y VNW pch L=4e-08 W=1.9e-07 
M12 Y A VDD VNW pch L=4e-08 W=1.9e-07 
M13 VDD B Y VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT NAND3XXB_X2M_A9TR Y VDD VNW VPW VSS A B CN
M0 VSS CN 1 VPW nch L=4e-08 W=1.7e-07 
M1 VSS 1 4 VPW nch L=4e-08 W=4e-07 
M2 4 1 VSS VPW nch L=4e-08 W=4e-07 
M3 9 B 4 VPW nch L=4e-08 W=4e-07 
M4 Y A 9 VPW nch L=4e-08 W=4e-07 
M5 10 A Y VPW nch L=4e-08 W=4e-07 
M6 4 B 10 VPW nch L=4e-08 W=4e-07 
M7 VDD CN 1 VNW pch L=4e-08 W=2.2e-07 
M8 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=2.65e-07 
M10 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M11 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M12 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M13 VDD B Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3XXB_X3M_A9TR Y VDD VNW VPW VSS A B CN
M0 VSS CN 1 VPW nch L=4e-08 W=2.5e-07 
M1 4 1 VSS VPW nch L=4e-08 W=4e-07 
M2 VSS 1 4 VPW nch L=4e-08 W=4e-07 
M3 4 1 VSS VPW nch L=4e-08 W=4e-07 
M4 9 B 4 VPW nch L=4e-08 W=4e-07 
M5 Y A 9 VPW nch L=4e-08 W=4e-07 
M6 10 A Y VPW nch L=4e-08 W=4e-07 
M7 4 B 10 VPW nch L=4e-08 W=4e-07 
M8 11 B 4 VPW nch L=4e-08 W=4e-07 
M9 Y A 11 VPW nch L=4e-08 W=4e-07 
M10 VDD CN 1 VNW pch L=4e-08 W=3.2e-07 
M11 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
M12 VDD 1 Y VNW pch L=4e-08 W=2.65e-07 
M13 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
M14 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M15 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M16 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M17 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M18 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M19 Y A VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3XXB_X4M_A9TR Y VDD VNW VPW VSS A B CN
M0 VSS CN 1 VPW nch L=4e-08 W=3.1e-07 
M1 VSS 1 4 VPW nch L=4e-08 W=4e-07 
M2 4 1 VSS VPW nch L=4e-08 W=4e-07 
M3 VSS 1 4 VPW nch L=4e-08 W=4e-07 
M4 4 1 VSS VPW nch L=4e-08 W=4e-07 
M5 9 B 4 VPW nch L=4e-08 W=4e-07 
M6 Y A 9 VPW nch L=4e-08 W=4e-07 
M7 10 A Y VPW nch L=4e-08 W=4e-07 
M8 4 B 10 VPW nch L=4e-08 W=4e-07 
M9 11 B 4 VPW nch L=4e-08 W=4e-07 
M10 Y A 11 VPW nch L=4e-08 W=4e-07 
M11 12 A Y VPW nch L=4e-08 W=4e-07 
M12 4 B 12 VPW nch L=4e-08 W=4e-07 
M13 VDD CN 1 VNW pch L=4e-08 W=4e-07 
M14 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
M15 VDD 1 Y VNW pch L=4e-08 W=2.65e-07 
M16 Y 1 VDD VNW pch L=4e-08 W=2.65e-07 
M17 VDD 1 Y VNW pch L=4e-08 W=2.65e-07 
M18 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M19 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M20 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M21 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M22 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M23 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M24 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M25 VDD B Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3XXB_X6M_A9TR Y VDD VNW VPW VSS A B CN
M0 3 CN VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS CN 3 VPW nch L=4e-08 W=2.45e-07 
M2 VSS 3 4 VPW nch L=4e-08 W=4e-07 
M3 4 3 VSS VPW nch L=4e-08 W=4e-07 
M4 VSS 3 4 VPW nch L=4e-08 W=4e-07 
M5 4 3 VSS VPW nch L=4e-08 W=4e-07 
M6 VSS 3 4 VPW nch L=4e-08 W=4e-07 
M7 4 3 VSS VPW nch L=4e-08 W=4e-07 
M8 9 B 4 VPW nch L=4e-08 W=4e-07 
M9 Y A 9 VPW nch L=4e-08 W=4e-07 
M10 10 A Y VPW nch L=4e-08 W=4e-07 
M11 4 B 10 VPW nch L=4e-08 W=4e-07 
M12 11 B 4 VPW nch L=4e-08 W=4e-07 
M13 Y A 11 VPW nch L=4e-08 W=4e-07 
M14 12 A Y VPW nch L=4e-08 W=4e-07 
M15 4 B 12 VPW nch L=4e-08 W=4e-07 
M16 13 B 4 VPW nch L=4e-08 W=4e-07 
M17 Y A 13 VPW nch L=4e-08 W=4e-07 
M18 14 A Y VPW nch L=4e-08 W=4e-07 
M19 4 B 14 VPW nch L=4e-08 W=4e-07 
M20 3 CN VDD VNW pch L=4e-08 W=3.15e-07 
M21 VDD CN 3 VNW pch L=4e-08 W=3.15e-07 
M22 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M23 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M24 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M25 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M26 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M27 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M28 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M29 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M30 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M31 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M32 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M33 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M34 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M35 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M36 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M37 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M38 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M39 VDD B Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3_X0P5A_A9TR Y VDD VNW VPW VSS A B C
M0 7 C VSS VPW nch L=4e-08 W=2e-07 
M1 8 B 7 VPW nch L=4e-08 W=2e-07 
M2 Y A 8 VPW nch L=4e-08 W=2e-07 
M3 Y C VDD VNW pch L=4e-08 W=2e-07 
M4 VDD B Y VNW pch L=4e-08 W=2e-07 
M5 Y A VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT NAND3_X0P5M_A9TR Y VDD VNW VPW VSS A B C
M0 7 C VSS VPW nch L=4e-08 W=2e-07 
M1 8 B 7 VPW nch L=4e-08 W=2e-07 
M2 Y A 8 VPW nch L=4e-08 W=2e-07 
M3 Y C VDD VNW pch L=4e-08 W=1.35e-07 
M4 VDD B Y VNW pch L=4e-08 W=1.35e-07 
M5 Y A VDD VNW pch L=4e-08 W=1.35e-07 
.ENDS


.SUBCKT NAND3_X0P7A_A9TR Y VDD VNW VPW VSS A B C
M0 7 C VSS VPW nch L=4e-08 W=2.85e-07 
M1 8 B 7 VPW nch L=4e-08 W=2.85e-07 
M2 Y A 8 VPW nch L=4e-08 W=2.85e-07 
M3 Y C VDD VNW pch L=4e-08 W=2.85e-07 
M4 VDD B Y VNW pch L=4e-08 W=2.85e-07 
M5 Y A VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NAND3_X0P7M_A9TR Y VDD VNW VPW VSS A B C
M0 7 C VSS VPW nch L=4e-08 W=2.85e-07 
M1 8 B 7 VPW nch L=4e-08 W=2.85e-07 
M2 Y A 8 VPW nch L=4e-08 W=2.85e-07 
M3 Y C VDD VNW pch L=4e-08 W=1.9e-07 
M4 VDD B Y VNW pch L=4e-08 W=1.9e-07 
M5 Y A VDD VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT NAND3_X1A_A9TR Y VDD VNW VPW VSS A B C
M0 7 C VSS VPW nch L=4e-08 W=3.9e-07 
M1 8 B 7 VPW nch L=4e-08 W=3.9e-07 
M2 Y A 8 VPW nch L=4e-08 W=3.9e-07 
M3 Y C VDD VNW pch L=4e-08 W=3.65e-07 
M4 VDD B Y VNW pch L=4e-08 W=3.65e-07 
M5 Y A VDD VNW pch L=4e-08 W=3.65e-07 
.ENDS


.SUBCKT NAND3_X1M_A9TR Y VDD VNW VPW VSS A B C
M0 7 C VSS VPW nch L=4e-08 W=4e-07 
M1 8 B 7 VPW nch L=4e-08 W=4e-07 
M2 Y A 8 VPW nch L=4e-08 W=4e-07 
M3 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M4 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M5 Y A VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3_X1P4A_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=2.85e-07 
M1 1 C VSS VPW nch L=4e-08 W=2.85e-07 
M2 8 B 1 VPW nch L=4e-08 W=2.85e-07 
M3 Y A 8 VPW nch L=4e-08 W=2.85e-07 
M4 9 A Y VPW nch L=4e-08 W=2.85e-07 
M5 1 B 9 VPW nch L=4e-08 W=2.85e-07 
M6 Y C VDD VNW pch L=4e-08 W=2.85e-07 
M7 VDD C Y VNW pch L=4e-08 W=2.85e-07 
M8 Y B VDD VNW pch L=4e-08 W=2.85e-07 
M9 VDD A Y VNW pch L=4e-08 W=2.85e-07 
M10 Y A VDD VNW pch L=4e-08 W=2.85e-07 
M11 VDD B Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NAND3_X1P4M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=2.85e-07 
M1 1 C VSS VPW nch L=4e-08 W=2.85e-07 
M2 8 B 1 VPW nch L=4e-08 W=2.85e-07 
M3 Y A 8 VPW nch L=4e-08 W=2.85e-07 
M4 9 A Y VPW nch L=4e-08 W=2.85e-07 
M5 1 B 9 VPW nch L=4e-08 W=2.85e-07 
M6 Y C VDD VNW pch L=4e-08 W=1.9e-07 
M7 VDD C Y VNW pch L=4e-08 W=1.9e-07 
M8 Y B VDD VNW pch L=4e-08 W=1.9e-07 
M9 VDD A Y VNW pch L=4e-08 W=1.9e-07 
M10 Y A VDD VNW pch L=4e-08 W=1.9e-07 
M11 VDD B Y VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT NAND3_X2A_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=3.9e-07 
M1 1 C VSS VPW nch L=4e-08 W=3.9e-07 
M2 8 B 1 VPW nch L=4e-08 W=3.9e-07 
M3 Y A 8 VPW nch L=4e-08 W=3.9e-07 
M4 9 A Y VPW nch L=4e-08 W=3.9e-07 
M5 1 B 9 VPW nch L=4e-08 W=3.9e-07 
M6 Y C VDD VNW pch L=4e-08 W=3.9e-07 
M7 VDD C Y VNW pch L=4e-08 W=3.9e-07 
M8 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M9 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M10 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M11 VDD B Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND3_X2M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=4e-07 
M1 1 C VSS VPW nch L=4e-08 W=4e-07 
M2 8 B 1 VPW nch L=4e-08 W=4e-07 
M3 Y A 8 VPW nch L=4e-08 W=4e-07 
M4 9 A Y VPW nch L=4e-08 W=4e-07 
M5 1 B 9 VPW nch L=4e-08 W=4e-07 
M6 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M7 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M8 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M9 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M10 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M11 VDD B Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3_X3A_A9TR Y VDD VNW VPW VSS A B C
M0 3 C VSS VPW nch L=4e-08 W=3.9e-07 
M1 VSS C 3 VPW nch L=4e-08 W=3.9e-07 
M2 3 C VSS VPW nch L=4e-08 W=3.9e-07 
M3 8 B 3 VPW nch L=4e-08 W=3.9e-07 
M4 Y A 8 VPW nch L=4e-08 W=3.9e-07 
M5 9 A Y VPW nch L=4e-08 W=3.9e-07 
M6 3 B 9 VPW nch L=4e-08 W=3.9e-07 
M7 10 B 3 VPW nch L=4e-08 W=3.9e-07 
M8 Y A 10 VPW nch L=4e-08 W=3.9e-07 
M9 Y C VDD VNW pch L=4e-08 W=3.9e-07 
M10 VDD C Y VNW pch L=4e-08 W=3.9e-07 
M11 Y C VDD VNW pch L=4e-08 W=3.9e-07 
M12 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M13 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M14 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M15 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M16 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M17 Y A VDD VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND3_X3M_A9TR Y VDD VNW VPW VSS A B C
M0 3 C VSS VPW nch L=4e-08 W=4e-07 
M1 VSS C 3 VPW nch L=4e-08 W=4e-07 
M2 3 C VSS VPW nch L=4e-08 W=4e-07 
M3 8 B 3 VPW nch L=4e-08 W=4e-07 
M4 Y A 8 VPW nch L=4e-08 W=4e-07 
M5 9 A Y VPW nch L=4e-08 W=4e-07 
M6 3 B 9 VPW nch L=4e-08 W=4e-07 
M7 10 B 3 VPW nch L=4e-08 W=4e-07 
M8 Y A 10 VPW nch L=4e-08 W=4e-07 
M9 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M10 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M11 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M12 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M13 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M14 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M15 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M16 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M17 Y A VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3_X4A_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=3.9e-07 
M1 1 C VSS VPW nch L=4e-08 W=3.9e-07 
M2 VSS C 1 VPW nch L=4e-08 W=3.9e-07 
M3 1 C VSS VPW nch L=4e-08 W=3.9e-07 
M4 8 B 1 VPW nch L=4e-08 W=3.9e-07 
M5 Y A 8 VPW nch L=4e-08 W=3.9e-07 
M6 9 A Y VPW nch L=4e-08 W=3.9e-07 
M7 1 B 9 VPW nch L=4e-08 W=3.9e-07 
M8 10 B 1 VPW nch L=4e-08 W=3.9e-07 
M9 Y A 10 VPW nch L=4e-08 W=3.9e-07 
M10 11 A Y VPW nch L=4e-08 W=3.9e-07 
M11 1 B 11 VPW nch L=4e-08 W=3.9e-07 
M12 Y C VDD VNW pch L=4e-08 W=3.9e-07 
M13 VDD C Y VNW pch L=4e-08 W=3.9e-07 
M14 Y C VDD VNW pch L=4e-08 W=3.9e-07 
M15 VDD C Y VNW pch L=4e-08 W=3.9e-07 
M16 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M17 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M18 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M19 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M20 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M21 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M22 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M23 VDD B Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND3_X4M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=4e-07 
M1 1 C VSS VPW nch L=4e-08 W=4e-07 
M2 VSS C 1 VPW nch L=4e-08 W=4e-07 
M3 1 C VSS VPW nch L=4e-08 W=4e-07 
M4 8 B 1 VPW nch L=4e-08 W=4e-07 
M5 Y A 8 VPW nch L=4e-08 W=4e-07 
M6 9 A Y VPW nch L=4e-08 W=4e-07 
M7 1 B 9 VPW nch L=4e-08 W=4e-07 
M8 10 B 1 VPW nch L=4e-08 W=4e-07 
M9 Y A 10 VPW nch L=4e-08 W=4e-07 
M10 11 A Y VPW nch L=4e-08 W=4e-07 
M11 1 B 11 VPW nch L=4e-08 W=4e-07 
M12 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M13 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M14 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M15 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M16 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M17 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M18 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M19 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M20 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M21 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M22 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M23 VDD B Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND3_X6A_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=3.9e-07 
M1 1 C VSS VPW nch L=4e-08 W=3.9e-07 
M2 VSS C 1 VPW nch L=4e-08 W=3.9e-07 
M3 1 C VSS VPW nch L=4e-08 W=3.9e-07 
M4 VSS C 1 VPW nch L=4e-08 W=3.9e-07 
M5 1 C VSS VPW nch L=4e-08 W=3.9e-07 
M6 8 B 1 VPW nch L=4e-08 W=3.9e-07 
M7 Y A 8 VPW nch L=4e-08 W=3.9e-07 
M8 9 A Y VPW nch L=4e-08 W=3.9e-07 
M9 1 B 9 VPW nch L=4e-08 W=3.9e-07 
M10 10 B 1 VPW nch L=4e-08 W=3.9e-07 
M11 Y A 10 VPW nch L=4e-08 W=3.9e-07 
M12 11 A Y VPW nch L=4e-08 W=3.9e-07 
M13 1 B 11 VPW nch L=4e-08 W=3.9e-07 
M14 12 B 1 VPW nch L=4e-08 W=3.9e-07 
M15 Y A 12 VPW nch L=4e-08 W=3.9e-07 
M16 13 A Y VPW nch L=4e-08 W=3.9e-07 
M17 1 B 13 VPW nch L=4e-08 W=3.9e-07 
M18 Y C VDD VNW pch L=4e-08 W=3.9e-07 
M19 VDD C Y VNW pch L=4e-08 W=3.9e-07 
M20 Y C VDD VNW pch L=4e-08 W=3.9e-07 
M21 VDD C Y VNW pch L=4e-08 W=3.9e-07 
M22 Y C VDD VNW pch L=4e-08 W=3.9e-07 
M23 VDD C Y VNW pch L=4e-08 W=3.9e-07 
M24 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M25 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M26 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M27 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M28 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M29 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M30 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M31 VDD B Y VNW pch L=4e-08 W=3.9e-07 
M32 Y B VDD VNW pch L=4e-08 W=3.9e-07 
M33 VDD A Y VNW pch L=4e-08 W=3.9e-07 
M34 Y A VDD VNW pch L=4e-08 W=3.9e-07 
M35 VDD B Y VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NAND3_X6M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=4e-07 
M1 1 C VSS VPW nch L=4e-08 W=4e-07 
M2 VSS C 1 VPW nch L=4e-08 W=4e-07 
M3 1 C VSS VPW nch L=4e-08 W=4e-07 
M4 VSS C 1 VPW nch L=4e-08 W=4e-07 
M5 1 C VSS VPW nch L=4e-08 W=4e-07 
M6 8 B 1 VPW nch L=4e-08 W=4e-07 
M7 Y A 8 VPW nch L=4e-08 W=4e-07 
M8 9 A Y VPW nch L=4e-08 W=4e-07 
M9 1 B 9 VPW nch L=4e-08 W=4e-07 
M10 10 B 1 VPW nch L=4e-08 W=4e-07 
M11 Y A 10 VPW nch L=4e-08 W=4e-07 
M12 11 A Y VPW nch L=4e-08 W=4e-07 
M13 1 B 11 VPW nch L=4e-08 W=4e-07 
M14 12 B 1 VPW nch L=4e-08 W=4e-07 
M15 Y A 12 VPW nch L=4e-08 W=4e-07 
M16 13 A Y VPW nch L=4e-08 W=4e-07 
M17 1 B 13 VPW nch L=4e-08 W=4e-07 
M18 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M19 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M20 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M21 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M22 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M23 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M24 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M25 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M26 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M27 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M28 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M29 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M30 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M31 VDD B Y VNW pch L=4e-08 W=2.65e-07 
M32 Y B VDD VNW pch L=4e-08 W=2.65e-07 
M33 VDD A Y VNW pch L=4e-08 W=2.65e-07 
M34 Y A VDD VNW pch L=4e-08 W=2.65e-07 
M35 VDD B Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND4BB_X0P5M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 2 AN VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=1.2e-07 
M2 10 D VSS VPW nch L=4e-08 W=2e-07 
M3 11 C 10 VPW nch L=4e-08 W=2e-07 
M4 Y 2 11 VPW nch L=4e-08 W=2e-07 
M5 9 AN 2 VNW pch L=4e-08 W=2.1e-07 
M6 VDD BN 9 VNW pch L=4e-08 W=2.1e-07 
M7 Y D VDD VNW pch L=4e-08 W=1.35e-07 
M8 VDD C Y VNW pch L=4e-08 W=1.35e-07 
M9 Y 2 VDD VNW pch L=4e-08 W=1.35e-07 
.ENDS


.SUBCKT NAND4BB_X0P7M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 2 AN VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=1.2e-07 
M2 10 D VSS VPW nch L=4e-08 W=2.85e-07 
M3 11 C 10 VPW nch L=4e-08 W=2.85e-07 
M4 Y 2 11 VPW nch L=4e-08 W=2.85e-07 
M5 9 AN 2 VNW pch L=4e-08 W=2.95e-07 
M6 VDD BN 9 VNW pch L=4e-08 W=2.95e-07 
M7 Y D VDD VNW pch L=4e-08 W=1.9e-07 
M8 VDD C Y VNW pch L=4e-08 W=1.9e-07 
M9 Y 2 VDD VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT NAND4BB_X1M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 2 AN VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=1.2e-07 
M2 10 D VSS VPW nch L=4e-08 W=3.9e-07 
M3 11 C 10 VPW nch L=4e-08 W=3.9e-07 
M4 Y 2 11 VPW nch L=4e-08 W=3.9e-07 
M5 9 AN 2 VNW pch L=4e-08 W=3e-07 
M6 VDD BN 9 VNW pch L=4e-08 W=3e-07 
M7 Y D VDD VNW pch L=4e-08 W=2.65e-07 
M8 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M9 Y 2 VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND4BB_X1P4M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 2 AN VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=1.6e-07 
M2 10 D VSS VPW nch L=4e-08 W=2.85e-07 
M3 11 C 10 VPW nch L=4e-08 W=2.85e-07 
M4 Y 2 11 VPW nch L=4e-08 W=2.85e-07 
M5 12 2 Y VPW nch L=4e-08 W=2.85e-07 
M6 13 C 12 VPW nch L=4e-08 W=2.85e-07 
M7 VSS D 13 VPW nch L=4e-08 W=2.85e-07 
M8 9 AN 2 VNW pch L=4e-08 W=4e-07 
M9 VDD BN 9 VNW pch L=4e-08 W=4e-07 
M10 Y D VDD VNW pch L=4e-08 W=1.9e-07 
M11 VDD C Y VNW pch L=4e-08 W=1.9e-07 
M12 Y 2 VDD VNW pch L=4e-08 W=1.9e-07 
M13 VDD 2 Y VNW pch L=4e-08 W=1.9e-07 
M14 Y C VDD VNW pch L=4e-08 W=1.9e-07 
M15 VDD D Y VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT NAND4BB_X2M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 3 BN VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS AN 3 VPW nch L=4e-08 W=1.2e-07 
M2 3 AN VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS BN 3 VPW nch L=4e-08 W=1.2e-07 
M4 11 D VSS VPW nch L=4e-08 W=4e-07 
M5 12 C 11 VPW nch L=4e-08 W=4e-07 
M6 Y 3 12 VPW nch L=4e-08 W=4e-07 
M7 13 3 Y VPW nch L=4e-08 W=4e-07 
M8 14 C 13 VPW nch L=4e-08 W=4e-07 
M9 VSS D 14 VPW nch L=4e-08 W=4e-07 
M10 9 BN VDD VNW pch L=4e-08 W=2.95e-07 
M11 3 AN 9 VNW pch L=4e-08 W=2.95e-07 
M12 10 AN 3 VNW pch L=4e-08 W=2.95e-07 
M13 VDD BN 10 VNW pch L=4e-08 W=2.95e-07 
M14 Y D VDD VNW pch L=4e-08 W=2.65e-07 
M15 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M16 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M17 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M18 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M19 VDD D Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND4BB_X3M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 3 BN VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS AN 3 VPW nch L=4e-08 W=1.6e-07 
M2 3 AN VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS BN 3 VPW nch L=4e-08 W=1.6e-07 
M4 4 D VSS VPW nch L=4e-08 W=4e-07 
M5 VSS D 4 VPW nch L=4e-08 W=4e-07 
M6 4 D VSS VPW nch L=4e-08 W=4e-07 
M7 12 C 4 VPW nch L=4e-08 W=4e-07 
M8 Y 3 12 VPW nch L=4e-08 W=4e-07 
M9 13 3 Y VPW nch L=4e-08 W=4e-07 
M10 4 C 13 VPW nch L=4e-08 W=4e-07 
M11 14 C 4 VPW nch L=4e-08 W=4e-07 
M12 Y 3 14 VPW nch L=4e-08 W=4e-07 
M13 10 BN VDD VNW pch L=4e-08 W=4e-07 
M14 3 AN 10 VNW pch L=4e-08 W=4e-07 
M15 11 AN 3 VNW pch L=4e-08 W=4e-07 
M16 VDD BN 11 VNW pch L=4e-08 W=4e-07 
M17 Y D VDD VNW pch L=4e-08 W=2.65e-07 
M18 VDD D Y VNW pch L=4e-08 W=2.65e-07 
M19 Y D VDD VNW pch L=4e-08 W=2.65e-07 
M20 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M21 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M22 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M23 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M24 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M25 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND4BB_X4M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 2 AN VSS VPW nch L=4e-08 W=1.55e-07 
M1 VSS BN 2 VPW nch L=4e-08 W=1.55e-07 
M2 2 BN VSS VPW nch L=4e-08 W=1.55e-07 
M3 VSS AN 2 VPW nch L=4e-08 W=1.55e-07 
M4 2 AN VSS VPW nch L=4e-08 W=1.55e-07 
M5 VSS BN 2 VPW nch L=4e-08 W=1.55e-07 
M6 12 D VSS VPW nch L=4e-08 W=3.8e-07 
M7 13 C 12 VPW nch L=4e-08 W=3.8e-07 
M8 Y 2 13 VPW nch L=4e-08 W=3.8e-07 
M9 14 2 Y VPW nch L=4e-08 W=3.8e-07 
M10 15 C 14 VPW nch L=4e-08 W=3.8e-07 
M11 VSS D 15 VPW nch L=4e-08 W=3.8e-07 
M12 16 D VSS VPW nch L=4e-08 W=3.8e-07 
M13 17 C 16 VPW nch L=4e-08 W=3.8e-07 
M14 Y 2 17 VPW nch L=4e-08 W=3.8e-07 
M15 18 2 Y VPW nch L=4e-08 W=3.8e-07 
M16 19 C 18 VPW nch L=4e-08 W=3.8e-07 
M17 VSS D 19 VPW nch L=4e-08 W=3.8e-07 
M18 9 AN 2 VNW pch L=4e-08 W=3.8e-07 
M19 VDD BN 9 VNW pch L=4e-08 W=3.8e-07 
M20 10 BN VDD VNW pch L=4e-08 W=3.8e-07 
M21 2 AN 10 VNW pch L=4e-08 W=3.8e-07 
M22 11 AN 2 VNW pch L=4e-08 W=3.8e-07 
M23 VDD BN 11 VNW pch L=4e-08 W=3.8e-07 
M24 Y D VDD VNW pch L=4e-08 W=2.65e-07 
M25 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M26 Y 2 VDD VNW pch L=4e-08 W=2.65e-07 
M27 VDD 2 Y VNW pch L=4e-08 W=2.65e-07 
M28 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M29 VDD D Y VNW pch L=4e-08 W=2.65e-07 
M30 Y D VDD VNW pch L=4e-08 W=2.65e-07 
M31 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M32 Y 2 VDD VNW pch L=4e-08 W=2.65e-07 
M33 VDD 2 Y VNW pch L=4e-08 W=2.65e-07 
M34 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M35 VDD D Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND4BB_X6M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 3 BN VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS AN 3 VPW nch L=4e-08 W=1.6e-07 
M2 3 AN VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS BN 3 VPW nch L=4e-08 W=1.6e-07 
M4 3 BN VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS AN 3 VPW nch L=4e-08 W=1.6e-07 
M6 3 AN VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS BN 3 VPW nch L=4e-08 W=1.6e-07 
M8 13 D VSS VPW nch L=4e-08 W=3.8e-07 
M9 14 C 13 VPW nch L=4e-08 W=3.8e-07 
M10 Y 3 14 VPW nch L=4e-08 W=3.8e-07 
M11 15 3 Y VPW nch L=4e-08 W=3.8e-07 
M12 16 C 15 VPW nch L=4e-08 W=3.8e-07 
M13 VSS D 16 VPW nch L=4e-08 W=3.8e-07 
M14 17 D VSS VPW nch L=4e-08 W=3.8e-07 
M15 18 C 17 VPW nch L=4e-08 W=3.8e-07 
M16 Y 3 18 VPW nch L=4e-08 W=3.8e-07 
M17 19 3 Y VPW nch L=4e-08 W=3.8e-07 
M18 20 C 19 VPW nch L=4e-08 W=3.8e-07 
M19 VSS D 20 VPW nch L=4e-08 W=3.8e-07 
M20 21 D VSS VPW nch L=4e-08 W=3.8e-07 
M21 22 C 21 VPW nch L=4e-08 W=3.8e-07 
M22 Y 3 22 VPW nch L=4e-08 W=3.8e-07 
M23 23 3 Y VPW nch L=4e-08 W=3.8e-07 
M24 24 C 23 VPW nch L=4e-08 W=3.8e-07 
M25 VSS D 24 VPW nch L=4e-08 W=3.8e-07 
M26 9 BN VDD VNW pch L=4e-08 W=4e-07 
M27 3 AN 9 VNW pch L=4e-08 W=4e-07 
M28 10 AN 3 VNW pch L=4e-08 W=4e-07 
M29 VDD BN 10 VNW pch L=4e-08 W=4e-07 
M30 11 BN VDD VNW pch L=4e-08 W=4e-07 
M31 3 AN 11 VNW pch L=4e-08 W=4e-07 
M32 12 AN 3 VNW pch L=4e-08 W=4e-07 
M33 VDD BN 12 VNW pch L=4e-08 W=4e-07 
M34 Y D VDD VNW pch L=4e-08 W=2.65e-07 
M35 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M36 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M37 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M38 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M39 VDD D Y VNW pch L=4e-08 W=2.65e-07 
M40 Y D VDD VNW pch L=4e-08 W=2.65e-07 
M41 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M42 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M43 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M44 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M45 VDD D Y VNW pch L=4e-08 W=2.65e-07 
M46 Y D VDD VNW pch L=4e-08 W=2.65e-07 
M47 VDD C Y VNW pch L=4e-08 W=2.65e-07 
M48 Y 3 VDD VNW pch L=4e-08 W=2.65e-07 
M49 VDD 3 Y VNW pch L=4e-08 W=2.65e-07 
M50 Y C VDD VNW pch L=4e-08 W=2.65e-07 
M51 VDD D Y VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT NAND4B_X0P5M_A9TR Y VDD VNW VPW VSS AN B C D
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 9 D VSS VPW nch L=4e-08 W=2.25e-07 
M2 10 C 9 VPW nch L=4e-08 W=2.25e-07 
M3 11 B 10 VPW nch L=4e-08 W=2.25e-07 
M4 Y 1 11 VPW nch L=4e-08 W=2.25e-07 
M5 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M6 Y D VDD VNW pch L=4e-08 W=1.2e-07 
M7 VDD C Y VNW pch L=4e-08 W=1.2e-07 
M8 Y B VDD VNW pch L=4e-08 W=1.2e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT NAND4B_X0P7M_A9TR Y VDD VNW VPW VSS AN B C D
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 9 D VSS VPW nch L=4e-08 W=2.85e-07 
M2 10 C 9 VPW nch L=4e-08 W=2.85e-07 
M3 11 B 10 VPW nch L=4e-08 W=2.85e-07 
M4 Y 1 11 VPW nch L=4e-08 W=2.85e-07 
M5 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M6 Y D VDD VNW pch L=4e-08 W=1.55e-07 
M7 VDD C Y VNW pch L=4e-08 W=1.55e-07 
M8 Y B VDD VNW pch L=4e-08 W=1.55e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=1.55e-07 
.ENDS


.SUBCKT NAND4B_X1M_A9TR Y VDD VNW VPW VSS AN B C D
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 9 D VSS VPW nch L=4e-08 W=3.8e-07 
M2 10 C 9 VPW nch L=4e-08 W=3.8e-07 
M3 11 B 10 VPW nch L=4e-08 W=3.8e-07 
M4 Y 1 11 VPW nch L=4e-08 W=3.8e-07 
M5 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M6 Y D VDD VNW pch L=4e-08 W=2.15e-07 
M7 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M8 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M9 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
.ENDS


.SUBCKT NAND4B_X1P4M_A9TR Y VDD VNW VPW VSS AN B C D
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 10 C 4 VPW nch L=4e-08 W=2.85e-07 
M2 VSS D 10 VPW nch L=4e-08 W=2.85e-07 
M3 11 D VSS VPW nch L=4e-08 W=2.85e-07 
M4 4 C 11 VPW nch L=4e-08 W=2.85e-07 
M5 12 B 4 VPW nch L=4e-08 W=2.85e-07 
M6 Y 1 12 VPW nch L=4e-08 W=2.85e-07 
M7 13 1 Y VPW nch L=4e-08 W=2.85e-07 
M8 4 B 13 VPW nch L=4e-08 W=2.85e-07 
M9 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M10 Y C VDD VNW pch L=4e-08 W=1.55e-07 
M11 VDD D Y VNW pch L=4e-08 W=1.55e-07 
M12 Y D VDD VNW pch L=4e-08 W=1.55e-07 
M13 VDD C Y VNW pch L=4e-08 W=1.55e-07 
M14 Y B VDD VNW pch L=4e-08 W=1.55e-07 
M15 VDD 1 Y VNW pch L=4e-08 W=1.55e-07 
M16 Y 1 VDD VNW pch L=4e-08 W=1.55e-07 
M17 VDD B Y VNW pch L=4e-08 W=1.55e-07 
.ENDS


.SUBCKT NAND4B_X2M_A9TR Y VDD VNW VPW VSS AN B C D
M0 VSS AN 1 VPW nch L=4e-08 W=1.6e-07 
M1 10 C 4 VPW nch L=4e-08 W=4e-07 
M2 VSS D 10 VPW nch L=4e-08 W=4e-07 
M3 11 D VSS VPW nch L=4e-08 W=4e-07 
M4 4 C 11 VPW nch L=4e-08 W=4e-07 
M5 12 B 4 VPW nch L=4e-08 W=4e-07 
M6 Y 1 12 VPW nch L=4e-08 W=4e-07 
M7 13 1 Y VPW nch L=4e-08 W=4e-07 
M8 4 B 13 VPW nch L=4e-08 W=4e-07 
M9 VDD AN 1 VNW pch L=4e-08 W=2.05e-07 
M10 Y C VDD VNW pch L=4e-08 W=2.15e-07 
M11 VDD D Y VNW pch L=4e-08 W=2.15e-07 
M12 Y D VDD VNW pch L=4e-08 W=2.15e-07 
M13 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M14 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M15 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
M16 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M17 VDD B Y VNW pch L=4e-08 W=2.15e-07 
.ENDS


.SUBCKT NAND4B_X3M_A9TR Y VDD VNW VPW VSS AN B C D
M0 VSS AN 1 VPW nch L=4e-08 W=2.3e-07 
M1 10 D VSS VPW nch L=4e-08 W=4e-07 
M2 5 C 10 VPW nch L=4e-08 W=4e-07 
M3 11 C 5 VPW nch L=4e-08 W=4e-07 
M4 VSS D 11 VPW nch L=4e-08 W=4e-07 
M5 12 D VSS VPW nch L=4e-08 W=4e-07 
M6 5 C 12 VPW nch L=4e-08 W=4e-07 
M7 13 B 5 VPW nch L=4e-08 W=4e-07 
M8 Y 1 13 VPW nch L=4e-08 W=4e-07 
M9 14 1 Y VPW nch L=4e-08 W=4e-07 
M10 5 B 14 VPW nch L=4e-08 W=4e-07 
M11 15 B 5 VPW nch L=4e-08 W=4e-07 
M12 Y 1 15 VPW nch L=4e-08 W=4e-07 
M13 VDD AN 1 VNW pch L=4e-08 W=3e-07 
M14 Y D VDD VNW pch L=4e-08 W=2.15e-07 
M15 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M16 Y C VDD VNW pch L=4e-08 W=2.15e-07 
M17 VDD D Y VNW pch L=4e-08 W=2.15e-07 
M18 Y D VDD VNW pch L=4e-08 W=2.15e-07 
M19 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M20 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M21 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M23 VDD B Y VNW pch L=4e-08 W=2.15e-07 
M24 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M25 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
.ENDS


.SUBCKT NAND4B_X4M_A9TR Y VDD VNW VPW VSS AN B C D
M0 VSS AN 1 VPW nch L=4e-08 W=3.05e-07 
M1 10 C 4 VPW nch L=4e-08 W=4e-07 
M2 VSS D 10 VPW nch L=4e-08 W=4e-07 
M3 11 D VSS VPW nch L=4e-08 W=4e-07 
M4 4 C 11 VPW nch L=4e-08 W=4e-07 
M5 12 C 4 VPW nch L=4e-08 W=4e-07 
M6 VSS D 12 VPW nch L=4e-08 W=4e-07 
M7 13 D VSS VPW nch L=4e-08 W=4e-07 
M8 4 C 13 VPW nch L=4e-08 W=4e-07 
M9 14 B 4 VPW nch L=4e-08 W=4e-07 
M10 Y 1 14 VPW nch L=4e-08 W=4e-07 
M11 15 1 Y VPW nch L=4e-08 W=4e-07 
M12 4 B 15 VPW nch L=4e-08 W=4e-07 
M13 16 B 4 VPW nch L=4e-08 W=4e-07 
M14 Y 1 16 VPW nch L=4e-08 W=4e-07 
M15 17 1 Y VPW nch L=4e-08 W=4e-07 
M16 4 B 17 VPW nch L=4e-08 W=4e-07 
M17 VDD AN 1 VNW pch L=4e-08 W=3.95e-07 
M18 Y C VDD VNW pch L=4e-08 W=2.15e-07 
M19 VDD D Y VNW pch L=4e-08 W=2.15e-07 
M20 Y D VDD VNW pch L=4e-08 W=2.15e-07 
M21 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M22 Y C VDD VNW pch L=4e-08 W=2.15e-07 
M23 VDD D Y VNW pch L=4e-08 W=2.15e-07 
M24 Y D VDD VNW pch L=4e-08 W=2.15e-07 
M25 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M26 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M27 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
M28 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M29 VDD B Y VNW pch L=4e-08 W=2.15e-07 
M30 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M31 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
M32 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M33 VDD B Y VNW pch L=4e-08 W=2.15e-07 
.ENDS


.SUBCKT NAND4XXXB_X0P5M_A9TR Y VDD VNW VPW VSS A B C DN
M0 VSS DN 1 VPW nch L=4e-08 W=1.2e-07 
M1 9 1 VSS VPW nch L=4e-08 W=2.25e-07 
M2 10 C 9 VPW nch L=4e-08 W=2.25e-07 
M3 11 B 10 VPW nch L=4e-08 W=2.25e-07 
M4 Y A 11 VPW nch L=4e-08 W=2.25e-07 
M5 VDD DN 1 VNW pch L=4e-08 W=1.55e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=1.2e-07 
M7 VDD C Y VNW pch L=4e-08 W=1.2e-07 
M8 Y B VDD VNW pch L=4e-08 W=1.2e-07 
M9 VDD A Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT NAND4XXXB_X0P7M_A9TR Y VDD VNW VPW VSS A B C DN
M0 VSS DN 1 VPW nch L=4e-08 W=1.2e-07 
M1 9 1 VSS VPW nch L=4e-08 W=2.85e-07 
M2 10 C 9 VPW nch L=4e-08 W=2.85e-07 
M3 11 B 10 VPW nch L=4e-08 W=2.85e-07 
M4 Y A 11 VPW nch L=4e-08 W=2.85e-07 
M5 VDD DN 1 VNW pch L=4e-08 W=1.55e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=1.55e-07 
M7 VDD C Y VNW pch L=4e-08 W=1.55e-07 
M8 Y B VDD VNW pch L=4e-08 W=1.55e-07 
M9 VDD A Y VNW pch L=4e-08 W=1.55e-07 
.ENDS


.SUBCKT NAND4XXXB_X1M_A9TR Y VDD VNW VPW VSS A B C DN
M0 VSS DN 1 VPW nch L=4e-08 W=1.2e-07 
M1 9 1 VSS VPW nch L=4e-08 W=4e-07 
M2 10 C 9 VPW nch L=4e-08 W=4e-07 
M3 11 B 10 VPW nch L=4e-08 W=4e-07 
M4 Y A 11 VPW nch L=4e-08 W=4e-07 
M5 VDD DN 1 VNW pch L=4e-08 W=1.55e-07 
M6 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M7 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M8 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M9 VDD A Y VNW pch L=4e-08 W=2.15e-07 
.ENDS


.SUBCKT NAND4XXXB_X1P4M_A9TR Y VDD VNW VPW VSS A B C DN
M0 VSS DN 1 VPW nch L=4e-08 W=1.2e-07 
M1 10 C 4 VPW nch L=4e-08 W=2.85e-07 
M2 VSS 1 10 VPW nch L=4e-08 W=2.85e-07 
M3 11 1 VSS VPW nch L=4e-08 W=2.85e-07 
M4 4 C 11 VPW nch L=4e-08 W=2.85e-07 
M5 12 B 4 VPW nch L=4e-08 W=2.85e-07 
M6 Y A 12 VPW nch L=4e-08 W=2.85e-07 
M7 13 A Y VPW nch L=4e-08 W=2.85e-07 
M8 4 B 13 VPW nch L=4e-08 W=2.85e-07 
M9 VDD DN 1 VNW pch L=4e-08 W=1.55e-07 
M10 Y C VDD VNW pch L=4e-08 W=1.55e-07 
M11 VDD 1 Y VNW pch L=4e-08 W=1.55e-07 
M12 Y 1 VDD VNW pch L=4e-08 W=1.55e-07 
M13 VDD C Y VNW pch L=4e-08 W=1.55e-07 
M14 Y B VDD VNW pch L=4e-08 W=1.55e-07 
M15 VDD A Y VNW pch L=4e-08 W=1.55e-07 
M16 Y A VDD VNW pch L=4e-08 W=1.55e-07 
M17 VDD B Y VNW pch L=4e-08 W=1.55e-07 
.ENDS


.SUBCKT NAND4XXXB_X2M_A9TR Y VDD VNW VPW VSS A B C DN
M0 VSS DN 1 VPW nch L=4e-08 W=1.6e-07 
M1 10 C 4 VPW nch L=4e-08 W=4e-07 
M2 VSS 1 10 VPW nch L=4e-08 W=4e-07 
M3 11 1 VSS VPW nch L=4e-08 W=4e-07 
M4 4 C 11 VPW nch L=4e-08 W=4e-07 
M5 12 B 4 VPW nch L=4e-08 W=4e-07 
M6 Y A 12 VPW nch L=4e-08 W=4e-07 
M7 13 A Y VPW nch L=4e-08 W=4e-07 
M8 4 B 13 VPW nch L=4e-08 W=4e-07 
M9 VDD DN 1 VNW pch L=4e-08 W=2.05e-07 
M10 Y C VDD VNW pch L=4e-08 W=2.15e-07 
M11 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
M12 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M13 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M14 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M15 VDD A Y VNW pch L=4e-08 W=2.15e-07 
M16 Y A VDD VNW pch L=4e-08 W=2.15e-07 
M17 VDD B Y VNW pch L=4e-08 W=2.15e-07 
.ENDS


.SUBCKT NAND4XXXB_X3M_A9TR Y VDD VNW VPW VSS A B C DN
M0 VSS DN 1 VPW nch L=4e-08 W=2.3e-07 
M1 10 1 VSS VPW nch L=4e-08 W=4e-07 
M2 5 C 10 VPW nch L=4e-08 W=4e-07 
M3 11 C 5 VPW nch L=4e-08 W=4e-07 
M4 VSS 1 11 VPW nch L=4e-08 W=4e-07 
M5 12 1 VSS VPW nch L=4e-08 W=4e-07 
M6 5 C 12 VPW nch L=4e-08 W=4e-07 
M7 13 B 5 VPW nch L=4e-08 W=4e-07 
M8 Y A 13 VPW nch L=4e-08 W=4e-07 
M9 14 A Y VPW nch L=4e-08 W=4e-07 
M10 5 B 14 VPW nch L=4e-08 W=4e-07 
M11 15 B 5 VPW nch L=4e-08 W=4e-07 
M12 Y A 15 VPW nch L=4e-08 W=4e-07 
M13 VDD DN 1 VNW pch L=4e-08 W=3e-07 
M14 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M15 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M16 Y C VDD VNW pch L=4e-08 W=2.15e-07 
M17 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
M18 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M19 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M20 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M21 VDD A Y VNW pch L=4e-08 W=2.15e-07 
M22 Y A VDD VNW pch L=4e-08 W=2.15e-07 
M23 VDD B Y VNW pch L=4e-08 W=2.15e-07 
M24 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M25 VDD A Y VNW pch L=4e-08 W=2.15e-07 
.ENDS


.SUBCKT NAND4XXXB_X4M_A9TR Y VDD VNW VPW VSS A B C DN
M0 VSS DN 1 VPW nch L=4e-08 W=3.05e-07 
M1 10 C 4 VPW nch L=4e-08 W=4e-07 
M2 VSS 1 10 VPW nch L=4e-08 W=4e-07 
M3 11 1 VSS VPW nch L=4e-08 W=4e-07 
M4 4 C 11 VPW nch L=4e-08 W=4e-07 
M5 12 C 4 VPW nch L=4e-08 W=4e-07 
M6 VSS 1 12 VPW nch L=4e-08 W=4e-07 
M7 13 1 VSS VPW nch L=4e-08 W=4e-07 
M8 4 C 13 VPW nch L=4e-08 W=4e-07 
M9 14 B 4 VPW nch L=4e-08 W=4e-07 
M10 Y A 14 VPW nch L=4e-08 W=4e-07 
M11 15 A Y VPW nch L=4e-08 W=4e-07 
M12 4 B 15 VPW nch L=4e-08 W=4e-07 
M13 16 B 4 VPW nch L=4e-08 W=4e-07 
M14 Y A 16 VPW nch L=4e-08 W=4e-07 
M15 17 A Y VPW nch L=4e-08 W=4e-07 
M16 4 B 17 VPW nch L=4e-08 W=4e-07 
M17 VDD DN 1 VNW pch L=4e-08 W=3.95e-07 
M18 Y C VDD VNW pch L=4e-08 W=2.15e-07 
M19 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
M20 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M21 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M22 Y C VDD VNW pch L=4e-08 W=2.15e-07 
M23 VDD 1 Y VNW pch L=4e-08 W=2.15e-07 
M24 Y 1 VDD VNW pch L=4e-08 W=2.15e-07 
M25 VDD C Y VNW pch L=4e-08 W=2.15e-07 
M26 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M27 VDD A Y VNW pch L=4e-08 W=2.15e-07 
M28 Y A VDD VNW pch L=4e-08 W=2.15e-07 
M29 VDD B Y VNW pch L=4e-08 W=2.15e-07 
M30 Y B VDD VNW pch L=4e-08 W=2.15e-07 
M31 VDD A Y VNW pch L=4e-08 W=2.15e-07 
M32 Y A VDD VNW pch L=4e-08 W=2.15e-07 
M33 VDD B Y VNW pch L=4e-08 W=2.15e-07 
.ENDS


.SUBCKT NAND4_X0P5A_A9TR Y VDD VNW VPW VSS A B C D
M0 8 D VSS VPW nch L=4e-08 W=2e-07 
M1 9 C 8 VPW nch L=4e-08 W=2e-07 
M2 10 B 9 VPW nch L=4e-08 W=2e-07 
M3 Y A 10 VPW nch L=4e-08 W=2e-07 
M4 Y D VDD VNW pch L=4e-08 W=1.7e-07 
M5 VDD C Y VNW pch L=4e-08 W=1.7e-07 
M6 Y B VDD VNW pch L=4e-08 W=1.7e-07 
M7 VDD A Y VNW pch L=4e-08 W=1.7e-07 
.ENDS


.SUBCKT NAND4_X0P5M_A9TR Y VDD VNW VPW VSS A B C D
M0 8 D VSS VPW nch L=4e-08 W=2.25e-07 
M1 9 C 8 VPW nch L=4e-08 W=2.25e-07 
M2 10 B 9 VPW nch L=4e-08 W=2.25e-07 
M3 Y A 10 VPW nch L=4e-08 W=2.25e-07 
M4 Y D VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD C Y VNW pch L=4e-08 W=1.2e-07 
M6 Y B VDD VNW pch L=4e-08 W=1.2e-07 
M7 VDD A Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT NAND4_X0P7A_A9TR Y VDD VNW VPW VSS A B C D
M0 8 D VSS VPW nch L=4e-08 W=2.85e-07 
M1 9 C 8 VPW nch L=4e-08 W=2.85e-07 
M2 10 B 9 VPW nch L=4e-08 W=2.85e-07 
M3 Y A 10 VPW nch L=4e-08 W=2.85e-07 
M4 Y D VDD VNW pch L=4e-08 W=2.4e-07 
M5 VDD C Y VNW pch L=4e-08 W=2.4e-07 
M6 Y B VDD VNW pch L=4e-08 W=2.4e-07 
M7 VDD A Y VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT NAND4_X0P7M_A9TR Y VDD VNW VPW VSS A B C D
M0 8 D VSS VPW nch L=4e-08 W=2.85e-07 
M1 9 C 8 VPW nch L=4e-08 W=2.85e-07 
M2 10 B 9 VPW nch L=4e-08 W=2.85e-07 
M3 Y A 10 VPW nch L=4e-08 W=2.85e-07 
M4 Y D VDD VNW pch L=4e-08 W=1.55e-07 
M5 VDD C Y VNW pch L=4e-08 W=1.55e-07 
M6 Y B VDD VNW pch L=4e-08 W=1.55e-07 
M7 VDD A Y VNW pch L=4e-08 W=1.55e-07 
.ENDS


.SUBCKT NAND4_X1A_A9TR Y VDD VNW VPW VSS A B C D
M0 8 D VSS VPW nch L=4e-08 W=4e-07 
M1 9 C 8 VPW nch L=4e-08 W=4e-07 
M2 10 B 9 VPW nch L=4e-08 W=4e-07 
M3 Y A 10 VPW nch L=4e-08 W=4e-07 
M4 Y D VDD VNW pch L=4e-08 W=3.35e-07 
M5 VDD C Y VNW pch L=4e-08 W=3.35e-07 
M6 Y B VDD VNW pch L=4e-08 W=3.35e-07 
M7 VDD A Y VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT NAND4_X1M_A9TR Y VDD VNW VPW VSS A B C D
M0 8 D VSS VPW nch L=4e-08 W=4e-07 
M1 9 C 8 VPW nch L=4e-08 W=4e-07 
M2 10 B 9 VPW nch L=4e-08 W=4e-07 
M3 Y A 10 VPW nch L=4e-08 W=4e-07 
M4 Y D VDD VNW pch L=4e-08 W=2.2e-07 
M5 VDD C Y VNW pch L=4e-08 W=2.2e-07 
M6 Y B VDD VNW pch L=4e-08 W=2.2e-07 
M7 VDD A Y VNW pch L=4e-08 W=2.2e-07 
.ENDS


.SUBCKT NAND4_X1P4A_A9TR Y VDD VNW VPW VSS A B C D
M0 9 C 1 VPW nch L=4e-08 W=2.85e-07 
M1 VSS D 9 VPW nch L=4e-08 W=2.85e-07 
M2 10 D VSS VPW nch L=4e-08 W=2.85e-07 
M3 1 C 10 VPW nch L=4e-08 W=2.85e-07 
M4 11 B 1 VPW nch L=4e-08 W=2.85e-07 
M5 Y A 11 VPW nch L=4e-08 W=2.85e-07 
M6 12 A Y VPW nch L=4e-08 W=2.85e-07 
M7 1 B 12 VPW nch L=4e-08 W=2.85e-07 
M8 Y C VDD VNW pch L=4e-08 W=2.4e-07 
M9 VDD D Y VNW pch L=4e-08 W=2.4e-07 
M10 Y D VDD VNW pch L=4e-08 W=2.4e-07 
M11 VDD C Y VNW pch L=4e-08 W=2.4e-07 
M12 Y B VDD VNW pch L=4e-08 W=2.4e-07 
M13 VDD A Y VNW pch L=4e-08 W=2.4e-07 
M14 Y A VDD VNW pch L=4e-08 W=2.4e-07 
M15 VDD B Y VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT NAND4_X1P4M_A9TR Y VDD VNW VPW VSS A B C D
M0 11 C 1 VPW nch L=4e-08 W=2.85e-07 
M1 VSS D 11 VPW nch L=4e-08 W=2.85e-07 
M2 12 D VSS VPW nch L=4e-08 W=2.85e-07 
M3 1 C 12 VPW nch L=4e-08 W=2.85e-07 
M4 13 B 1 VPW nch L=4e-08 W=2.85e-07 
M5 Y A 13 VPW nch L=4e-08 W=2.85e-07 
M6 14 A Y VPW nch L=4e-08 W=2.85e-07 
M7 1 B 14 VPW nch L=4e-08 W=2.85e-07 
M8 Y D VDD VNW pch L=4e-08 W=3.1e-07 
M9 VDD C Y VNW pch L=4e-08 W=3.1e-07 
M10 Y B VDD VNW pch L=4e-08 W=3.1e-07 
M11 VDD A Y VNW pch L=4e-08 W=3.1e-07 
.ENDS


.SUBCKT NAND4_X2A_A9TR Y VDD VNW VPW VSS A B C D
M0 9 C 1 VPW nch L=4e-08 W=4e-07 
M1 VSS D 9 VPW nch L=4e-08 W=4e-07 
M2 10 D VSS VPW nch L=4e-08 W=4e-07 
M3 1 C 10 VPW nch L=4e-08 W=4e-07 
M4 11 B 1 VPW nch L=4e-08 W=4e-07 
M5 Y A 11 VPW nch L=4e-08 W=4e-07 
M6 12 A Y VPW nch L=4e-08 W=4e-07 
M7 1 B 12 VPW nch L=4e-08 W=4e-07 
M8 Y C VDD VNW pch L=4e-08 W=3.35e-07 
M9 VDD D Y VNW pch L=4e-08 W=3.35e-07 
M10 Y D VDD VNW pch L=4e-08 W=3.35e-07 
M11 VDD C Y VNW pch L=4e-08 W=3.35e-07 
M12 Y B VDD VNW pch L=4e-08 W=3.35e-07 
M13 VDD A Y VNW pch L=4e-08 W=3.35e-07 
M14 Y A VDD VNW pch L=4e-08 W=3.35e-07 
M15 VDD B Y VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT NAND4_X2M_A9TR Y VDD VNW VPW VSS A B C D
M0 9 C 1 VPW nch L=4e-08 W=4e-07 
M1 VSS D 9 VPW nch L=4e-08 W=4e-07 
M2 10 D VSS VPW nch L=4e-08 W=4e-07 
M3 1 C 10 VPW nch L=4e-08 W=4e-07 
M4 11 B 1 VPW nch L=4e-08 W=4e-07 
M5 Y A 11 VPW nch L=4e-08 W=4e-07 
M6 12 A Y VPW nch L=4e-08 W=4e-07 
M7 1 B 12 VPW nch L=4e-08 W=4e-07 
M8 Y C VDD VNW pch L=4e-08 W=2.2e-07 
M9 VDD D Y VNW pch L=4e-08 W=2.2e-07 
M10 Y D VDD VNW pch L=4e-08 W=2.2e-07 
M11 VDD C Y VNW pch L=4e-08 W=2.2e-07 
M12 Y B VDD VNW pch L=4e-08 W=2.2e-07 
M13 VDD A Y VNW pch L=4e-08 W=2.2e-07 
M14 Y A VDD VNW pch L=4e-08 W=2.2e-07 
M15 VDD B Y VNW pch L=4e-08 W=2.2e-07 
.ENDS


.SUBCKT NAND4_X3A_A9TR Y VDD VNW VPW VSS A B C D
M0 9 D VSS VPW nch L=4e-08 W=4e-07 
M1 4 C 9 VPW nch L=4e-08 W=4e-07 
M2 10 C 4 VPW nch L=4e-08 W=4e-07 
M3 VSS D 10 VPW nch L=4e-08 W=4e-07 
M4 11 D VSS VPW nch L=4e-08 W=4e-07 
M5 4 C 11 VPW nch L=4e-08 W=4e-07 
M6 12 B 4 VPW nch L=4e-08 W=4e-07 
M7 Y A 12 VPW nch L=4e-08 W=4e-07 
M8 13 A Y VPW nch L=4e-08 W=4e-07 
M9 4 B 13 VPW nch L=4e-08 W=4e-07 
M10 14 B 4 VPW nch L=4e-08 W=4e-07 
M11 Y A 14 VPW nch L=4e-08 W=4e-07 
M12 Y D VDD VNW pch L=4e-08 W=3.35e-07 
M13 VDD C Y VNW pch L=4e-08 W=3.35e-07 
M14 Y C VDD VNW pch L=4e-08 W=3.35e-07 
M15 VDD D Y VNW pch L=4e-08 W=3.35e-07 
M16 Y D VDD VNW pch L=4e-08 W=3.35e-07 
M17 VDD C Y VNW pch L=4e-08 W=3.35e-07 
M18 Y B VDD VNW pch L=4e-08 W=3.35e-07 
M19 VDD A Y VNW pch L=4e-08 W=3.35e-07 
M20 Y A VDD VNW pch L=4e-08 W=3.35e-07 
M21 VDD B Y VNW pch L=4e-08 W=3.35e-07 
M22 Y B VDD VNW pch L=4e-08 W=3.35e-07 
M23 VDD A Y VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT NAND4_X3M_A9TR Y VDD VNW VPW VSS A B C D
M0 11 D VSS VPW nch L=4e-08 W=4e-07 
M1 2 C 11 VPW nch L=4e-08 W=4e-07 
M2 12 C 2 VPW nch L=4e-08 W=4e-07 
M3 VSS D 12 VPW nch L=4e-08 W=4e-07 
M4 13 D VSS VPW nch L=4e-08 W=4e-07 
M5 2 C 13 VPW nch L=4e-08 W=4e-07 
M6 14 B 2 VPW nch L=4e-08 W=4e-07 
M7 Y A 14 VPW nch L=4e-08 W=4e-07 
M8 15 A Y VPW nch L=4e-08 W=4e-07 
M9 2 B 15 VPW nch L=4e-08 W=4e-07 
M10 16 B 2 VPW nch L=4e-08 W=4e-07 
M11 Y A 16 VPW nch L=4e-08 W=4e-07 
M12 Y C VDD VNW pch L=4e-08 W=3.25e-07 
M13 VDD D Y VNW pch L=4e-08 W=3.25e-07 
M14 Y D VDD VNW pch L=4e-08 W=3.25e-07 
M15 VDD C Y VNW pch L=4e-08 W=3.25e-07 
M16 Y B VDD VNW pch L=4e-08 W=3.25e-07 
M17 VDD A Y VNW pch L=4e-08 W=3.25e-07 
M18 Y A VDD VNW pch L=4e-08 W=3.25e-07 
M19 VDD B Y VNW pch L=4e-08 W=3.25e-07 
.ENDS


.SUBCKT NAND4_X4A_A9TR Y VDD VNW VPW VSS A B C D
M0 9 C 1 VPW nch L=4e-08 W=4e-07 
M1 VSS D 9 VPW nch L=4e-08 W=4e-07 
M2 10 D VSS VPW nch L=4e-08 W=4e-07 
M3 1 C 10 VPW nch L=4e-08 W=4e-07 
M4 11 C 1 VPW nch L=4e-08 W=4e-07 
M5 VSS D 11 VPW nch L=4e-08 W=4e-07 
M6 12 D VSS VPW nch L=4e-08 W=4e-07 
M7 1 C 12 VPW nch L=4e-08 W=4e-07 
M8 13 B 1 VPW nch L=4e-08 W=4e-07 
M9 Y A 13 VPW nch L=4e-08 W=4e-07 
M10 14 A Y VPW nch L=4e-08 W=4e-07 
M11 1 B 14 VPW nch L=4e-08 W=4e-07 
M12 15 B 1 VPW nch L=4e-08 W=4e-07 
M13 Y A 15 VPW nch L=4e-08 W=4e-07 
M14 16 A Y VPW nch L=4e-08 W=4e-07 
M15 1 B 16 VPW nch L=4e-08 W=4e-07 
M16 Y C VDD VNW pch L=4e-08 W=3.35e-07 
M17 VDD D Y VNW pch L=4e-08 W=3.35e-07 
M18 Y D VDD VNW pch L=4e-08 W=3.35e-07 
M19 VDD C Y VNW pch L=4e-08 W=3.35e-07 
M20 Y C VDD VNW pch L=4e-08 W=3.35e-07 
M21 VDD D Y VNW pch L=4e-08 W=3.35e-07 
M22 Y D VDD VNW pch L=4e-08 W=3.35e-07 
M23 VDD C Y VNW pch L=4e-08 W=3.35e-07 
M24 Y B VDD VNW pch L=4e-08 W=3.35e-07 
M25 VDD A Y VNW pch L=4e-08 W=3.35e-07 
M26 Y A VDD VNW pch L=4e-08 W=3.35e-07 
M27 VDD B Y VNW pch L=4e-08 W=3.35e-07 
M28 Y B VDD VNW pch L=4e-08 W=3.35e-07 
M29 VDD A Y VNW pch L=4e-08 W=3.35e-07 
M30 Y A VDD VNW pch L=4e-08 W=3.35e-07 
M31 VDD B Y VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT NAND4_X4M_A9TR Y VDD VNW VPW VSS A B C D
M0 11 C 1 VPW nch L=4e-08 W=4e-07 
M1 VSS D 11 VPW nch L=4e-08 W=4e-07 
M2 12 D VSS VPW nch L=4e-08 W=4e-07 
M3 1 C 12 VPW nch L=4e-08 W=4e-07 
M4 13 C 1 VPW nch L=4e-08 W=4e-07 
M5 VSS D 13 VPW nch L=4e-08 W=4e-07 
M6 14 D VSS VPW nch L=4e-08 W=4e-07 
M7 1 C 14 VPW nch L=4e-08 W=4e-07 
M8 15 B 1 VPW nch L=4e-08 W=4e-07 
M9 Y A 15 VPW nch L=4e-08 W=4e-07 
M10 16 A Y VPW nch L=4e-08 W=4e-07 
M11 1 B 16 VPW nch L=4e-08 W=4e-07 
M12 17 B 1 VPW nch L=4e-08 W=4e-07 
M13 Y A 17 VPW nch L=4e-08 W=4e-07 
M14 18 A Y VPW nch L=4e-08 W=4e-07 
M15 1 B 18 VPW nch L=4e-08 W=4e-07 
M16 Y D VDD VNW pch L=4e-08 W=2.9e-07 
M17 VDD C Y VNW pch L=4e-08 W=2.9e-07 
M18 Y C VDD VNW pch L=4e-08 W=2.9e-07 
M19 VDD D Y VNW pch L=4e-08 W=2.9e-07 
M20 Y D VDD VNW pch L=4e-08 W=2.9e-07 
M21 VDD C Y VNW pch L=4e-08 W=2.9e-07 
M22 Y B VDD VNW pch L=4e-08 W=2.9e-07 
M23 VDD A Y VNW pch L=4e-08 W=2.9e-07 
M24 Y A VDD VNW pch L=4e-08 W=2.9e-07 
M25 VDD B Y VNW pch L=4e-08 W=2.9e-07 
M26 Y B VDD VNW pch L=4e-08 W=2.9e-07 
M27 VDD A Y VNW pch L=4e-08 W=2.9e-07 
.ENDS


.SUBCKT NOR2B_X0P5M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y B VSS VPW nch L=4e-08 W=1.2e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=1.2e-07 
M3 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M4 7 B VDD VNW pch L=4e-08 W=2e-07 
M5 Y 1 7 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT NOR2B_X0P7M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y B VSS VPW nch L=4e-08 W=1.2e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=1.2e-07 
M3 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M4 7 B VDD VNW pch L=4e-08 W=2.95e-07 
M5 Y 1 7 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT NOR2B_X1M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y B VSS VPW nch L=4e-08 W=1.6e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M3 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M4 7 B VDD VNW pch L=4e-08 W=4e-07 
M5 Y 1 7 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2B_X1P4M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.3e-07 
M2 VSS B Y VPW nch L=4e-08 W=2.3e-07 
M3 VDD AN 1 VNW pch L=4e-08 W=1.55e-07 
M4 7 B VDD VNW pch L=4e-08 W=2.85e-07 
M5 Y 1 7 VNW pch L=4e-08 W=2.85e-07 
M6 8 1 Y VNW pch L=4e-08 W=2.85e-07 
M7 VDD B 8 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR2B_X2M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=1.45e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=3.2e-07 
M2 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M3 VDD AN 1 VNW pch L=4e-08 W=1.9e-07 
M4 7 B VDD VNW pch L=4e-08 W=4e-07 
M5 Y 1 7 VNW pch L=4e-08 W=4e-07 
M6 8 1 Y VNW pch L=4e-08 W=4e-07 
M7 VDD B 8 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2B_X3M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=2.15e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS B Y VPW nch L=4e-08 W=2.4e-07 
M3 Y B VSS VPW nch L=4e-08 W=2.4e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=2.4e-07 
M5 VDD AN 1 VNW pch L=4e-08 W=2.75e-07 
M6 7 B VDD VNW pch L=4e-08 W=4e-07 
M7 Y 1 7 VNW pch L=4e-08 W=4e-07 
M8 8 1 Y VNW pch L=4e-08 W=4e-07 
M9 VDD B 8 VNW pch L=4e-08 W=4e-07 
M10 9 B VDD VNW pch L=4e-08 W=4e-07 
M11 Y 1 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2B_X4M_A9TR Y VDD VNW VPW VSS AN B
M0 VSS AN 1 VPW nch L=4e-08 W=2.8e-07 
M1 Y B VSS VPW nch L=4e-08 W=3.2e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=3.2e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=3.2e-07 
M4 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M5 VDD AN 1 VNW pch L=4e-08 W=3.6e-07 
M6 7 B VDD VNW pch L=4e-08 W=4e-07 
M7 Y 1 7 VNW pch L=4e-08 W=4e-07 
M8 8 1 Y VNW pch L=4e-08 W=4e-07 
M9 VDD B 8 VNW pch L=4e-08 W=4e-07 
M10 9 B VDD VNW pch L=4e-08 W=4e-07 
M11 Y 1 9 VNW pch L=4e-08 W=4e-07 
M12 10 1 Y VNW pch L=4e-08 W=4e-07 
M13 VDD B 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2B_X6M_A9TR Y VDD VNW VPW VSS AN B
M0 3 AN VSS VPW nch L=4e-08 W=2.1e-07 
M1 VSS AN 3 VPW nch L=4e-08 W=2.1e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M4 Y B VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M7 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M8 3 AN VDD VNW pch L=4e-08 W=2.75e-07 
M9 VDD AN 3 VNW pch L=4e-08 W=2.75e-07 
M10 7 B VDD VNW pch L=4e-08 W=4e-07 
M11 Y 3 7 VNW pch L=4e-08 W=4e-07 
M12 8 3 Y VNW pch L=4e-08 W=4e-07 
M13 VDD B 8 VNW pch L=4e-08 W=4e-07 
M14 9 B VDD VNW pch L=4e-08 W=4e-07 
M15 Y 3 9 VNW pch L=4e-08 W=4e-07 
M16 10 3 Y VNW pch L=4e-08 W=4e-07 
M17 VDD B 10 VNW pch L=4e-08 W=4e-07 
M18 11 B VDD VNW pch L=4e-08 W=4e-07 
M19 Y 3 11 VNW pch L=4e-08 W=4e-07 
M20 12 3 Y VNW pch L=4e-08 W=4e-07 
M21 VDD B 12 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2B_X8M_A9TR Y VDD VNW VPW VSS AN B
M0 3 AN VSS VPW nch L=4e-08 W=2.8e-07 
M1 VSS AN 3 VPW nch L=4e-08 W=2.8e-07 
M2 Y B VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M6 Y B VSS VPW nch L=4e-08 W=3.2e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M9 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M10 3 AN VDD VNW pch L=4e-08 W=3.6e-07 
M11 VDD AN 3 VNW pch L=4e-08 W=3.6e-07 
M12 7 B VDD VNW pch L=4e-08 W=4e-07 
M13 Y 3 7 VNW pch L=4e-08 W=4e-07 
M14 8 3 Y VNW pch L=4e-08 W=4e-07 
M15 VDD B 8 VNW pch L=4e-08 W=4e-07 
M16 9 B VDD VNW pch L=4e-08 W=4e-07 
M17 Y 3 9 VNW pch L=4e-08 W=4e-07 
M18 10 3 Y VNW pch L=4e-08 W=4e-07 
M19 VDD B 10 VNW pch L=4e-08 W=4e-07 
M20 11 B VDD VNW pch L=4e-08 W=4e-07 
M21 Y 3 11 VNW pch L=4e-08 W=4e-07 
M22 12 3 Y VNW pch L=4e-08 W=4e-07 
M23 VDD B 12 VNW pch L=4e-08 W=4e-07 
M24 13 B VDD VNW pch L=4e-08 W=4e-07 
M25 Y 3 13 VNW pch L=4e-08 W=4e-07 
M26 14 3 Y VNW pch L=4e-08 W=4e-07 
M27 VDD B 14 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2XB_X0P5M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 VSS A Y VPW nch L=4e-08 W=1.2e-07 
M3 VDD BN 1 VNW pch L=4e-08 W=1.55e-07 
M4 7 1 VDD VNW pch L=4e-08 W=2e-07 
M5 Y A 7 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT NOR2XB_X0P7M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 VSS A Y VPW nch L=4e-08 W=1.2e-07 
M3 VDD BN 1 VNW pch L=4e-08 W=1.55e-07 
M4 7 1 VDD VNW pch L=4e-08 W=2.95e-07 
M5 Y A 7 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT NOR2XB_X1M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M2 VSS A Y VPW nch L=4e-08 W=1.6e-07 
M3 VDD BN 1 VNW pch L=4e-08 W=1.55e-07 
M4 7 1 VDD VNW pch L=4e-08 W=4e-07 
M5 Y A 7 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2XB_X1P4M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y A VSS VPW nch L=4e-08 W=2.3e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.3e-07 
M3 VDD BN 1 VNW pch L=4e-08 W=1.55e-07 
M4 7 1 VDD VNW pch L=4e-08 W=2.85e-07 
M5 Y A 7 VNW pch L=4e-08 W=2.85e-07 
M6 8 A Y VNW pch L=4e-08 W=2.85e-07 
M7 VDD 1 8 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR2XB_X2M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=1.45e-07 
M1 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=3.2e-07 
M3 VDD BN 1 VNW pch L=4e-08 W=1.9e-07 
M4 7 1 VDD VNW pch L=4e-08 W=4e-07 
M5 Y A 7 VNW pch L=4e-08 W=4e-07 
M6 8 A Y VNW pch L=4e-08 W=4e-07 
M7 VDD 1 8 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2XB_X3M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=2.15e-07 
M1 Y A VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS 1 Y VPW nch L=4e-08 W=2.4e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.4e-07 
M4 VSS A Y VPW nch L=4e-08 W=2.4e-07 
M5 VDD BN 1 VNW pch L=4e-08 W=2.75e-07 
M6 7 1 VDD VNW pch L=4e-08 W=4e-07 
M7 Y A 7 VNW pch L=4e-08 W=4e-07 
M8 8 A Y VNW pch L=4e-08 W=4e-07 
M9 VDD 1 8 VNW pch L=4e-08 W=4e-07 
M10 9 1 VDD VNW pch L=4e-08 W=4e-07 
M11 Y A 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2XB_X4M_A9TR Y VDD VNW VPW VSS A BN
M0 VSS BN 1 VPW nch L=4e-08 W=2.8e-07 
M1 Y 1 VSS VPW nch L=4e-08 W=3.2e-07 
M2 VSS A Y VPW nch L=4e-08 W=3.2e-07 
M3 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=3.2e-07 
M5 VDD BN 1 VNW pch L=4e-08 W=3.6e-07 
M6 7 1 VDD VNW pch L=4e-08 W=4e-07 
M7 Y A 7 VNW pch L=4e-08 W=4e-07 
M8 8 A Y VNW pch L=4e-08 W=4e-07 
M9 VDD 1 8 VNW pch L=4e-08 W=4e-07 
M10 9 1 VDD VNW pch L=4e-08 W=4e-07 
M11 Y A 9 VNW pch L=4e-08 W=4e-07 
M12 10 A Y VNW pch L=4e-08 W=4e-07 
M13 VDD 1 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2XB_X6M_A9TR Y VDD VNW VPW VSS A BN
M0 3 BN VSS VPW nch L=4e-08 W=2.1e-07 
M1 VSS BN 3 VPW nch L=4e-08 W=2.1e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS A Y VPW nch L=4e-08 W=3.2e-07 
M6 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M8 3 BN VDD VNW pch L=4e-08 W=2.75e-07 
M9 VDD BN 3 VNW pch L=4e-08 W=2.75e-07 
M10 7 3 VDD VNW pch L=4e-08 W=4e-07 
M11 Y A 7 VNW pch L=4e-08 W=4e-07 
M12 8 A Y VNW pch L=4e-08 W=4e-07 
M13 VDD 3 8 VNW pch L=4e-08 W=4e-07 
M14 9 3 VDD VNW pch L=4e-08 W=4e-07 
M15 Y A 9 VNW pch L=4e-08 W=4e-07 
M16 10 A Y VNW pch L=4e-08 W=4e-07 
M17 VDD 3 10 VNW pch L=4e-08 W=4e-07 
M18 11 3 VDD VNW pch L=4e-08 W=4e-07 
M19 Y A 11 VNW pch L=4e-08 W=4e-07 
M20 12 A Y VNW pch L=4e-08 W=4e-07 
M21 VDD 3 12 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2XB_X8M_A9TR Y VDD VNW VPW VSS A BN
M0 3 BN VSS VPW nch L=4e-08 W=2.8e-07 
M1 VSS BN 3 VPW nch L=4e-08 W=2.8e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.2e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M7 VSS A Y VPW nch L=4e-08 W=3.2e-07 
M8 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M9 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M10 3 BN VDD VNW pch L=4e-08 W=3.6e-07 
M11 VDD BN 3 VNW pch L=4e-08 W=3.6e-07 
M12 7 3 VDD VNW pch L=4e-08 W=4e-07 
M13 Y A 7 VNW pch L=4e-08 W=4e-07 
M14 8 A Y VNW pch L=4e-08 W=4e-07 
M15 VDD 3 8 VNW pch L=4e-08 W=4e-07 
M16 9 3 VDD VNW pch L=4e-08 W=4e-07 
M17 Y A 9 VNW pch L=4e-08 W=4e-07 
M18 10 A Y VNW pch L=4e-08 W=4e-07 
M19 VDD 3 10 VNW pch L=4e-08 W=4e-07 
M20 11 3 VDD VNW pch L=4e-08 W=4e-07 
M21 Y A 11 VNW pch L=4e-08 W=4e-07 
M22 12 A Y VNW pch L=4e-08 W=4e-07 
M23 VDD 3 12 VNW pch L=4e-08 W=4e-07 
M24 13 3 VDD VNW pch L=4e-08 W=4e-07 
M25 Y A 13 VNW pch L=4e-08 W=4e-07 
M26 14 A Y VNW pch L=4e-08 W=4e-07 
M27 VDD 3 14 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X0P5A_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=1.45e-07 
M1 VSS A Y VPW nch L=4e-08 W=1.45e-07 
M2 6 B VDD VNW pch L=4e-08 W=2e-07 
M3 Y A 6 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT NOR2_X0P5B_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS A Y VPW nch L=4e-08 W=1.2e-07 
M2 6 B VDD VNW pch L=4e-08 W=3.6e-07 
M3 Y A 6 VNW pch L=4e-08 W=3.6e-07 
.ENDS


.SUBCKT NOR2_X0P5M_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS A Y VPW nch L=4e-08 W=1.2e-07 
M2 6 B VDD VNW pch L=4e-08 W=2e-07 
M3 Y A 6 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT NOR2_X0P7A_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=2.05e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.05e-07 
M2 6 B VDD VNW pch L=4e-08 W=2.85e-07 
M3 Y A 6 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR2_X0P7B_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=1.25e-07 
M1 VSS A Y VPW nch L=4e-08 W=1.25e-07 
M2 6 B VDD VNW pch L=4e-08 W=3.75e-07 
M3 Y A 6 VNW pch L=4e-08 W=3.75e-07 
.ENDS


.SUBCKT NOR2_X0P7M_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS A Y VPW nch L=4e-08 W=1.2e-07 
M2 6 B VDD VNW pch L=4e-08 W=2.95e-07 
M3 Y A 6 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT NOR2_X1A_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M2 6 B VDD VNW pch L=4e-08 W=4e-07 
M3 Y A 6 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X1B_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=1.35e-07 
M1 VSS A Y VPW nch L=4e-08 W=1.35e-07 
M2 6 B VDD VNW pch L=4e-08 W=4e-07 
M3 Y A 6 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X1M_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS A Y VPW nch L=4e-08 W=1.6e-07 
M2 6 B VDD VNW pch L=4e-08 W=4e-07 
M3 Y A 6 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X1P4A_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=2.05e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.05e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.05e-07 
M3 VSS B Y VPW nch L=4e-08 W=2.05e-07 
M4 6 B VDD VNW pch L=4e-08 W=2.85e-07 
M5 Y A 6 VNW pch L=4e-08 W=2.85e-07 
M6 7 A Y VNW pch L=4e-08 W=2.85e-07 
M7 VDD B 7 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR2_X1P4B_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=1.9e-07 
M1 VSS B Y VPW nch L=4e-08 W=1.9e-07 
M2 6 B VDD VNW pch L=4e-08 W=2.85e-07 
M3 Y A 6 VNW pch L=4e-08 W=2.85e-07 
M4 7 A Y VNW pch L=4e-08 W=2.85e-07 
M5 VDD B 7 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR2_X1P4M_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=2.3e-07 
M1 VSS B Y VPW nch L=4e-08 W=2.3e-07 
M2 6 B VDD VNW pch L=4e-08 W=2.85e-07 
M3 Y A 6 VNW pch L=4e-08 W=2.85e-07 
M4 7 A Y VNW pch L=4e-08 W=2.85e-07 
M5 VDD B 7 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR2_X2A_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M3 VSS B Y VPW nch L=4e-08 W=2.85e-07 
M4 6 B VDD VNW pch L=4e-08 W=4e-07 
M5 Y A 6 VNW pch L=4e-08 W=4e-07 
M6 7 A Y VNW pch L=4e-08 W=4e-07 
M7 VDD B 7 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X2B_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=2.7e-07 
M1 VSS B Y VPW nch L=4e-08 W=2.7e-07 
M2 6 B VDD VNW pch L=4e-08 W=4e-07 
M3 Y A 6 VNW pch L=4e-08 W=4e-07 
M4 7 A Y VNW pch L=4e-08 W=4e-07 
M5 VDD B 7 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X2M_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M2 6 B VDD VNW pch L=4e-08 W=4e-07 
M3 Y A 6 VNW pch L=4e-08 W=4e-07 
M4 7 A Y VNW pch L=4e-08 W=4e-07 
M5 VDD B 7 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X3A_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M3 VSS B Y VPW nch L=4e-08 W=2.85e-07 
M4 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M5 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M6 6 B VDD VNW pch L=4e-08 W=4e-07 
M7 Y A 6 VNW pch L=4e-08 W=4e-07 
M8 7 A Y VNW pch L=4e-08 W=4e-07 
M9 VDD B 7 VNW pch L=4e-08 W=4e-07 
M10 8 B VDD VNW pch L=4e-08 W=4e-07 
M11 Y A 8 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X3B_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=2e-07 
M1 VSS B Y VPW nch L=4e-08 W=2e-07 
M2 Y B VSS VPW nch L=4e-08 W=2e-07 
M3 VSS A Y VPW nch L=4e-08 W=2e-07 
M4 6 B VDD VNW pch L=4e-08 W=4e-07 
M5 Y A 6 VNW pch L=4e-08 W=4e-07 
M6 7 A Y VNW pch L=4e-08 W=4e-07 
M7 VDD B 7 VNW pch L=4e-08 W=4e-07 
M8 8 B VDD VNW pch L=4e-08 W=4e-07 
M9 Y A 8 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X3M_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=2.4e-07 
M1 VSS B Y VPW nch L=4e-08 W=2.4e-07 
M2 Y B VSS VPW nch L=4e-08 W=2.4e-07 
M3 VSS A Y VPW nch L=4e-08 W=2.4e-07 
M4 6 B VDD VNW pch L=4e-08 W=4e-07 
M5 Y A 6 VNW pch L=4e-08 W=4e-07 
M6 7 A Y VNW pch L=4e-08 W=4e-07 
M7 VDD B 7 VNW pch L=4e-08 W=4e-07 
M8 8 B VDD VNW pch L=4e-08 W=4e-07 
M9 Y A 8 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X4A_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=3.8e-07 
M1 VSS B Y VPW nch L=4e-08 W=3.8e-07 
M2 Y B VSS VPW nch L=4e-08 W=3.8e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.8e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.8e-07 
M5 VSS B Y VPW nch L=4e-08 W=3.8e-07 
M6 6 B VDD VNW pch L=4e-08 W=4e-07 
M7 Y A 6 VNW pch L=4e-08 W=4e-07 
M8 7 A Y VNW pch L=4e-08 W=4e-07 
M9 VDD B 7 VNW pch L=4e-08 W=4e-07 
M10 8 B VDD VNW pch L=4e-08 W=4e-07 
M11 Y A 8 VNW pch L=4e-08 W=4e-07 
M12 9 A Y VNW pch L=4e-08 W=4e-07 
M13 VDD B 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X4B_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=2.7e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.7e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.7e-07 
M3 VSS B Y VPW nch L=4e-08 W=2.7e-07 
M4 6 B VDD VNW pch L=4e-08 W=4e-07 
M5 Y A 6 VNW pch L=4e-08 W=4e-07 
M6 7 A Y VNW pch L=4e-08 W=4e-07 
M7 VDD B 7 VNW pch L=4e-08 W=4e-07 
M8 8 B VDD VNW pch L=4e-08 W=4e-07 
M9 Y A 8 VNW pch L=4e-08 W=4e-07 
M10 9 A Y VNW pch L=4e-08 W=4e-07 
M11 VDD B 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X4M_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.2e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M4 6 B VDD VNW pch L=4e-08 W=4e-07 
M5 Y A 6 VNW pch L=4e-08 W=4e-07 
M6 7 A Y VNW pch L=4e-08 W=4e-07 
M7 VDD B 7 VNW pch L=4e-08 W=4e-07 
M8 8 B VDD VNW pch L=4e-08 W=4e-07 
M9 Y A 8 VNW pch L=4e-08 W=4e-07 
M10 9 A Y VNW pch L=4e-08 W=4e-07 
M11 VDD B 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X6A_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M3 VSS B Y VPW nch L=4e-08 W=2.85e-07 
M4 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M5 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M6 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M7 VSS B Y VPW nch L=4e-08 W=2.85e-07 
M8 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M9 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M10 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M11 VSS B Y VPW nch L=4e-08 W=2.85e-07 
M12 6 B VDD VNW pch L=4e-08 W=4e-07 
M13 Y A 6 VNW pch L=4e-08 W=4e-07 
M14 7 A Y VNW pch L=4e-08 W=4e-07 
M15 VDD B 7 VNW pch L=4e-08 W=4e-07 
M16 8 B VDD VNW pch L=4e-08 W=4e-07 
M17 Y A 8 VNW pch L=4e-08 W=4e-07 
M18 9 A Y VNW pch L=4e-08 W=4e-07 
M19 VDD B 9 VNW pch L=4e-08 W=4e-07 
M20 10 B VDD VNW pch L=4e-08 W=4e-07 
M21 Y A 10 VNW pch L=4e-08 W=4e-07 
M22 11 A Y VNW pch L=4e-08 W=4e-07 
M23 VDD B 11 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X6B_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=2.65e-07 
M1 VSS B Y VPW nch L=4e-08 W=2.65e-07 
M2 Y B VSS VPW nch L=4e-08 W=2.65e-07 
M3 VSS A Y VPW nch L=4e-08 W=2.65e-07 
M4 Y A VSS VPW nch L=4e-08 W=2.65e-07 
M5 VSS B Y VPW nch L=4e-08 W=2.65e-07 
M6 6 B VDD VNW pch L=4e-08 W=4e-07 
M7 Y A 6 VNW pch L=4e-08 W=4e-07 
M8 7 A Y VNW pch L=4e-08 W=4e-07 
M9 VDD B 7 VNW pch L=4e-08 W=4e-07 
M10 8 B VDD VNW pch L=4e-08 W=4e-07 
M11 Y A 8 VNW pch L=4e-08 W=4e-07 
M12 9 A Y VNW pch L=4e-08 W=4e-07 
M13 VDD B 9 VNW pch L=4e-08 W=4e-07 
M14 10 B VDD VNW pch L=4e-08 W=4e-07 
M15 Y A 10 VNW pch L=4e-08 W=4e-07 
M16 11 A Y VNW pch L=4e-08 W=4e-07 
M17 VDD B 11 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X6M_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M2 Y B VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.2e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M6 6 B VDD VNW pch L=4e-08 W=4e-07 
M7 Y A 6 VNW pch L=4e-08 W=4e-07 
M8 7 A Y VNW pch L=4e-08 W=4e-07 
M9 VDD B 7 VNW pch L=4e-08 W=4e-07 
M10 8 B VDD VNW pch L=4e-08 W=4e-07 
M11 Y A 8 VNW pch L=4e-08 W=4e-07 
M12 9 A Y VNW pch L=4e-08 W=4e-07 
M13 VDD B 9 VNW pch L=4e-08 W=4e-07 
M14 10 B VDD VNW pch L=4e-08 W=4e-07 
M15 Y A 10 VNW pch L=4e-08 W=4e-07 
M16 11 A Y VNW pch L=4e-08 W=4e-07 
M17 VDD B 11 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X8A_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M3 VSS B Y VPW nch L=4e-08 W=2.85e-07 
M4 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M5 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M6 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M7 VSS B Y VPW nch L=4e-08 W=2.85e-07 
M8 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M9 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M10 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M11 VSS B Y VPW nch L=4e-08 W=2.85e-07 
M12 Y B VSS VPW nch L=4e-08 W=2.85e-07 
M13 VSS A Y VPW nch L=4e-08 W=2.85e-07 
M14 Y A VSS VPW nch L=4e-08 W=2.85e-07 
M15 VSS B Y VPW nch L=4e-08 W=2.85e-07 
M16 6 B VDD VNW pch L=4e-08 W=4e-07 
M17 Y A 6 VNW pch L=4e-08 W=4e-07 
M18 7 A Y VNW pch L=4e-08 W=4e-07 
M19 VDD B 7 VNW pch L=4e-08 W=4e-07 
M20 8 B VDD VNW pch L=4e-08 W=4e-07 
M21 Y A 8 VNW pch L=4e-08 W=4e-07 
M22 9 A Y VNW pch L=4e-08 W=4e-07 
M23 VDD B 9 VNW pch L=4e-08 W=4e-07 
M24 10 B VDD VNW pch L=4e-08 W=4e-07 
M25 Y A 10 VNW pch L=4e-08 W=4e-07 
M26 11 A Y VNW pch L=4e-08 W=4e-07 
M27 VDD B 11 VNW pch L=4e-08 W=4e-07 
M28 12 B VDD VNW pch L=4e-08 W=4e-07 
M29 Y A 12 VNW pch L=4e-08 W=4e-07 
M30 13 A Y VNW pch L=4e-08 W=4e-07 
M31 VDD B 13 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X8B_A9TR Y VDD VNW VPW VSS A B
M0 Y A VSS VPW nch L=4e-08 W=3.6e-07 
M1 VSS B Y VPW nch L=4e-08 W=3.6e-07 
M2 Y B VSS VPW nch L=4e-08 W=3.6e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.6e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.6e-07 
M5 VSS B Y VPW nch L=4e-08 W=3.6e-07 
M6 6 B VDD VNW pch L=4e-08 W=4e-07 
M7 Y A 6 VNW pch L=4e-08 W=4e-07 
M8 7 A Y VNW pch L=4e-08 W=4e-07 
M9 VDD B 7 VNW pch L=4e-08 W=4e-07 
M10 8 B VDD VNW pch L=4e-08 W=4e-07 
M11 Y A 8 VNW pch L=4e-08 W=4e-07 
M12 9 A Y VNW pch L=4e-08 W=4e-07 
M13 VDD B 9 VNW pch L=4e-08 W=4e-07 
M14 10 B VDD VNW pch L=4e-08 W=4e-07 
M15 Y A 10 VNW pch L=4e-08 W=4e-07 
M16 11 A Y VNW pch L=4e-08 W=4e-07 
M17 VDD B 11 VNW pch L=4e-08 W=4e-07 
M18 12 B VDD VNW pch L=4e-08 W=4e-07 
M19 Y A 12 VNW pch L=4e-08 W=4e-07 
M20 13 A Y VNW pch L=4e-08 W=4e-07 
M21 VDD B 13 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR2_X8M_A9TR Y VDD VNW VPW VSS A B
M0 Y B VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS A Y VPW nch L=4e-08 W=3.2e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M4 Y B VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS A Y VPW nch L=4e-08 W=3.2e-07 
M6 Y A VSS VPW nch L=4e-08 W=3.2e-07 
M7 VSS B Y VPW nch L=4e-08 W=3.2e-07 
M8 6 B VDD VNW pch L=4e-08 W=4e-07 
M9 Y A 6 VNW pch L=4e-08 W=4e-07 
M10 7 A Y VNW pch L=4e-08 W=4e-07 
M11 VDD B 7 VNW pch L=4e-08 W=4e-07 
M12 8 B VDD VNW pch L=4e-08 W=4e-07 
M13 Y A 8 VNW pch L=4e-08 W=4e-07 
M14 9 A Y VNW pch L=4e-08 W=4e-07 
M15 VDD B 9 VNW pch L=4e-08 W=4e-07 
M16 10 B VDD VNW pch L=4e-08 W=4e-07 
M17 Y A 10 VNW pch L=4e-08 W=4e-07 
M18 11 A Y VNW pch L=4e-08 W=4e-07 
M19 VDD B 11 VNW pch L=4e-08 W=4e-07 
M20 12 B VDD VNW pch L=4e-08 W=4e-07 
M21 Y A 12 VNW pch L=4e-08 W=4e-07 
M22 13 A Y VNW pch L=4e-08 W=4e-07 
M23 VDD B 13 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3BB_X0P5M_A9TR Y VDD VNW VPW VSS AN BN C
M0 9 AN 1 VPW nch L=4e-08 W=1.3e-07 
M1 VSS BN 9 VPW nch L=4e-08 W=1.3e-07 
M2 Y C VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=1.2e-07 
M4 1 AN VDD VNW pch L=4e-08 W=1.2e-07 
M5 VDD BN 1 VNW pch L=4e-08 W=1.2e-07 
M6 8 C VDD VNW pch L=4e-08 W=2e-07 
M7 Y 1 8 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT NOR3BB_X0P7M_A9TR Y VDD VNW VPW VSS AN BN C
M0 9 AN 1 VPW nch L=4e-08 W=1.45e-07 
M1 VSS BN 9 VPW nch L=4e-08 W=1.45e-07 
M2 Y C VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=1.2e-07 
M4 1 AN VDD VNW pch L=4e-08 W=1.25e-07 
M5 VDD BN 1 VNW pch L=4e-08 W=1.25e-07 
M6 8 C VDD VNW pch L=4e-08 W=2.95e-07 
M7 Y 1 8 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT NOR3BB_X1M_A9TR Y VDD VNW VPW VSS AN BN C
M0 9 AN 1 VPW nch L=4e-08 W=1.7e-07 
M1 VSS BN 9 VPW nch L=4e-08 W=1.7e-07 
M2 Y C VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M4 1 AN VDD VNW pch L=4e-08 W=1.5e-07 
M5 VDD BN 1 VNW pch L=4e-08 W=1.5e-07 
M6 8 C VDD VNW pch L=4e-08 W=3.9e-07 
M7 Y 1 8 VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT NOR3BB_X1P4M_A9TR Y VDD VNW VPW VSS AN BN C
M0 10 AN 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS BN 10 VPW nch L=4e-08 W=1.2e-07 
M2 Y C VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=1.2e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M5 VSS C Y VPW nch L=4e-08 W=1.2e-07 
M6 1 AN VDD VNW pch L=4e-08 W=1.55e-07 
M7 VDD BN 1 VNW pch L=4e-08 W=1.55e-07 
M8 8 C VDD VNW pch L=4e-08 W=2.85e-07 
M9 Y 1 8 VNW pch L=4e-08 W=2.85e-07 
M10 9 1 Y VNW pch L=4e-08 W=2.85e-07 
M11 VDD C 9 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR3BB_X2M_A9TR Y VDD VNW VPW VSS AN BN C
M0 10 AN 1 VPW nch L=4e-08 W=2.9e-07 
M1 VSS BN 10 VPW nch L=4e-08 W=2.9e-07 
M2 Y C VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS C Y VPW nch L=4e-08 W=1.6e-07 
M6 1 AN VDD VNW pch L=4e-08 W=2.5e-07 
M7 VDD BN 1 VNW pch L=4e-08 W=2.5e-07 
M8 8 C VDD VNW pch L=4e-08 W=4e-07 
M9 Y 1 8 VNW pch L=4e-08 W=4e-07 
M10 9 1 Y VNW pch L=4e-08 W=4e-07 
M11 VDD C 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3BB_X3M_A9TR Y VDD VNW VPW VSS AN BN C
M0 11 AN 1 VPW nch L=4e-08 W=4e-07 
M1 VSS BN 11 VPW nch L=4e-08 W=4e-07 
M2 Y C VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS C Y VPW nch L=4e-08 W=1.6e-07 
M6 Y C VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M8 1 AN VDD VNW pch L=4e-08 W=3.5e-07 
M9 VDD BN 1 VNW pch L=4e-08 W=3.5e-07 
M10 8 C VDD VNW pch L=4e-08 W=4e-07 
M11 Y 1 8 VNW pch L=4e-08 W=4e-07 
M12 9 1 Y VNW pch L=4e-08 W=4e-07 
M13 VDD C 9 VNW pch L=4e-08 W=4e-07 
M14 10 C VDD VNW pch L=4e-08 W=4e-07 
M15 Y 1 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3BB_X4M_A9TR Y VDD VNW VPW VSS AN BN C
M0 12 BN VSS VPW nch L=4e-08 W=2.9e-07 
M1 3 AN 12 VPW nch L=4e-08 W=2.9e-07 
M2 13 AN 3 VPW nch L=4e-08 W=2.9e-07 
M3 VSS BN 13 VPW nch L=4e-08 W=2.9e-07 
M4 Y C VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M7 VSS C Y VPW nch L=4e-08 W=3.2e-07 
M8 3 BN VDD VNW pch L=4e-08 W=2.5e-07 
M9 VDD AN 3 VNW pch L=4e-08 W=2.5e-07 
M10 3 AN VDD VNW pch L=4e-08 W=2.5e-07 
M11 VDD BN 3 VNW pch L=4e-08 W=2.5e-07 
M12 8 C VDD VNW pch L=4e-08 W=4e-07 
M13 Y 3 8 VNW pch L=4e-08 W=4e-07 
M14 9 3 Y VNW pch L=4e-08 W=4e-07 
M15 VDD C 9 VNW pch L=4e-08 W=4e-07 
M16 10 C VDD VNW pch L=4e-08 W=4e-07 
M17 Y 3 10 VNW pch L=4e-08 W=4e-07 
M18 11 3 Y VNW pch L=4e-08 W=4e-07 
M19 VDD C 11 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3BB_X6M_A9TR Y VDD VNW VPW VSS AN BN C
M0 14 BN VSS VPW nch L=4e-08 W=4e-07 
M1 3 AN 14 VPW nch L=4e-08 W=4e-07 
M2 15 AN 3 VPW nch L=4e-08 W=4e-07 
M3 VSS BN 15 VPW nch L=4e-08 W=4e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS C Y VPW nch L=4e-08 W=3.2e-07 
M6 Y C VSS VPW nch L=4e-08 W=3.2e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=3.2e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=3.2e-07 
M9 VSS C Y VPW nch L=4e-08 W=3.2e-07 
M10 3 BN VDD VNW pch L=4e-08 W=3.45e-07 
M11 VDD AN 3 VNW pch L=4e-08 W=3.45e-07 
M12 3 AN VDD VNW pch L=4e-08 W=3.45e-07 
M13 VDD BN 3 VNW pch L=4e-08 W=3.45e-07 
M14 8 C VDD VNW pch L=4e-08 W=4e-07 
M15 Y 3 8 VNW pch L=4e-08 W=4e-07 
M16 9 3 Y VNW pch L=4e-08 W=4e-07 
M17 VDD C 9 VNW pch L=4e-08 W=4e-07 
M18 10 C VDD VNW pch L=4e-08 W=4e-07 
M19 Y 3 10 VNW pch L=4e-08 W=4e-07 
M20 11 3 Y VNW pch L=4e-08 W=4e-07 
M21 VDD C 11 VNW pch L=4e-08 W=4e-07 
M22 12 C VDD VNW pch L=4e-08 W=4e-07 
M23 Y 3 12 VNW pch L=4e-08 W=4e-07 
M24 13 3 Y VNW pch L=4e-08 W=4e-07 
M25 VDD C 13 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3BB_X8M_A9TR Y VDD VNW VPW VSS AN BN C
M0 16 AN 1 VPW nch L=4e-08 W=3.8e-07 
M1 VSS BN 16 VPW nch L=4e-08 W=3.8e-07 
M2 17 BN VSS VPW nch L=4e-08 W=3.8e-07 
M3 1 AN 17 VPW nch L=4e-08 W=3.8e-07 
M4 18 AN 1 VPW nch L=4e-08 W=3.8e-07 
M5 VSS BN 18 VPW nch L=4e-08 W=3.8e-07 
M6 Y C VSS VPW nch L=4e-08 W=3.2e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.2e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.2e-07 
M9 VSS C Y VPW nch L=4e-08 W=3.2e-07 
M10 Y C VSS VPW nch L=4e-08 W=3.2e-07 
M11 VSS 1 Y VPW nch L=4e-08 W=3.2e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=3.2e-07 
M13 VSS C Y VPW nch L=4e-08 W=3.2e-07 
M14 1 AN VDD VNW pch L=4e-08 W=3.3e-07 
M15 VDD BN 1 VNW pch L=4e-08 W=3.3e-07 
M16 1 BN VDD VNW pch L=4e-08 W=3.3e-07 
M17 VDD AN 1 VNW pch L=4e-08 W=3.3e-07 
M18 1 AN VDD VNW pch L=4e-08 W=3.3e-07 
M19 VDD BN 1 VNW pch L=4e-08 W=3.3e-07 
M20 8 C VDD VNW pch L=4e-08 W=4e-07 
M21 Y 1 8 VNW pch L=4e-08 W=4e-07 
M22 9 1 Y VNW pch L=4e-08 W=4e-07 
M23 VDD C 9 VNW pch L=4e-08 W=4e-07 
M24 10 C VDD VNW pch L=4e-08 W=4e-07 
M25 Y 1 10 VNW pch L=4e-08 W=4e-07 
M26 11 1 Y VNW pch L=4e-08 W=4e-07 
M27 VDD C 11 VNW pch L=4e-08 W=4e-07 
M28 12 C VDD VNW pch L=4e-08 W=4e-07 
M29 Y 1 12 VNW pch L=4e-08 W=4e-07 
M30 13 1 Y VNW pch L=4e-08 W=4e-07 
M31 VDD C 13 VNW pch L=4e-08 W=4e-07 
M32 14 C VDD VNW pch L=4e-08 W=4e-07 
M33 Y 1 14 VNW pch L=4e-08 W=4e-07 
M34 15 1 Y VNW pch L=4e-08 W=4e-07 
M35 VDD C 15 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3_X0P5A_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B Y VPW nch L=4e-08 W=1.2e-07 
M2 Y A VSS VPW nch L=4e-08 W=1.2e-07 
M3 7 C VDD VNW pch L=4e-08 W=2.2e-07 
M4 8 B 7 VNW pch L=4e-08 W=2.2e-07 
M5 Y A 8 VNW pch L=4e-08 W=2.2e-07 
.ENDS


.SUBCKT NOR3_X0P5M_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B Y VPW nch L=4e-08 W=1.2e-07 
M2 Y A VSS VPW nch L=4e-08 W=1.2e-07 
M3 7 C VDD VNW pch L=4e-08 W=2e-07 
M4 8 B 7 VNW pch L=4e-08 W=2e-07 
M5 Y A 8 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT NOR3_X0P7A_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=1.55e-07 
M1 VSS B Y VPW nch L=4e-08 W=1.55e-07 
M2 Y A VSS VPW nch L=4e-08 W=1.55e-07 
M3 7 C VDD VNW pch L=4e-08 W=2.85e-07 
M4 8 B 7 VNW pch L=4e-08 W=2.85e-07 
M5 Y A 8 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR3_X0P7M_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B Y VPW nch L=4e-08 W=1.2e-07 
M2 Y A VSS VPW nch L=4e-08 W=1.2e-07 
M3 7 C VDD VNW pch L=4e-08 W=2.85e-07 
M4 8 B 7 VNW pch L=4e-08 W=2.85e-07 
M5 Y A 8 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR3_X1A_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS B Y VPW nch L=4e-08 W=2.2e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.2e-07 
M3 7 C VDD VNW pch L=4e-08 W=4e-07 
M4 8 B 7 VNW pch L=4e-08 W=4e-07 
M5 Y A 8 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3_X1M_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B Y VPW nch L=4e-08 W=1.2e-07 
M2 Y A VSS VPW nch L=4e-08 W=1.2e-07 
M3 7 C VDD VNW pch L=4e-08 W=4e-07 
M4 8 B 7 VNW pch L=4e-08 W=4e-07 
M5 Y A 8 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3_X1P4A_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS B Y VPW nch L=4e-08 W=3.1e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.1e-07 
M3 VDD C 1 VNW pch L=4e-08 W=2.85e-07 
M4 1 C VDD VNW pch L=4e-08 W=2.85e-07 
M5 8 B 1 VNW pch L=4e-08 W=2.85e-07 
M6 Y A 8 VNW pch L=4e-08 W=2.85e-07 
M7 9 A Y VNW pch L=4e-08 W=2.85e-07 
M8 1 B 9 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR3_X1P4M_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=1.5e-07 
M1 VSS B Y VPW nch L=4e-08 W=1.5e-07 
M2 Y A VSS VPW nch L=4e-08 W=1.5e-07 
M3 VDD C 1 VNW pch L=4e-08 W=2.85e-07 
M4 1 C VDD VNW pch L=4e-08 W=2.85e-07 
M5 8 B 1 VNW pch L=4e-08 W=2.85e-07 
M6 Y A 8 VNW pch L=4e-08 W=2.85e-07 
M7 9 A Y VNW pch L=4e-08 W=2.85e-07 
M8 1 B 9 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR3_X2A_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS C Y VPW nch L=4e-08 W=2.2e-07 
M2 Y B VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS A Y VPW nch L=4e-08 W=2.2e-07 
M4 Y A VSS VPW nch L=4e-08 W=2.2e-07 
M5 VSS B Y VPW nch L=4e-08 W=2.2e-07 
M6 VDD C 2 VNW pch L=4e-08 W=4e-07 
M7 2 C VDD VNW pch L=4e-08 W=4e-07 
M8 8 B 2 VNW pch L=4e-08 W=4e-07 
M9 Y A 8 VNW pch L=4e-08 W=4e-07 
M10 9 A Y VNW pch L=4e-08 W=4e-07 
M11 2 B 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3_X2M_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS B Y VPW nch L=4e-08 W=2.2e-07 
M2 Y A VSS VPW nch L=4e-08 W=2.2e-07 
M3 VDD C 1 VNW pch L=4e-08 W=4e-07 
M4 1 C VDD VNW pch L=4e-08 W=4e-07 
M5 8 B 1 VNW pch L=4e-08 W=4e-07 
M6 Y A 8 VNW pch L=4e-08 W=4e-07 
M7 9 A Y VNW pch L=4e-08 W=4e-07 
M8 1 B 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3_X3A_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=3.3e-07 
M1 VSS C Y VPW nch L=4e-08 W=3.3e-07 
M2 Y B VSS VPW nch L=4e-08 W=3.3e-07 
M3 VSS A Y VPW nch L=4e-08 W=3.3e-07 
M4 Y A VSS VPW nch L=4e-08 W=3.3e-07 
M5 VSS B Y VPW nch L=4e-08 W=3.3e-07 
M6 3 C VDD VNW pch L=4e-08 W=4e-07 
M7 VDD C 3 VNW pch L=4e-08 W=4e-07 
M8 3 C VDD VNW pch L=4e-08 W=4e-07 
M9 8 B 3 VNW pch L=4e-08 W=4e-07 
M10 Y A 8 VNW pch L=4e-08 W=4e-07 
M11 9 A Y VNW pch L=4e-08 W=4e-07 
M12 3 B 9 VNW pch L=4e-08 W=4e-07 
M13 10 B 3 VNW pch L=4e-08 W=4e-07 
M14 Y A 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3_X3M_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=3.3e-07 
M1 VSS B Y VPW nch L=4e-08 W=3.3e-07 
M2 Y A VSS VPW nch L=4e-08 W=3.3e-07 
M3 2 C VDD VNW pch L=4e-08 W=4e-07 
M4 VDD C 2 VNW pch L=4e-08 W=4e-07 
M5 2 C VDD VNW pch L=4e-08 W=4e-07 
M6 8 B 2 VNW pch L=4e-08 W=4e-07 
M7 Y A 8 VNW pch L=4e-08 W=4e-07 
M8 9 A Y VNW pch L=4e-08 W=4e-07 
M9 2 B 9 VNW pch L=4e-08 W=4e-07 
M10 10 B 2 VNW pch L=4e-08 W=4e-07 
M11 Y A 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3_X4A_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS C Y VPW nch L=4e-08 W=2.2e-07 
M2 Y C VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS C Y VPW nch L=4e-08 W=2.2e-07 
M4 Y B VSS VPW nch L=4e-08 W=2.2e-07 
M5 VSS A Y VPW nch L=4e-08 W=2.2e-07 
M6 Y A VSS VPW nch L=4e-08 W=2.2e-07 
M7 VSS B Y VPW nch L=4e-08 W=2.2e-07 
M8 Y B VSS VPW nch L=4e-08 W=2.2e-07 
M9 VSS A Y VPW nch L=4e-08 W=2.2e-07 
M10 Y A VSS VPW nch L=4e-08 W=2.2e-07 
M11 VSS B Y VPW nch L=4e-08 W=2.2e-07 
M12 VDD C 2 VNW pch L=4e-08 W=4e-07 
M13 2 C VDD VNW pch L=4e-08 W=4e-07 
M14 VDD C 2 VNW pch L=4e-08 W=4e-07 
M15 2 C VDD VNW pch L=4e-08 W=4e-07 
M16 8 B 2 VNW pch L=4e-08 W=4e-07 
M17 Y A 8 VNW pch L=4e-08 W=4e-07 
M18 9 A Y VNW pch L=4e-08 W=4e-07 
M19 2 B 9 VNW pch L=4e-08 W=4e-07 
M20 10 B 2 VNW pch L=4e-08 W=4e-07 
M21 Y A 10 VNW pch L=4e-08 W=4e-07 
M22 11 A Y VNW pch L=4e-08 W=4e-07 
M23 2 B 11 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR3_X4M_A9TR Y VDD VNW VPW VSS A B C
M0 Y C VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS C Y VPW nch L=4e-08 W=2.2e-07 
M2 Y B VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS A Y VPW nch L=4e-08 W=2.2e-07 
M4 Y A VSS VPW nch L=4e-08 W=2.2e-07 
M5 VSS B Y VPW nch L=4e-08 W=2.2e-07 
M6 VDD C 1 VNW pch L=4e-08 W=4e-07 
M7 1 C VDD VNW pch L=4e-08 W=4e-07 
M8 VDD C 1 VNW pch L=4e-08 W=4e-07 
M9 1 C VDD VNW pch L=4e-08 W=4e-07 
M10 8 B 1 VNW pch L=4e-08 W=4e-07 
M11 Y A 8 VNW pch L=4e-08 W=4e-07 
M12 9 A Y VNW pch L=4e-08 W=4e-07 
M13 1 B 9 VNW pch L=4e-08 W=4e-07 
M14 10 B 1 VNW pch L=4e-08 W=4e-07 
M15 Y A 10 VNW pch L=4e-08 W=4e-07 
M16 11 A Y VNW pch L=4e-08 W=4e-07 
M17 1 B 11 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR4BB_X0P5M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 11 AN 1 VPW nch L=4e-08 W=1.3e-07 
M1 VSS BN 11 VPW nch L=4e-08 W=1.3e-07 
M2 Y D VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS C Y VPW nch L=4e-08 W=1.2e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M5 1 AN VDD VNW pch L=4e-08 W=1.2e-07 
M6 VDD BN 1 VNW pch L=4e-08 W=1.2e-07 
M7 9 D VDD VNW pch L=4e-08 W=2e-07 
M8 10 C 9 VNW pch L=4e-08 W=2e-07 
M9 Y 1 10 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT NOR4BB_X0P7M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 11 AN 1 VPW nch L=4e-08 W=1.45e-07 
M1 VSS BN 11 VPW nch L=4e-08 W=1.45e-07 
M2 Y D VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS C Y VPW nch L=4e-08 W=1.2e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M5 1 AN VDD VNW pch L=4e-08 W=1.25e-07 
M6 VDD BN 1 VNW pch L=4e-08 W=1.25e-07 
M7 9 D VDD VNW pch L=4e-08 W=2.85e-07 
M8 10 C 9 VNW pch L=4e-08 W=2.85e-07 
M9 Y 1 10 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR4BB_X1M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 11 AN 1 VPW nch L=4e-08 W=1.65e-07 
M1 VSS BN 11 VPW nch L=4e-08 W=1.65e-07 
M2 Y D VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS C Y VPW nch L=4e-08 W=1.2e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M5 1 AN VDD VNW pch L=4e-08 W=1.4e-07 
M6 VDD BN 1 VNW pch L=4e-08 W=1.4e-07 
M7 9 D VDD VNW pch L=4e-08 W=4e-07 
M8 10 C 9 VNW pch L=4e-08 W=4e-07 
M9 Y 1 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR4BB_X1P4M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 13 AN 1 VPW nch L=4e-08 W=2.1e-07 
M1 VSS BN 13 VPW nch L=4e-08 W=2.1e-07 
M2 Y D VSS VPW nch L=4e-08 W=1.5e-07 
M3 VSS C Y VPW nch L=4e-08 W=1.5e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.5e-07 
M5 1 AN VDD VNW pch L=4e-08 W=1.8e-07 
M6 VDD BN 1 VNW pch L=4e-08 W=1.8e-07 
M7 9 D VDD VNW pch L=4e-08 W=2.85e-07 
M8 10 C 9 VNW pch L=4e-08 W=2.85e-07 
M9 Y 1 10 VNW pch L=4e-08 W=2.85e-07 
M10 11 1 Y VNW pch L=4e-08 W=2.85e-07 
M11 12 C 11 VNW pch L=4e-08 W=2.85e-07 
M12 VDD D 12 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT NOR4BB_X2M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 13 AN 1 VPW nch L=4e-08 W=2.7e-07 
M1 VSS BN 13 VPW nch L=4e-08 W=2.7e-07 
M2 Y D VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS C Y VPW nch L=4e-08 W=1.2e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M5 VSS 1 Y VPW nch L=4e-08 W=1.2e-07 
M6 Y C VSS VPW nch L=4e-08 W=1.2e-07 
M7 VSS D Y VPW nch L=4e-08 W=1.2e-07 
M8 1 AN VDD VNW pch L=4e-08 W=2.3e-07 
M9 VDD BN 1 VNW pch L=4e-08 W=2.3e-07 
M10 9 D VDD VNW pch L=4e-08 W=4e-07 
M11 10 C 9 VNW pch L=4e-08 W=4e-07 
M12 Y 1 10 VNW pch L=4e-08 W=4e-07 
M13 11 1 Y VNW pch L=4e-08 W=4e-07 
M14 12 C 11 VNW pch L=4e-08 W=4e-07 
M15 VDD D 12 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR4BB_X3M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 13 AN 1 VPW nch L=4e-08 W=3.8e-07 
M1 VSS BN 13 VPW nch L=4e-08 W=3.8e-07 
M2 Y D VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS D Y VPW nch L=4e-08 W=1.2e-07 
M4 Y D VSS VPW nch L=4e-08 W=1.2e-07 
M5 VSS C Y VPW nch L=4e-08 W=1.2e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=1.2e-07 
M8 Y C VSS VPW nch L=4e-08 W=1.2e-07 
M9 VSS C Y VPW nch L=4e-08 W=1.2e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=1.2e-07 
M11 1 AN VDD VNW pch L=4e-08 W=3.3e-07 
M12 VDD BN 1 VNW pch L=4e-08 W=3.3e-07 
M13 5 D VDD VNW pch L=4e-08 W=4e-07 
M14 VDD D 5 VNW pch L=4e-08 W=4e-07 
M15 5 D VDD VNW pch L=4e-08 W=4e-07 
M16 10 C 5 VNW pch L=4e-08 W=4e-07 
M17 Y 1 10 VNW pch L=4e-08 W=4e-07 
M18 11 1 Y VNW pch L=4e-08 W=4e-07 
M19 5 C 11 VNW pch L=4e-08 W=4e-07 
M20 12 C 5 VNW pch L=4e-08 W=4e-07 
M21 Y 1 12 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT NOR4BB_X4M_A9TR Y VDD VNW VPW VSS AN BN C D
M0 17 BN VSS VPW nch L=4e-08 W=2.7e-07 
M1 3 AN 17 VPW nch L=4e-08 W=2.7e-07 
M2 18 AN 3 VPW nch L=4e-08 W=2.7e-07 
M3 VSS BN 18 VPW nch L=4e-08 W=2.7e-07 
M4 Y D VSS VPW nch L=4e-08 W=2.2e-07 
M5 VSS C Y VPW nch L=4e-08 W=2.2e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=2.2e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=2.2e-07 
M8 Y C VSS VPW nch L=4e-08 W=2.2e-07 
M9 VSS D Y VPW nch L=4e-08 W=2.2e-07 
M10 3 BN VDD VNW pch L=4e-08 W=2.3e-07 
M11 VDD AN 3 VNW pch L=4e-08 W=2.3e-07 
M12 3 AN VDD VNW pch L=4e-08 W=2.3e-07 
M13 VDD BN 3 VNW pch L=4e-08 W=2.3e-07 
M14 9 D VDD VNW pch L=4e-08 W=4e-07 
M15 10 C 9 VNW pch L=4e-08 W=4e-07 
M16 Y 3 10 VNW pch L=4e-08 W=4e-07 
M17 11 3 Y VNW pch L=4e-08 W=4e-07 
M18 12 C 11 VNW pch L=4e-08 W=4e-07 
M19 VDD D 12 VNW pch L=4e-08 W=4e-07 
M20 13 D VDD VNW pch L=4e-08 W=4e-07 
M21 14 C 13 VNW pch L=4e-08 W=4e-07 
M22 Y 3 14 VNW pch L=4e-08 W=4e-07 
M23 15 3 Y VNW pch L=4e-08 W=4e-07 
M24 16 C 15 VNW pch L=4e-08 W=4e-07 
M25 VDD D 16 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA1B2_X0P5M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 2 B0 VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B1 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y A0N VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS 2 Y VPW nch L=4e-08 W=1.2e-07 
M4 8 B0 2 VNW pch L=4e-08 W=2e-07 
M5 VDD B1 8 VNW pch L=4e-08 W=2e-07 
M6 9 A0N VDD VNW pch L=4e-08 W=2e-07 
M7 Y 2 9 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OA1B2_X0P7M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 2 B0 VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B1 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y A0N VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS 2 Y VPW nch L=4e-08 W=1.2e-07 
M4 8 B0 2 VNW pch L=4e-08 W=2.3e-07 
M5 VDD B1 8 VNW pch L=4e-08 W=2.3e-07 
M6 9 A0N VDD VNW pch L=4e-08 W=2.95e-07 
M7 Y 2 9 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT OA1B2_X1M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 2 B0 VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B1 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS 2 Y VPW nch L=4e-08 W=1.6e-07 
M4 8 B0 2 VNW pch L=4e-08 W=2.7e-07 
M5 VDD B1 8 VNW pch L=4e-08 W=2.7e-07 
M6 9 A0N VDD VNW pch L=4e-08 W=4e-07 
M7 Y 2 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA1B2_X1P4M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 2 B0 VSS VPW nch L=4e-08 W=1.4e-07 
M1 VSS B1 2 VPW nch L=4e-08 W=1.4e-07 
M2 Y A0N VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS 2 Y VPW nch L=4e-08 W=1.2e-07 
M4 Y 2 VSS VPW nch L=4e-08 W=1.2e-07 
M5 VSS A0N Y VPW nch L=4e-08 W=1.2e-07 
M6 8 B0 2 VNW pch L=4e-08 W=3.55e-07 
M7 VDD B1 8 VNW pch L=4e-08 W=3.55e-07 
M8 9 A0N VDD VNW pch L=4e-08 W=2.85e-07 
M9 Y 2 9 VNW pch L=4e-08 W=2.85e-07 
M10 10 2 Y VNW pch L=4e-08 W=2.85e-07 
M11 VDD A0N 10 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA1B2_X2M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 2 B0 VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS B1 2 VPW nch L=4e-08 W=1.6e-07 
M2 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS 2 Y VPW nch L=4e-08 W=1.6e-07 
M4 Y 2 VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M6 8 B0 2 VNW pch L=4e-08 W=4e-07 
M7 VDD B1 8 VNW pch L=4e-08 W=4e-07 
M8 9 A0N VDD VNW pch L=4e-08 W=4e-07 
M9 Y 2 9 VNW pch L=4e-08 W=4e-07 
M10 10 2 Y VNW pch L=4e-08 W=4e-07 
M11 VDD A0N 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA1B2_X3M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 3 B1 VSS VPW nch L=4e-08 W=1.45e-07 
M1 VSS B0 3 VPW nch L=4e-08 W=1.45e-07 
M2 3 B0 VSS VPW nch L=4e-08 W=1.45e-07 
M3 VSS B1 3 VPW nch L=4e-08 W=1.45e-07 
M4 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M8 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M10 8 B1 VDD VNW pch L=4e-08 W=3.6e-07 
M11 3 B0 8 VNW pch L=4e-08 W=3.6e-07 
M12 9 B0 3 VNW pch L=4e-08 W=3.6e-07 
M13 VDD B1 9 VNW pch L=4e-08 W=3.6e-07 
M14 10 A0N VDD VNW pch L=4e-08 W=4e-07 
M15 Y 3 10 VNW pch L=4e-08 W=4e-07 
M16 11 3 Y VNW pch L=4e-08 W=4e-07 
M17 VDD A0N 11 VNW pch L=4e-08 W=4e-07 
M18 12 A0N VDD VNW pch L=4e-08 W=4e-07 
M19 Y 3 12 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA1B2_X4M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 2 B0 VSS VPW nch L=4e-08 W=1.4e-07 
M1 VSS B1 2 VPW nch L=4e-08 W=1.4e-07 
M2 2 B1 VSS VPW nch L=4e-08 W=1.4e-07 
M3 VSS B0 2 VPW nch L=4e-08 W=1.4e-07 
M4 2 B0 VSS VPW nch L=4e-08 W=1.4e-07 
M5 VSS B1 2 VPW nch L=4e-08 W=1.4e-07 
M6 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS 2 Y VPW nch L=4e-08 W=1.6e-07 
M8 Y 2 VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M10 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M11 VSS 2 Y VPW nch L=4e-08 W=1.6e-07 
M12 Y 2 VSS VPW nch L=4e-08 W=1.6e-07 
M13 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M14 8 B0 2 VNW pch L=4e-08 W=3.4e-07 
M15 VDD B1 8 VNW pch L=4e-08 W=3.4e-07 
M16 9 B1 VDD VNW pch L=4e-08 W=3.4e-07 
M17 2 B0 9 VNW pch L=4e-08 W=3.4e-07 
M18 10 B0 2 VNW pch L=4e-08 W=3.4e-07 
M19 VDD B1 10 VNW pch L=4e-08 W=3.4e-07 
M20 11 A0N VDD VNW pch L=4e-08 W=4e-07 
M21 Y 2 11 VNW pch L=4e-08 W=4e-07 
M22 12 2 Y VNW pch L=4e-08 W=4e-07 
M23 VDD A0N 12 VNW pch L=4e-08 W=4e-07 
M24 13 A0N VDD VNW pch L=4e-08 W=4e-07 
M25 Y 2 13 VNW pch L=4e-08 W=4e-07 
M26 14 2 Y VNW pch L=4e-08 W=4e-07 
M27 VDD A0N 14 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA1B2_X6M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 3 B0 VSS VPW nch L=4e-08 W=2e-07 
M1 VSS B1 3 VPW nch L=4e-08 W=2e-07 
M2 3 B1 VSS VPW nch L=4e-08 W=2e-07 
M3 VSS B0 3 VPW nch L=4e-08 W=2e-07 
M4 3 B0 VSS VPW nch L=4e-08 W=2e-07 
M5 VSS B1 3 VPW nch L=4e-08 W=2e-07 
M6 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M10 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M11 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M12 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M13 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M14 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M15 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M16 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M17 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M18 8 B1 VDD VNW pch L=4e-08 W=3.7e-07 
M19 3 B0 8 VNW pch L=4e-08 W=3.7e-07 
M20 9 B0 3 VNW pch L=4e-08 W=3.7e-07 
M21 VDD B1 9 VNW pch L=4e-08 W=3.7e-07 
M22 10 B1 VDD VNW pch L=4e-08 W=3.7e-07 
M23 3 B0 10 VNW pch L=4e-08 W=3.7e-07 
M24 11 B0 3 VNW pch L=4e-08 W=3.7e-07 
M25 VDD B1 11 VNW pch L=4e-08 W=3.7e-07 
M26 12 A0N VDD VNW pch L=4e-08 W=4e-07 
M27 Y 3 12 VNW pch L=4e-08 W=4e-07 
M28 13 3 Y VNW pch L=4e-08 W=4e-07 
M29 VDD A0N 13 VNW pch L=4e-08 W=4e-07 
M30 14 A0N VDD VNW pch L=4e-08 W=4e-07 
M31 Y 3 14 VNW pch L=4e-08 W=4e-07 
M32 15 3 Y VNW pch L=4e-08 W=4e-07 
M33 VDD A0N 15 VNW pch L=4e-08 W=4e-07 
M34 16 A0N VDD VNW pch L=4e-08 W=4e-07 
M35 Y 3 16 VNW pch L=4e-08 W=4e-07 
M36 17 3 Y VNW pch L=4e-08 W=4e-07 
M37 VDD A0N 17 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA1B2_X8M_A9TR Y VDD VNW VPW VSS A0N B0 B1
M0 1 B0 VSS VPW nch L=4e-08 W=2.5e-07 
M1 VSS B1 1 VPW nch L=4e-08 W=2.5e-07 
M2 1 B1 VSS VPW nch L=4e-08 W=2.5e-07 
M3 VSS B0 1 VPW nch L=4e-08 W=2.5e-07 
M4 1 B0 VSS VPW nch L=4e-08 W=2.5e-07 
M5 VSS B1 1 VPW nch L=4e-08 W=2.5e-07 
M6 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M10 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M11 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M13 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M14 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M15 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M16 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M17 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M18 Y A0N VSS VPW nch L=4e-08 W=1.6e-07 
M19 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M20 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M21 VSS A0N Y VPW nch L=4e-08 W=1.6e-07 
M22 8 B0 1 VNW pch L=4e-08 W=3.7e-07 
M23 VDD B1 8 VNW pch L=4e-08 W=3.7e-07 
M24 9 B1 VDD VNW pch L=4e-08 W=3.7e-07 
M25 1 B0 9 VNW pch L=4e-08 W=3.7e-07 
M26 10 B0 1 VNW pch L=4e-08 W=3.7e-07 
M27 VDD B1 10 VNW pch L=4e-08 W=3.7e-07 
M28 11 B1 VDD VNW pch L=4e-08 W=3.7e-07 
M29 1 B0 11 VNW pch L=4e-08 W=3.7e-07 
M30 12 B0 1 VNW pch L=4e-08 W=3.7e-07 
M31 VDD B1 12 VNW pch L=4e-08 W=3.7e-07 
M32 13 A0N VDD VNW pch L=4e-08 W=4e-07 
M33 Y 1 13 VNW pch L=4e-08 W=4e-07 
M34 14 1 Y VNW pch L=4e-08 W=4e-07 
M35 VDD A0N 14 VNW pch L=4e-08 W=4e-07 
M36 15 A0N VDD VNW pch L=4e-08 W=4e-07 
M37 Y 1 15 VNW pch L=4e-08 W=4e-07 
M38 16 1 Y VNW pch L=4e-08 W=4e-07 
M39 VDD A0N 16 VNW pch L=4e-08 W=4e-07 
M40 17 A0N VDD VNW pch L=4e-08 W=4e-07 
M41 Y 1 17 VNW pch L=4e-08 W=4e-07 
M42 18 1 Y VNW pch L=4e-08 W=4e-07 
M43 VDD A0N 18 VNW pch L=4e-08 W=4e-07 
M44 19 A0N VDD VNW pch L=4e-08 W=4e-07 
M45 Y 1 19 VNW pch L=4e-08 W=4e-07 
M46 20 1 Y VNW pch L=4e-08 W=4e-07 
M47 VDD A0N 20 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA211_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=2.05e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.05e-07 
M2 11 B0 1 VPW nch L=4e-08 W=2.05e-07 
M3 4 C0 11 VPW nch L=4e-08 W=2.05e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=1.55e-07 
M5 10 A1 VDD VNW pch L=4e-08 W=2.6e-07 
M6 4 A0 10 VNW pch L=4e-08 W=2.6e-07 
M7 VDD B0 4 VNW pch L=4e-08 W=1.35e-07 
M8 4 C0 VDD VNW pch L=4e-08 W=1.35e-07 
M9 Y 4 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OA211_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=2.5e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.5e-07 
M2 11 B0 1 VPW nch L=4e-08 W=2.5e-07 
M3 4 C0 11 VPW nch L=4e-08 W=2.5e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=2.2e-07 
M5 10 A1 VDD VNW pch L=4e-08 W=3.25e-07 
M6 4 A0 10 VNW pch L=4e-08 W=3.25e-07 
M7 VDD B0 4 VNW pch L=4e-08 W=1.7e-07 
M8 4 C0 VDD VNW pch L=4e-08 W=1.7e-07 
M9 Y 4 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA211_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 11 B0 1 VPW nch L=4e-08 W=3.1e-07 
M3 4 C0 11 VPW nch L=4e-08 W=3.1e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M5 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M6 4 A0 10 VNW pch L=4e-08 W=4e-07 
M7 VDD B0 4 VNW pch L=4e-08 W=2.1e-07 
M8 4 C0 VDD VNW pch L=4e-08 W=2.1e-07 
M9 Y 4 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA211_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=2.35e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.35e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.35e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.35e-07 
M4 12 B0 1 VPW nch L=4e-08 W=2.35e-07 
M5 4 C0 12 VPW nch L=4e-08 W=2.35e-07 
M6 13 C0 4 VPW nch L=4e-08 W=2.35e-07 
M7 1 B0 13 VPW nch L=4e-08 W=2.35e-07 
M8 Y 4 VSS VPW nch L=4e-08 W=2.2e-07 
M9 VSS 4 Y VPW nch L=4e-08 W=2.2e-07 
M10 10 A1 VDD VNW pch L=4e-08 W=3.05e-07 
M11 4 A0 10 VNW pch L=4e-08 W=3.05e-07 
M12 11 A0 4 VNW pch L=4e-08 W=3.05e-07 
M13 VDD A1 11 VNW pch L=4e-08 W=3.05e-07 
M14 4 B0 VDD VNW pch L=4e-08 W=1.6e-07 
M15 VDD C0 4 VNW pch L=4e-08 W=1.6e-07 
M16 4 C0 VDD VNW pch L=4e-08 W=1.6e-07 
M17 VDD B0 4 VNW pch L=4e-08 W=1.6e-07 
M18 Y 4 VDD VNW pch L=4e-08 W=2.85e-07 
M19 VDD 4 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA211_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.05e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.05e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.05e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.05e-07 
M4 12 B0 1 VPW nch L=4e-08 W=3.05e-07 
M5 4 C0 12 VPW nch L=4e-08 W=3.05e-07 
M6 13 C0 4 VPW nch L=4e-08 W=3.05e-07 
M7 1 B0 13 VPW nch L=4e-08 W=3.05e-07 
M8 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M10 10 A1 VDD VNW pch L=4e-08 W=3.9e-07 
M11 4 A0 10 VNW pch L=4e-08 W=3.9e-07 
M12 11 A0 4 VNW pch L=4e-08 W=3.9e-07 
M13 VDD A1 11 VNW pch L=4e-08 W=3.9e-07 
M14 4 B0 VDD VNW pch L=4e-08 W=2e-07 
M15 VDD C0 4 VNW pch L=4e-08 W=2e-07 
M16 4 C0 VDD VNW pch L=4e-08 W=2e-07 
M17 VDD B0 4 VNW pch L=4e-08 W=2e-07 
M18 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA211_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 13 B0 1 VPW nch L=4e-08 W=3.1e-07 
M7 4 C0 13 VPW nch L=4e-08 W=3.1e-07 
M8 14 C0 4 VPW nch L=4e-08 W=3.1e-07 
M9 1 B0 14 VPW nch L=4e-08 W=3.1e-07 
M10 15 B0 1 VPW nch L=4e-08 W=3.1e-07 
M11 4 C0 15 VPW nch L=4e-08 W=3.1e-07 
M12 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M15 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M16 4 A0 10 VNW pch L=4e-08 W=4e-07 
M17 11 A0 4 VNW pch L=4e-08 W=4e-07 
M18 VDD A1 11 VNW pch L=4e-08 W=4e-07 
M19 12 A1 VDD VNW pch L=4e-08 W=4e-07 
M20 4 A0 12 VNW pch L=4e-08 W=4e-07 
M21 VDD B0 4 VNW pch L=4e-08 W=2.1e-07 
M22 4 C0 VDD VNW pch L=4e-08 W=2.1e-07 
M23 VDD C0 4 VNW pch L=4e-08 W=2.1e-07 
M24 4 B0 VDD VNW pch L=4e-08 W=2.1e-07 
M25 VDD B0 4 VNW pch L=4e-08 W=2.1e-07 
M26 4 C0 VDD VNW pch L=4e-08 W=2.1e-07 
M27 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M29 Y 4 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA211_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M8 14 B0 1 VPW nch L=4e-08 W=3.1e-07 
M9 4 C0 14 VPW nch L=4e-08 W=3.1e-07 
M10 15 C0 4 VPW nch L=4e-08 W=3.1e-07 
M11 1 B0 15 VPW nch L=4e-08 W=3.1e-07 
M12 16 B0 1 VPW nch L=4e-08 W=3.1e-07 
M13 4 C0 16 VPW nch L=4e-08 W=3.1e-07 
M14 17 C0 4 VPW nch L=4e-08 W=3.1e-07 
M15 1 B0 17 VPW nch L=4e-08 W=3.1e-07 
M16 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M18 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M20 10 A1 VDD VNW pch L=4e-08 W=3.95e-07 
M21 4 A0 10 VNW pch L=4e-08 W=3.95e-07 
M22 11 A0 4 VNW pch L=4e-08 W=3.95e-07 
M23 VDD A1 11 VNW pch L=4e-08 W=3.95e-07 
M24 12 A1 VDD VNW pch L=4e-08 W=3.95e-07 
M25 4 A0 12 VNW pch L=4e-08 W=3.95e-07 
M26 13 A0 4 VNW pch L=4e-08 W=3.95e-07 
M27 VDD A1 13 VNW pch L=4e-08 W=3.95e-07 
M28 4 B0 VDD VNW pch L=4e-08 W=2.05e-07 
M29 VDD C0 4 VNW pch L=4e-08 W=2.05e-07 
M30 4 C0 VDD VNW pch L=4e-08 W=2.05e-07 
M31 VDD B0 4 VNW pch L=4e-08 W=2.05e-07 
M32 4 B0 VDD VNW pch L=4e-08 W=2.05e-07 
M33 VDD C0 4 VNW pch L=4e-08 W=2.05e-07 
M34 4 C0 VDD VNW pch L=4e-08 W=2.05e-07 
M35 VDD B0 4 VNW pch L=4e-08 W=2.05e-07 
M36 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M38 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA211_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M8 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M9 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M11 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M12 16 B0 1 VPW nch L=4e-08 W=3.7e-07 
M13 4 C0 16 VPW nch L=4e-08 W=3.7e-07 
M14 17 C0 4 VPW nch L=4e-08 W=3.7e-07 
M15 1 B0 17 VPW nch L=4e-08 W=3.7e-07 
M16 18 B0 1 VPW nch L=4e-08 W=3.7e-07 
M17 4 C0 18 VPW nch L=4e-08 W=3.7e-07 
M18 19 C0 4 VPW nch L=4e-08 W=3.7e-07 
M19 1 B0 19 VPW nch L=4e-08 W=3.7e-07 
M20 20 B0 1 VPW nch L=4e-08 W=3.7e-07 
M21 4 C0 20 VPW nch L=4e-08 W=3.7e-07 
M22 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M23 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M24 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M25 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M26 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M27 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M28 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M29 4 A0 10 VNW pch L=4e-08 W=4e-07 
M30 11 A0 4 VNW pch L=4e-08 W=4e-07 
M31 VDD A1 11 VNW pch L=4e-08 W=4e-07 
M32 12 A1 VDD VNW pch L=4e-08 W=4e-07 
M33 4 A0 12 VNW pch L=4e-08 W=4e-07 
M34 13 A0 4 VNW pch L=4e-08 W=4e-07 
M35 VDD A1 13 VNW pch L=4e-08 W=4e-07 
M36 14 A1 VDD VNW pch L=4e-08 W=4e-07 
M37 4 A0 14 VNW pch L=4e-08 W=4e-07 
M38 15 A0 4 VNW pch L=4e-08 W=4e-07 
M39 VDD A1 15 VNW pch L=4e-08 W=4e-07 
M40 4 B0 VDD VNW pch L=4e-08 W=2.5e-07 
M41 VDD C0 4 VNW pch L=4e-08 W=2.5e-07 
M42 4 C0 VDD VNW pch L=4e-08 W=2.5e-07 
M43 VDD B0 4 VNW pch L=4e-08 W=2.5e-07 
M44 4 B0 VDD VNW pch L=4e-08 W=2.5e-07 
M45 VDD C0 4 VNW pch L=4e-08 W=2.5e-07 
M46 4 C0 VDD VNW pch L=4e-08 W=2.5e-07 
M47 VDD B0 4 VNW pch L=4e-08 W=2.5e-07 
M48 4 B0 VDD VNW pch L=4e-08 W=2.5e-07 
M49 VDD C0 4 VNW pch L=4e-08 W=2.5e-07 
M50 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M51 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M52 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M53 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M54 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M55 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21A1OI2_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A0 1 VPW nch L=4e-08 W=1.2e-07 
M1 1 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 Y B0 1 VPW nch L=4e-08 W=1.2e-07 
M3 VSS C0 Y VPW nch L=4e-08 W=1.2e-07 
M4 10 A0 2 VNW pch L=4e-08 W=2e-07 
M5 VDD A1 10 VNW pch L=4e-08 W=2e-07 
M6 2 B0 VDD VNW pch L=4e-08 W=1.35e-07 
M7 Y C0 2 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OA21A1OI2_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A0 1 VPW nch L=4e-08 W=1.2e-07 
M1 1 A1 VSS VPW nch L=4e-08 W=1.2e-07 
M2 Y B0 1 VPW nch L=4e-08 W=1.2e-07 
M3 VSS C0 Y VPW nch L=4e-08 W=1.2e-07 
M4 10 A0 2 VNW pch L=4e-08 W=2.85e-07 
M5 VDD A1 10 VNW pch L=4e-08 W=2.85e-07 
M6 2 B0 VDD VNW pch L=4e-08 W=1.9e-07 
M7 Y C0 2 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA21A1OI2_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=1.8e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=1.8e-07 
M2 Y B0 1 VPW nch L=4e-08 W=1.8e-07 
M3 Y C0 VSS VPW nch L=4e-08 W=1.2e-07 
M4 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M5 4 A0 10 VNW pch L=4e-08 W=4e-07 
M6 VDD B0 4 VNW pch L=4e-08 W=3e-07 
M7 Y C0 4 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21A1OI2_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A0 2 VPW nch L=4e-08 W=2.3e-07 
M1 2 A1 VSS VPW nch L=4e-08 W=2.3e-07 
M2 Y B0 2 VPW nch L=4e-08 W=2.3e-07 
M3 VSS C0 Y VPW nch L=4e-08 W=1.5e-07 
M4 10 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M5 3 A0 10 VNW pch L=4e-08 W=2.85e-07 
M6 11 A0 3 VNW pch L=4e-08 W=2.85e-07 
M7 VDD A1 11 VNW pch L=4e-08 W=2.85e-07 
M8 3 B0 VDD VNW pch L=4e-08 W=3.8e-07 
M9 Y C0 3 VNW pch L=4e-08 W=2.85e-07 
M10 3 C0 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA21A1OI2_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A0 1 VPW nch L=4e-08 W=1.6e-07 
M1 1 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M2 VSS A1 1 VPW nch L=4e-08 W=1.6e-07 
M3 1 A0 VSS VPW nch L=4e-08 W=1.6e-07 
M4 Y B0 1 VPW nch L=4e-08 W=1.6e-07 
M5 1 B0 Y VPW nch L=4e-08 W=1.6e-07 
M6 VSS C0 Y VPW nch L=4e-08 W=2.1e-07 
M7 10 A0 2 VNW pch L=4e-08 W=4e-07 
M8 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M9 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M10 2 A0 11 VNW pch L=4e-08 W=4e-07 
M11 VDD B0 2 VNW pch L=4e-08 W=2.65e-07 
M12 2 B0 VDD VNW pch L=4e-08 W=2.65e-07 
M13 Y C0 2 VNW pch L=4e-08 W=4e-07 
M14 2 C0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21A1OI2_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 4 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1 4 VPW nch L=4e-08 W=2.4e-07 
M2 VSS A0 4 VPW nch L=4e-08 W=2.4e-07 
M3 4 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M4 Y B0 4 VPW nch L=4e-08 W=2.4e-07 
M5 4 B0 Y VPW nch L=4e-08 W=2.4e-07 
M6 Y C0 VSS VPW nch L=4e-08 W=3.15e-07 
M7 3 A1 VDD VNW pch L=4e-08 W=4e-07 
M8 VDD A1 3 VNW pch L=4e-08 W=4e-07 
M9 3 A1 VDD VNW pch L=4e-08 W=4e-07 
M10 5 A0 3 VNW pch L=4e-08 W=4e-07 
M11 3 A0 5 VNW pch L=4e-08 W=4e-07 
M12 5 A0 3 VNW pch L=4e-08 W=4e-07 
M13 VDD B0 5 VNW pch L=4e-08 W=4e-07 
M14 5 B0 VDD VNW pch L=4e-08 W=4e-07 
M15 Y C0 5 VNW pch L=4e-08 W=4e-07 
M16 5 C0 Y VNW pch L=4e-08 W=4e-07 
M17 Y C0 5 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21A1OI2_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 3 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS A1 3 VPW nch L=4e-08 W=1.6e-07 
M2 3 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS A1 3 VPW nch L=4e-08 W=1.6e-07 
M4 3 A0 VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS A0 3 VPW nch L=4e-08 W=1.6e-07 
M6 3 A0 VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS A0 3 VPW nch L=4e-08 W=1.6e-07 
M8 Y B0 3 VPW nch L=4e-08 W=2.2e-07 
M9 3 B0 Y VPW nch L=4e-08 W=2.2e-07 
M10 Y B0 3 VPW nch L=4e-08 W=2.2e-07 
M11 VSS C0 Y VPW nch L=4e-08 W=2.1e-07 
M12 Y C0 VSS VPW nch L=4e-08 W=2.1e-07 
M13 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M14 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M16 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M17 5 A0 2 VNW pch L=4e-08 W=4e-07 
M18 2 A0 5 VNW pch L=4e-08 W=4e-07 
M19 5 A0 2 VNW pch L=4e-08 W=4e-07 
M20 2 A0 5 VNW pch L=4e-08 W=4e-07 
M21 5 B0 VDD VNW pch L=4e-08 W=3.6e-07 
M22 VDD B0 5 VNW pch L=4e-08 W=3.6e-07 
M23 5 B0 VDD VNW pch L=4e-08 W=3.6e-07 
M24 Y C0 5 VNW pch L=4e-08 W=4e-07 
M25 5 C0 Y VNW pch L=4e-08 W=4e-07 
M26 Y C0 5 VNW pch L=4e-08 W=4e-07 
M27 5 C0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21A1OI2_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 3 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS A1 3 VPW nch L=4e-08 W=1.6e-07 
M2 3 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS A1 3 VPW nch L=4e-08 W=1.6e-07 
M4 3 A1 VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS A1 3 VPW nch L=4e-08 W=1.6e-07 
M6 3 A0 VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS A0 3 VPW nch L=4e-08 W=1.6e-07 
M8 3 A0 VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS A0 3 VPW nch L=4e-08 W=1.6e-07 
M10 3 A0 VSS VPW nch L=4e-08 W=1.6e-07 
M11 VSS A0 3 VPW nch L=4e-08 W=1.6e-07 
M12 Y B0 3 VPW nch L=4e-08 W=3.2e-07 
M13 3 B0 Y VPW nch L=4e-08 W=3.2e-07 
M14 Y B0 3 VPW nch L=4e-08 W=3.2e-07 
M15 Y C0 VSS VPW nch L=4e-08 W=3.15e-07 
M16 VSS C0 Y VPW nch L=4e-08 W=3.15e-07 
M17 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M18 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M20 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD A1 2 VNW pch L=4e-08 W=4e-07 
M22 2 A1 VDD VNW pch L=4e-08 W=4e-07 
M23 5 A0 2 VNW pch L=4e-08 W=4e-07 
M24 2 A0 5 VNW pch L=4e-08 W=4e-07 
M25 5 A0 2 VNW pch L=4e-08 W=4e-07 
M26 2 A0 5 VNW pch L=4e-08 W=4e-07 
M27 5 A0 2 VNW pch L=4e-08 W=4e-07 
M28 2 A0 5 VNW pch L=4e-08 W=4e-07 
M29 VDD B0 5 VNW pch L=4e-08 W=3.95e-07 
M30 5 B0 VDD VNW pch L=4e-08 W=3.95e-07 
M31 VDD B0 5 VNW pch L=4e-08 W=3.95e-07 
M32 5 B0 VDD VNW pch L=4e-08 W=3.95e-07 
M33 Y C0 5 VNW pch L=4e-08 W=4e-07 
M34 5 C0 Y VNW pch L=4e-08 W=4e-07 
M35 Y C0 5 VNW pch L=4e-08 W=4e-07 
M36 5 C0 Y VNW pch L=4e-08 W=4e-07 
M37 Y C0 5 VNW pch L=4e-08 W=4e-07 
M38 5 C0 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21B_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 2 A0 VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS A1 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS B0N Y VPW nch L=4e-08 W=1.2e-07 
M4 8 A0 2 VNW pch L=4e-08 W=2e-07 
M5 VDD A1 8 VNW pch L=4e-08 W=2e-07 
M6 9 2 VDD VNW pch L=4e-08 W=2e-07 
M7 Y B0N 9 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OA21B_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 2 A0 VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS A1 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS B0N Y VPW nch L=4e-08 W=1.2e-07 
M4 8 A0 2 VNW pch L=4e-08 W=2.3e-07 
M5 VDD A1 8 VNW pch L=4e-08 W=2.3e-07 
M6 9 2 VDD VNW pch L=4e-08 W=2.95e-07 
M7 Y B0N 9 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT OA21B_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 2 A0 VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS A1 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M4 8 A0 2 VNW pch L=4e-08 W=2.7e-07 
M5 VDD A1 8 VNW pch L=4e-08 W=2.7e-07 
M6 9 2 VDD VNW pch L=4e-08 W=4e-07 
M7 Y B0N 9 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21B_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 2 A0 VSS VPW nch L=4e-08 W=1.4e-07 
M1 VSS A1 2 VPW nch L=4e-08 W=1.4e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=1.2e-07 
M3 VSS B0N Y VPW nch L=4e-08 W=1.2e-07 
M4 Y B0N VSS VPW nch L=4e-08 W=1.2e-07 
M5 VSS 2 Y VPW nch L=4e-08 W=1.2e-07 
M6 8 A0 2 VNW pch L=4e-08 W=3.55e-07 
M7 VDD A1 8 VNW pch L=4e-08 W=3.55e-07 
M8 9 2 VDD VNW pch L=4e-08 W=2.85e-07 
M9 Y B0N 9 VNW pch L=4e-08 W=2.85e-07 
M10 10 B0N Y VNW pch L=4e-08 W=2.85e-07 
M11 VDD 2 10 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA21B_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 2 A0 VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS A1 2 VPW nch L=4e-08 W=1.6e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M4 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS 2 Y VPW nch L=4e-08 W=1.6e-07 
M6 8 A0 2 VNW pch L=4e-08 W=4e-07 
M7 VDD A1 8 VNW pch L=4e-08 W=4e-07 
M8 9 2 VDD VNW pch L=4e-08 W=4e-07 
M9 Y B0N 9 VNW pch L=4e-08 W=4e-07 
M10 10 B0N Y VNW pch L=4e-08 W=4e-07 
M11 VDD 2 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21B_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 A1 VSS VPW nch L=4e-08 W=1.45e-07 
M1 VSS A0 3 VPW nch L=4e-08 W=1.45e-07 
M2 3 A0 VSS VPW nch L=4e-08 W=1.45e-07 
M3 VSS A1 3 VPW nch L=4e-08 W=1.45e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M5 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M6 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M8 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M10 8 A1 VDD VNW pch L=4e-08 W=3.6e-07 
M11 3 A0 8 VNW pch L=4e-08 W=3.6e-07 
M12 9 A0 3 VNW pch L=4e-08 W=3.6e-07 
M13 VDD A1 9 VNW pch L=4e-08 W=3.6e-07 
M14 10 3 VDD VNW pch L=4e-08 W=4e-07 
M15 Y B0N 10 VNW pch L=4e-08 W=4e-07 
M16 11 B0N Y VNW pch L=4e-08 W=4e-07 
M17 VDD 3 11 VNW pch L=4e-08 W=4e-07 
M18 12 3 VDD VNW pch L=4e-08 W=4e-07 
M19 Y B0N 12 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21B_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 2 A0 VSS VPW nch L=4e-08 W=1.4e-07 
M1 VSS A1 2 VPW nch L=4e-08 W=1.4e-07 
M2 2 A1 VSS VPW nch L=4e-08 W=1.4e-07 
M3 VSS A0 2 VPW nch L=4e-08 W=1.4e-07 
M4 2 A0 VSS VPW nch L=4e-08 W=1.4e-07 
M5 VSS A1 2 VPW nch L=4e-08 W=1.4e-07 
M6 Y 2 VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M8 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS 2 Y VPW nch L=4e-08 W=1.6e-07 
M10 Y 2 VSS VPW nch L=4e-08 W=1.6e-07 
M11 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M12 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M13 VSS 2 Y VPW nch L=4e-08 W=1.6e-07 
M14 8 A0 2 VNW pch L=4e-08 W=3.4e-07 
M15 VDD A1 8 VNW pch L=4e-08 W=3.4e-07 
M16 9 A1 VDD VNW pch L=4e-08 W=3.4e-07 
M17 2 A0 9 VNW pch L=4e-08 W=3.4e-07 
M18 10 A0 2 VNW pch L=4e-08 W=3.4e-07 
M19 VDD A1 10 VNW pch L=4e-08 W=3.4e-07 
M20 11 2 VDD VNW pch L=4e-08 W=4e-07 
M21 Y B0N 11 VNW pch L=4e-08 W=4e-07 
M22 12 B0N Y VNW pch L=4e-08 W=4e-07 
M23 VDD 2 12 VNW pch L=4e-08 W=4e-07 
M24 13 2 VDD VNW pch L=4e-08 W=4e-07 
M25 Y B0N 13 VNW pch L=4e-08 W=4e-07 
M26 14 B0N Y VNW pch L=4e-08 W=4e-07 
M27 VDD 2 14 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21B_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 3 A0 VSS VPW nch L=4e-08 W=2e-07 
M1 VSS A1 3 VPW nch L=4e-08 W=2e-07 
M2 3 A1 VSS VPW nch L=4e-08 W=2e-07 
M3 VSS A0 3 VPW nch L=4e-08 W=2e-07 
M4 3 A0 VSS VPW nch L=4e-08 W=2e-07 
M5 VSS A1 3 VPW nch L=4e-08 W=2e-07 
M6 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M8 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M10 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M11 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M12 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M13 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M14 Y 3 VSS VPW nch L=4e-08 W=1.6e-07 
M15 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M16 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M17 VSS 3 Y VPW nch L=4e-08 W=1.6e-07 
M18 8 A1 VDD VNW pch L=4e-08 W=3.7e-07 
M19 3 A0 8 VNW pch L=4e-08 W=3.7e-07 
M20 9 A0 3 VNW pch L=4e-08 W=3.7e-07 
M21 VDD A1 9 VNW pch L=4e-08 W=3.7e-07 
M22 10 A1 VDD VNW pch L=4e-08 W=3.7e-07 
M23 3 A0 10 VNW pch L=4e-08 W=3.7e-07 
M24 11 A0 3 VNW pch L=4e-08 W=3.7e-07 
M25 VDD A1 11 VNW pch L=4e-08 W=3.7e-07 
M26 12 3 VDD VNW pch L=4e-08 W=4e-07 
M27 Y B0N 12 VNW pch L=4e-08 W=4e-07 
M28 13 B0N Y VNW pch L=4e-08 W=4e-07 
M29 VDD 3 13 VNW pch L=4e-08 W=4e-07 
M30 14 3 VDD VNW pch L=4e-08 W=4e-07 
M31 Y B0N 14 VNW pch L=4e-08 W=4e-07 
M32 15 B0N Y VNW pch L=4e-08 W=4e-07 
M33 VDD 3 15 VNW pch L=4e-08 W=4e-07 
M34 16 3 VDD VNW pch L=4e-08 W=4e-07 
M35 Y B0N 16 VNW pch L=4e-08 W=4e-07 
M36 17 B0N Y VNW pch L=4e-08 W=4e-07 
M37 VDD 3 17 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21B_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 1 A0 VSS VPW nch L=4e-08 W=2.5e-07 
M1 VSS A1 1 VPW nch L=4e-08 W=2.5e-07 
M2 1 A1 VSS VPW nch L=4e-08 W=2.5e-07 
M3 VSS A0 1 VPW nch L=4e-08 W=2.5e-07 
M4 1 A0 VSS VPW nch L=4e-08 W=2.5e-07 
M5 VSS A1 1 VPW nch L=4e-08 W=2.5e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M7 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M8 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M11 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M12 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M13 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M14 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M15 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M16 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M17 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M18 Y 1 VSS VPW nch L=4e-08 W=1.6e-07 
M19 VSS B0N Y VPW nch L=4e-08 W=1.6e-07 
M20 Y B0N VSS VPW nch L=4e-08 W=1.6e-07 
M21 VSS 1 Y VPW nch L=4e-08 W=1.6e-07 
M22 8 A0 1 VNW pch L=4e-08 W=3.7e-07 
M23 VDD A1 8 VNW pch L=4e-08 W=3.7e-07 
M24 9 A1 VDD VNW pch L=4e-08 W=3.7e-07 
M25 1 A0 9 VNW pch L=4e-08 W=3.7e-07 
M26 10 A0 1 VNW pch L=4e-08 W=3.7e-07 
M27 VDD A1 10 VNW pch L=4e-08 W=3.7e-07 
M28 11 A1 VDD VNW pch L=4e-08 W=3.7e-07 
M29 1 A0 11 VNW pch L=4e-08 W=3.7e-07 
M30 12 A0 1 VNW pch L=4e-08 W=3.7e-07 
M31 VDD A1 12 VNW pch L=4e-08 W=3.7e-07 
M32 13 1 VDD VNW pch L=4e-08 W=4e-07 
M33 Y B0N 13 VNW pch L=4e-08 W=4e-07 
M34 14 B0N Y VNW pch L=4e-08 W=4e-07 
M35 VDD 1 14 VNW pch L=4e-08 W=4e-07 
M36 15 1 VDD VNW pch L=4e-08 W=4e-07 
M37 Y B0N 15 VNW pch L=4e-08 W=4e-07 
M38 16 B0N Y VNW pch L=4e-08 W=4e-07 
M39 VDD 1 16 VNW pch L=4e-08 W=4e-07 
M40 17 1 VDD VNW pch L=4e-08 W=4e-07 
M41 Y B0N 17 VNW pch L=4e-08 W=4e-07 
M42 18 B0N Y VNW pch L=4e-08 W=4e-07 
M43 VDD 1 18 VNW pch L=4e-08 W=4e-07 
M44 19 1 VDD VNW pch L=4e-08 W=4e-07 
M45 Y B0N 19 VNW pch L=4e-08 W=4e-07 
M46 20 B0N Y VNW pch L=4e-08 W=4e-07 
M47 VDD 1 20 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=1.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=1.4e-07 
M2 4 B0 1 VPW nch L=4e-08 W=1.4e-07 
M3 Y 4 VSS VPW nch L=4e-08 W=1.55e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=2.3e-07 
M5 4 A0 9 VNW pch L=4e-08 W=2.3e-07 
M6 VDD B0 4 VNW pch L=4e-08 W=1.2e-07 
M7 Y 4 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OA21_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=1.6e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=1.6e-07 
M2 4 B0 1 VPW nch L=4e-08 W=1.6e-07 
M3 Y 4 VSS VPW nch L=4e-08 W=2.2e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=2.7e-07 
M5 4 A0 9 VNW pch L=4e-08 W=2.7e-07 
M6 VDD B0 4 VNW pch L=4e-08 W=1.4e-07 
M7 Y 4 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA21_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=2.05e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.05e-07 
M2 4 B0 1 VPW nch L=4e-08 W=2.05e-07 
M3 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=3.4e-07 
M5 4 A0 9 VNW pch L=4e-08 W=3.4e-07 
M6 VDD B0 4 VNW pch L=4e-08 W=1.75e-07 
M7 Y 4 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 2 B0 1 VPW nch L=4e-08 W=3e-07 
M1 VSS A1 2 VPW nch L=4e-08 W=3e-07 
M2 2 A0 VSS VPW nch L=4e-08 W=3e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=2.2e-07 
M5 VDD B0 1 VNW pch L=4e-08 W=2.6e-07 
M6 9 A1 VDD VNW pch L=4e-08 W=2.5e-07 
M7 1 A0 9 VNW pch L=4e-08 W=2.5e-07 
M8 10 A0 1 VNW pch L=4e-08 W=2.5e-07 
M9 VDD A1 10 VNW pch L=4e-08 W=2.5e-07 
M10 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
M11 VDD 1 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA21_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=1.95e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=1.95e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=1.95e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=1.95e-07 
M4 4 B0 1 VPW nch L=4e-08 W=3.9e-07 
M5 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M7 9 A1 VDD VNW pch L=4e-08 W=3.2e-07 
M8 4 A0 9 VNW pch L=4e-08 W=3.2e-07 
M9 10 A0 4 VNW pch L=4e-08 W=3.2e-07 
M10 VDD A1 10 VNW pch L=4e-08 W=3.2e-07 
M11 4 B0 VDD VNW pch L=4e-08 W=3.3e-07 
M12 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M13 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 2 VPW nch L=4e-08 W=2.95e-07 
M1 2 A0 VSS VPW nch L=4e-08 W=2.95e-07 
M2 VSS A0 2 VPW nch L=4e-08 W=2.95e-07 
M3 2 A1 VSS VPW nch L=4e-08 W=2.95e-07 
M4 1 B0 2 VPW nch L=4e-08 W=2.95e-07 
M5 2 B0 1 VPW nch L=4e-08 W=2.95e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M9 9 A0 1 VNW pch L=4e-08 W=3.25e-07 
M10 VDD A1 9 VNW pch L=4e-08 W=3.25e-07 
M11 10 A1 VDD VNW pch L=4e-08 W=3.25e-07 
M12 1 A0 10 VNW pch L=4e-08 W=3.25e-07 
M13 11 A0 1 VNW pch L=4e-08 W=3.25e-07 
M14 VDD A1 11 VNW pch L=4e-08 W=3.25e-07 
M15 1 B0 VDD VNW pch L=4e-08 W=2.55e-07 
M16 VDD B0 1 VNW pch L=4e-08 W=2.55e-07 
M17 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M19 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 2 VPW nch L=4e-08 W=3.6e-07 
M1 2 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M2 VSS A0 2 VPW nch L=4e-08 W=3.6e-07 
M3 2 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M4 1 B0 2 VPW nch L=4e-08 W=3.6e-07 
M5 2 B0 1 VPW nch L=4e-08 W=3.6e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M10 9 A0 1 VNW pch L=4e-08 W=4e-07 
M11 VDD A1 9 VNW pch L=4e-08 W=4e-07 
M12 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 1 A0 10 VNW pch L=4e-08 W=4e-07 
M14 11 A0 1 VNW pch L=4e-08 W=4e-07 
M15 VDD A1 11 VNW pch L=4e-08 W=4e-07 
M16 1 B0 VDD VNW pch L=4e-08 W=3.15e-07 
M17 VDD B0 1 VNW pch L=4e-08 W=3.15e-07 
M18 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M20 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A0 3 VPW nch L=4e-08 W=3.75e-07 
M1 3 A1 VSS VPW nch L=4e-08 W=3.75e-07 
M2 VSS A1 3 VPW nch L=4e-08 W=3.75e-07 
M3 3 A0 VSS VPW nch L=4e-08 W=3.75e-07 
M4 VSS A0 3 VPW nch L=4e-08 W=3.75e-07 
M5 3 A1 VSS VPW nch L=4e-08 W=3.75e-07 
M6 1 B0 3 VPW nch L=4e-08 W=3.75e-07 
M7 3 B0 1 VPW nch L=4e-08 W=3.75e-07 
M8 1 B0 3 VPW nch L=4e-08 W=3.75e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M13 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M15 9 A0 1 VNW pch L=4e-08 W=3.75e-07 
M16 VDD A1 9 VNW pch L=4e-08 W=3.75e-07 
M17 10 A1 VDD VNW pch L=4e-08 W=3.75e-07 
M18 1 A0 10 VNW pch L=4e-08 W=3.75e-07 
M19 11 A0 1 VNW pch L=4e-08 W=3.75e-07 
M20 VDD A1 11 VNW pch L=4e-08 W=3.75e-07 
M21 12 A1 VDD VNW pch L=4e-08 W=3.75e-07 
M22 1 A0 12 VNW pch L=4e-08 W=3.75e-07 
M23 13 A0 1 VNW pch L=4e-08 W=3.75e-07 
M24 VDD A1 13 VNW pch L=4e-08 W=3.75e-07 
M25 1 B0 VDD VNW pch L=4e-08 W=3.25e-07 
M26 VDD B0 1 VNW pch L=4e-08 W=3.25e-07 
M27 1 B0 VDD VNW pch L=4e-08 W=3.25e-07 
M28 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M30 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M32 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M33 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA21_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 3 VPW nch L=4e-08 W=3.6e-07 
M1 3 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M2 VSS A0 3 VPW nch L=4e-08 W=3.6e-07 
M3 3 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M4 VSS A1 3 VPW nch L=4e-08 W=3.6e-07 
M5 3 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M6 VSS A0 3 VPW nch L=4e-08 W=3.6e-07 
M7 3 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M8 2 B0 3 VPW nch L=4e-08 W=3.6e-07 
M9 3 B0 2 VPW nch L=4e-08 W=3.6e-07 
M10 2 B0 3 VPW nch L=4e-08 W=3.6e-07 
M11 3 B0 2 VPW nch L=4e-08 W=3.6e-07 
M12 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M16 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M18 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M20 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M21 2 A0 9 VNW pch L=4e-08 W=4e-07 
M22 10 A0 2 VNW pch L=4e-08 W=4e-07 
M23 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M24 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M25 2 A0 11 VNW pch L=4e-08 W=4e-07 
M26 12 A0 2 VNW pch L=4e-08 W=4e-07 
M27 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M28 13 A1 VDD VNW pch L=4e-08 W=4e-07 
M29 2 A0 13 VNW pch L=4e-08 W=4e-07 
M30 14 A0 2 VNW pch L=4e-08 W=4e-07 
M31 VDD A1 14 VNW pch L=4e-08 W=4e-07 
M32 2 B0 VDD VNW pch L=4e-08 W=3.15e-07 
M33 VDD B0 2 VNW pch L=4e-08 W=3.15e-07 
M34 2 B0 VDD VNW pch L=4e-08 W=3.15e-07 
M35 VDD B0 2 VNW pch L=4e-08 W=3.15e-07 
M36 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M38 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M40 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M41 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M42 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M43 VDD 2 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA22_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=1.35e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=1.35e-07 
M2 4 B0 1 VPW nch L=4e-08 W=1.35e-07 
M3 1 B1 4 VPW nch L=4e-08 W=1.35e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=1.55e-07 
M5 10 A1 VDD VNW pch L=4e-08 W=2.25e-07 
M6 4 A0 10 VNW pch L=4e-08 W=2.25e-07 
M7 11 B0 4 VNW pch L=4e-08 W=2.25e-07 
M8 VDD B1 11 VNW pch L=4e-08 W=2.25e-07 
M9 Y 4 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OA22_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=1.8e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=1.8e-07 
M2 4 B0 1 VPW nch L=4e-08 W=1.8e-07 
M3 1 B1 4 VPW nch L=4e-08 W=1.8e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=2.2e-07 
M5 10 A1 VDD VNW pch L=4e-08 W=2.8e-07 
M6 4 A0 10 VNW pch L=4e-08 W=2.8e-07 
M7 11 B0 4 VNW pch L=4e-08 W=2.8e-07 
M8 VDD B1 11 VNW pch L=4e-08 W=2.8e-07 
M9 Y 4 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA22_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=2.15e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.15e-07 
M2 4 B0 1 VPW nch L=4e-08 W=2.15e-07 
M3 1 B1 4 VPW nch L=4e-08 W=2.15e-07 
M4 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M5 10 A1 VDD VNW pch L=4e-08 W=3.5e-07 
M6 4 A0 10 VNW pch L=4e-08 W=3.5e-07 
M7 11 B0 4 VNW pch L=4e-08 W=3.5e-07 
M8 VDD B1 11 VNW pch L=4e-08 W=3.5e-07 
M9 Y 4 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA22_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A0 2 VPW nch L=4e-08 W=3.4e-07 
M1 2 A1 VSS VPW nch L=4e-08 W=3.4e-07 
M2 3 B1 2 VPW nch L=4e-08 W=3.4e-07 
M3 2 B0 3 VPW nch L=4e-08 W=3.4e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=2.2e-07 
M5 VSS 3 Y VPW nch L=4e-08 W=2.2e-07 
M6 10 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M7 3 A0 10 VNW pch L=4e-08 W=2.85e-07 
M8 11 A0 3 VNW pch L=4e-08 W=2.85e-07 
M9 VDD A1 11 VNW pch L=4e-08 W=2.85e-07 
M10 12 B1 VDD VNW pch L=4e-08 W=2.85e-07 
M11 3 B0 12 VNW pch L=4e-08 W=2.85e-07 
M12 13 B0 3 VNW pch L=4e-08 W=2.85e-07 
M13 VDD B1 13 VNW pch L=4e-08 W=2.85e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=2.85e-07 
M15 VDD 3 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OA22_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=2.15e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.15e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.15e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.15e-07 
M4 4 B1 1 VPW nch L=4e-08 W=2.15e-07 
M5 1 B0 4 VPW nch L=4e-08 W=2.15e-07 
M6 4 B0 1 VPW nch L=4e-08 W=2.15e-07 
M7 1 B1 4 VPW nch L=4e-08 W=2.15e-07 
M8 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M10 10 A1 VDD VNW pch L=4e-08 W=3.55e-07 
M11 4 A0 10 VNW pch L=4e-08 W=3.55e-07 
M12 11 A0 4 VNW pch L=4e-08 W=3.55e-07 
M13 VDD A1 11 VNW pch L=4e-08 W=3.55e-07 
M14 12 B1 VDD VNW pch L=4e-08 W=3.55e-07 
M15 4 B0 12 VNW pch L=4e-08 W=3.55e-07 
M16 13 B0 4 VNW pch L=4e-08 W=3.55e-07 
M17 VDD B1 13 VNW pch L=4e-08 W=3.55e-07 
M18 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA22_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=2.25e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.25e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.25e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.25e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=2.25e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=2.25e-07 
M6 4 B0 1 VPW nch L=4e-08 W=2.25e-07 
M7 1 B1 4 VPW nch L=4e-08 W=2.25e-07 
M8 4 B1 1 VPW nch L=4e-08 W=2.25e-07 
M9 1 B0 4 VPW nch L=4e-08 W=2.25e-07 
M10 4 B0 1 VPW nch L=4e-08 W=2.25e-07 
M11 1 B1 4 VPW nch L=4e-08 W=2.25e-07 
M12 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M15 10 A1 VDD VNW pch L=4e-08 W=3.75e-07 
M16 4 A0 10 VNW pch L=4e-08 W=3.75e-07 
M17 11 A0 4 VNW pch L=4e-08 W=3.75e-07 
M18 VDD A1 11 VNW pch L=4e-08 W=3.75e-07 
M19 12 A1 VDD VNW pch L=4e-08 W=3.75e-07 
M20 4 A0 12 VNW pch L=4e-08 W=3.75e-07 
M21 13 B0 4 VNW pch L=4e-08 W=3.75e-07 
M22 VDD B1 13 VNW pch L=4e-08 W=3.75e-07 
M23 14 B1 VDD VNW pch L=4e-08 W=3.75e-07 
M24 4 B0 14 VNW pch L=4e-08 W=3.75e-07 
M25 15 B0 4 VNW pch L=4e-08 W=3.75e-07 
M26 VDD B1 15 VNW pch L=4e-08 W=3.75e-07 
M27 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M29 Y 4 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA22_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A0 2 VPW nch L=4e-08 W=2.85e-07 
M1 2 A1 VSS VPW nch L=4e-08 W=2.85e-07 
M2 VSS A1 2 VPW nch L=4e-08 W=2.85e-07 
M3 2 A0 VSS VPW nch L=4e-08 W=2.85e-07 
M4 VSS A0 2 VPW nch L=4e-08 W=2.85e-07 
M5 2 A1 VSS VPW nch L=4e-08 W=2.85e-07 
M6 3 B1 2 VPW nch L=4e-08 W=2.85e-07 
M7 2 B0 3 VPW nch L=4e-08 W=2.85e-07 
M8 3 B0 2 VPW nch L=4e-08 W=2.85e-07 
M9 2 B1 3 VPW nch L=4e-08 W=2.85e-07 
M10 3 B1 2 VPW nch L=4e-08 W=2.85e-07 
M11 2 B0 3 VPW nch L=4e-08 W=2.85e-07 
M12 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M13 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M16 10 A1 VDD VNW pch L=4e-08 W=3.6e-07 
M17 3 A0 10 VNW pch L=4e-08 W=3.6e-07 
M18 11 A0 3 VNW pch L=4e-08 W=3.6e-07 
M19 VDD A1 11 VNW pch L=4e-08 W=3.6e-07 
M20 12 A1 VDD VNW pch L=4e-08 W=3.6e-07 
M21 3 A0 12 VNW pch L=4e-08 W=3.6e-07 
M22 13 A0 3 VNW pch L=4e-08 W=3.6e-07 
M23 VDD A1 13 VNW pch L=4e-08 W=3.6e-07 
M24 14 B1 VDD VNW pch L=4e-08 W=3.6e-07 
M25 3 B0 14 VNW pch L=4e-08 W=3.6e-07 
M26 15 B0 3 VNW pch L=4e-08 W=3.6e-07 
M27 VDD B1 15 VNW pch L=4e-08 W=3.6e-07 
M28 16 B1 VDD VNW pch L=4e-08 W=3.6e-07 
M29 3 B0 16 VNW pch L=4e-08 W=3.6e-07 
M30 17 B0 3 VNW pch L=4e-08 W=3.6e-07 
M31 VDD B1 17 VNW pch L=4e-08 W=3.6e-07 
M32 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M33 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M34 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA22_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A0 2 VPW nch L=4e-08 W=2.6e-07 
M1 2 A1 VSS VPW nch L=4e-08 W=2.6e-07 
M2 VSS A1 2 VPW nch L=4e-08 W=2.6e-07 
M3 2 A0 VSS VPW nch L=4e-08 W=2.6e-07 
M4 VSS A0 2 VPW nch L=4e-08 W=2.6e-07 
M5 2 A1 VSS VPW nch L=4e-08 W=2.6e-07 
M6 VSS A1 2 VPW nch L=4e-08 W=2.6e-07 
M7 2 A0 VSS VPW nch L=4e-08 W=2.6e-07 
M8 VSS A0 2 VPW nch L=4e-08 W=2.6e-07 
M9 2 A1 VSS VPW nch L=4e-08 W=2.6e-07 
M10 3 B1 2 VPW nch L=4e-08 W=2.6e-07 
M11 2 B0 3 VPW nch L=4e-08 W=2.6e-07 
M12 3 B0 2 VPW nch L=4e-08 W=2.6e-07 
M13 2 B1 3 VPW nch L=4e-08 W=2.6e-07 
M14 3 B1 2 VPW nch L=4e-08 W=2.6e-07 
M15 2 B0 3 VPW nch L=4e-08 W=2.6e-07 
M16 3 B0 2 VPW nch L=4e-08 W=2.6e-07 
M17 2 B1 3 VPW nch L=4e-08 W=2.6e-07 
M18 3 B1 2 VPW nch L=4e-08 W=2.6e-07 
M19 2 B0 3 VPW nch L=4e-08 W=2.6e-07 
M20 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M21 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M22 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M23 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M24 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M25 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M26 10 A1 VDD VNW pch L=4e-08 W=3.55e-07 
M27 3 A0 10 VNW pch L=4e-08 W=3.55e-07 
M28 11 A0 3 VNW pch L=4e-08 W=3.55e-07 
M29 VDD A1 11 VNW pch L=4e-08 W=3.55e-07 
M30 12 A1 VDD VNW pch L=4e-08 W=3.55e-07 
M31 3 A0 12 VNW pch L=4e-08 W=3.55e-07 
M32 13 A0 3 VNW pch L=4e-08 W=3.55e-07 
M33 VDD A1 13 VNW pch L=4e-08 W=3.55e-07 
M34 14 A1 VDD VNW pch L=4e-08 W=3.55e-07 
M35 3 A0 14 VNW pch L=4e-08 W=3.55e-07 
M36 15 A0 3 VNW pch L=4e-08 W=3.55e-07 
M37 VDD A1 15 VNW pch L=4e-08 W=3.55e-07 
M38 16 B1 VDD VNW pch L=4e-08 W=3.55e-07 
M39 3 B0 16 VNW pch L=4e-08 W=3.55e-07 
M40 17 B0 3 VNW pch L=4e-08 W=3.55e-07 
M41 VDD B1 17 VNW pch L=4e-08 W=3.55e-07 
M42 18 B1 VDD VNW pch L=4e-08 W=3.55e-07 
M43 3 B0 18 VNW pch L=4e-08 W=3.55e-07 
M44 19 B0 3 VNW pch L=4e-08 W=3.55e-07 
M45 VDD B1 19 VNW pch L=4e-08 W=3.55e-07 
M46 20 B1 VDD VNW pch L=4e-08 W=3.55e-07 
M47 3 B0 20 VNW pch L=4e-08 W=3.55e-07 
M48 21 B0 3 VNW pch L=4e-08 W=3.55e-07 
M49 VDD B1 21 VNW pch L=4e-08 W=3.55e-07 
M50 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M51 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M52 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M53 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M54 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M55 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OA22_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M4 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M6 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M7 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M8 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M9 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M10 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M11 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M12 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M13 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M14 2 B1 1 VPW nch L=4e-08 W=2.4e-07 
M15 1 B0 2 VPW nch L=4e-08 W=2.4e-07 
M16 2 B0 1 VPW nch L=4e-08 W=2.4e-07 
M17 1 B1 2 VPW nch L=4e-08 W=2.4e-07 
M18 2 B1 1 VPW nch L=4e-08 W=2.4e-07 
M19 1 B0 2 VPW nch L=4e-08 W=2.4e-07 
M20 2 B0 1 VPW nch L=4e-08 W=2.4e-07 
M21 1 B1 2 VPW nch L=4e-08 W=2.4e-07 
M22 2 B1 1 VPW nch L=4e-08 W=2.4e-07 
M23 1 B0 2 VPW nch L=4e-08 W=2.4e-07 
M24 2 B0 1 VPW nch L=4e-08 W=2.4e-07 
M25 1 B1 2 VPW nch L=4e-08 W=2.4e-07 
M26 2 B1 1 VPW nch L=4e-08 W=2.4e-07 
M27 1 B0 2 VPW nch L=4e-08 W=2.4e-07 
M28 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M29 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M30 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M31 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M32 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M33 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M34 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M35 VSS 2 Y VPW nch L=4e-08 W=3.1e-07 
M36 10 A0 2 VNW pch L=4e-08 W=4e-07 
M37 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M38 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M39 2 A0 11 VNW pch L=4e-08 W=4e-07 
M40 12 A0 2 VNW pch L=4e-08 W=4e-07 
M41 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M42 13 A1 VDD VNW pch L=4e-08 W=4e-07 
M43 2 A0 13 VNW pch L=4e-08 W=4e-07 
M44 14 A0 2 VNW pch L=4e-08 W=4e-07 
M45 VDD A1 14 VNW pch L=4e-08 W=4e-07 
M46 15 A1 VDD VNW pch L=4e-08 W=4e-07 
M47 2 A0 15 VNW pch L=4e-08 W=4e-07 
M48 16 A0 2 VNW pch L=4e-08 W=4e-07 
M49 VDD A1 16 VNW pch L=4e-08 W=4e-07 
M50 17 B1 VDD VNW pch L=4e-08 W=4e-07 
M51 2 B0 17 VNW pch L=4e-08 W=4e-07 
M52 18 B0 2 VNW pch L=4e-08 W=4e-07 
M53 VDD B1 18 VNW pch L=4e-08 W=4e-07 
M54 19 B1 VDD VNW pch L=4e-08 W=4e-07 
M55 2 B0 19 VNW pch L=4e-08 W=4e-07 
M56 20 B0 2 VNW pch L=4e-08 W=4e-07 
M57 VDD B1 20 VNW pch L=4e-08 W=4e-07 
M58 21 B1 VDD VNW pch L=4e-08 W=4e-07 
M59 2 B0 21 VNW pch L=4e-08 W=4e-07 
M60 22 B0 2 VNW pch L=4e-08 W=4e-07 
M61 VDD B1 22 VNW pch L=4e-08 W=4e-07 
M62 23 B1 VDD VNW pch L=4e-08 W=4e-07 
M63 2 B0 23 VNW pch L=4e-08 W=4e-07 
M64 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M65 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M66 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M67 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M68 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M69 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M70 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M71 VDD 2 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI211_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=1.8e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=1.8e-07 
M2 10 B0 1 VPW nch L=4e-08 W=1.8e-07 
M3 Y C0 10 VPW nch L=4e-08 W=1.8e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=2.3e-07 
M5 Y A0 9 VNW pch L=4e-08 W=2.3e-07 
M6 VDD B0 Y VNW pch L=4e-08 W=1.2e-07 
M7 Y C0 VDD VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT OAI211_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=2.2e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.2e-07 
M2 10 B0 1 VPW nch L=4e-08 W=2.2e-07 
M3 Y C0 10 VPW nch L=4e-08 W=2.2e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M5 Y A0 9 VNW pch L=4e-08 W=2.85e-07 
M6 VDD B0 Y VNW pch L=4e-08 W=1.5e-07 
M7 Y C0 VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT OAI211_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 10 B0 1 VPW nch L=4e-08 W=3.1e-07 
M3 Y C0 10 VPW nch L=4e-08 W=3.1e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M5 Y A0 9 VNW pch L=4e-08 W=4e-07 
M6 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
M7 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI211_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=2.2e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.2e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.2e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.2e-07 
M4 11 B0 1 VPW nch L=4e-08 W=2.2e-07 
M5 Y C0 11 VPW nch L=4e-08 W=2.2e-07 
M6 12 C0 Y VPW nch L=4e-08 W=2.2e-07 
M7 1 B0 12 VPW nch L=4e-08 W=2.2e-07 
M8 9 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M9 Y A0 9 VNW pch L=4e-08 W=2.85e-07 
M10 10 A0 Y VNW pch L=4e-08 W=2.85e-07 
M11 VDD A1 10 VNW pch L=4e-08 W=2.85e-07 
M12 Y B0 VDD VNW pch L=4e-08 W=1.5e-07 
M13 VDD C0 Y VNW pch L=4e-08 W=1.5e-07 
M14 Y C0 VDD VNW pch L=4e-08 W=1.5e-07 
M15 VDD B0 Y VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT OAI211_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 11 B0 1 VPW nch L=4e-08 W=3.1e-07 
M5 Y C0 11 VPW nch L=4e-08 W=3.1e-07 
M6 12 C0 Y VPW nch L=4e-08 W=3.1e-07 
M7 1 B0 12 VPW nch L=4e-08 W=3.1e-07 
M8 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M9 Y A0 9 VNW pch L=4e-08 W=4e-07 
M10 10 A0 Y VNW pch L=4e-08 W=4e-07 
M11 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M12 Y B0 VDD VNW pch L=4e-08 W=2.1e-07 
M13 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
M14 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
M15 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI211_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 12 B0 1 VPW nch L=4e-08 W=3.1e-07 
M7 Y C0 12 VPW nch L=4e-08 W=3.1e-07 
M8 13 C0 Y VPW nch L=4e-08 W=3.1e-07 
M9 1 B0 13 VPW nch L=4e-08 W=3.1e-07 
M10 14 B0 1 VPW nch L=4e-08 W=3.1e-07 
M11 Y C0 14 VPW nch L=4e-08 W=3.1e-07 
M12 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y A0 9 VNW pch L=4e-08 W=4e-07 
M14 10 A0 Y VNW pch L=4e-08 W=4e-07 
M15 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M16 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M17 Y A0 11 VNW pch L=4e-08 W=4e-07 
M18 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
M19 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
M20 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
M21 Y B0 VDD VNW pch L=4e-08 W=2.1e-07 
M22 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
M23 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI211_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M8 13 B0 1 VPW nch L=4e-08 W=3.1e-07 
M9 Y C0 13 VPW nch L=4e-08 W=3.1e-07 
M10 14 C0 Y VPW nch L=4e-08 W=3.1e-07 
M11 1 B0 14 VPW nch L=4e-08 W=3.1e-07 
M12 15 B0 1 VPW nch L=4e-08 W=3.1e-07 
M13 Y C0 15 VPW nch L=4e-08 W=3.1e-07 
M14 16 C0 Y VPW nch L=4e-08 W=3.1e-07 
M15 1 B0 16 VPW nch L=4e-08 W=3.1e-07 
M16 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M17 Y A0 9 VNW pch L=4e-08 W=4e-07 
M18 10 A0 Y VNW pch L=4e-08 W=4e-07 
M19 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M20 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M21 Y A0 11 VNW pch L=4e-08 W=4e-07 
M22 12 A0 Y VNW pch L=4e-08 W=4e-07 
M23 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M24 Y B0 VDD VNW pch L=4e-08 W=2.1e-07 
M25 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
M26 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
M27 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
M28 Y B0 VDD VNW pch L=4e-08 W=2.1e-07 
M29 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
M30 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
M31 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI21B_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 VSS B0N 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A1 4 VPW nch L=4e-08 W=1.4e-07 
M2 4 A0 VSS VPW nch L=4e-08 W=1.4e-07 
M3 Y 1 4 VPW nch L=4e-08 W=1.4e-07 
M4 VDD B0N 1 VNW pch L=4e-08 W=1.55e-07 
M5 9 A1 VDD VNW pch L=4e-08 W=2.3e-07 
M6 Y A0 9 VNW pch L=4e-08 W=2.3e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT OAI21B_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 VSS B0N 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A1 4 VPW nch L=4e-08 W=1.7e-07 
M2 4 A0 VSS VPW nch L=4e-08 W=1.7e-07 
M3 Y 1 4 VPW nch L=4e-08 W=1.7e-07 
M4 VDD B0N 1 VNW pch L=4e-08 W=1.55e-07 
M5 9 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M6 Y A0 9 VNW pch L=4e-08 W=2.85e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT OAI21B_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 VSS B0N 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS A1 4 VPW nch L=4e-08 W=2.4e-07 
M2 4 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y 1 4 VPW nch L=4e-08 W=2.4e-07 
M4 VDD B0N 1 VNW pch L=4e-08 W=1.55e-07 
M5 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M6 Y A0 9 VNW pch L=4e-08 W=4e-07 
M7 VDD 1 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI21B_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 VSS A0 2 VPW nch L=4e-08 W=3.4e-07 
M1 2 A1 VSS VPW nch L=4e-08 W=3.4e-07 
M2 Y 5 2 VPW nch L=4e-08 W=3.4e-07 
M3 VSS B0N 5 VPW nch L=4e-08 W=1.2e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M5 Y A0 9 VNW pch L=4e-08 W=2.85e-07 
M6 10 A0 Y VNW pch L=4e-08 W=2.85e-07 
M7 VDD A1 10 VNW pch L=4e-08 W=2.85e-07 
M8 Y 5 VDD VNW pch L=4e-08 W=3e-07 
M9 VDD B0N 5 VNW pch L=4e-08 W=1.55e-07 
.ENDS


.SUBCKT OAI21B_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M4 Y 5 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 5 Y VPW nch L=4e-08 W=2.4e-07 
M6 VSS B0N 5 VPW nch L=4e-08 W=1.2e-07 
M7 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M8 Y A0 9 VNW pch L=4e-08 W=4e-07 
M9 10 A0 Y VNW pch L=4e-08 W=4e-07 
M10 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M11 Y 5 VDD VNW pch L=4e-08 W=2.1e-07 
M12 VDD 5 Y VNW pch L=4e-08 W=2.1e-07 
M13 VDD B0N 5 VNW pch L=4e-08 W=1.55e-07 
.ENDS


.SUBCKT OAI21B_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 VSS A1 2 VPW nch L=4e-08 W=3.6e-07 
M1 2 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M2 VSS A0 2 VPW nch L=4e-08 W=3.6e-07 
M3 2 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M4 Y 5 2 VPW nch L=4e-08 W=3.6e-07 
M5 2 5 Y VPW nch L=4e-08 W=3.6e-07 
M6 5 B0N VSS VPW nch L=4e-08 W=1.75e-07 
M7 9 A0 Y VNW pch L=4e-08 W=4e-07 
M8 VDD A1 9 VNW pch L=4e-08 W=4e-07 
M9 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M10 Y A0 10 VNW pch L=4e-08 W=4e-07 
M11 11 A0 Y VNW pch L=4e-08 W=4e-07 
M12 VDD A1 11 VNW pch L=4e-08 W=4e-07 
M13 Y 5 VDD VNW pch L=4e-08 W=3.15e-07 
M14 VDD 5 Y VNW pch L=4e-08 W=3.15e-07 
M15 5 B0N VDD VNW pch L=4e-08 W=2.3e-07 
.ENDS


.SUBCKT OAI21B_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M6 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M7 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M8 Y 5 1 VPW nch L=4e-08 W=3.2e-07 
M9 1 5 Y VPW nch L=4e-08 W=3.2e-07 
M10 Y 5 1 VPW nch L=4e-08 W=3.2e-07 
M11 5 B0N VSS VPW nch L=4e-08 W=2.35e-07 
M12 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y A0 9 VNW pch L=4e-08 W=4e-07 
M14 10 A0 Y VNW pch L=4e-08 W=4e-07 
M15 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M16 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M17 Y A0 11 VNW pch L=4e-08 W=4e-07 
M18 12 A0 Y VNW pch L=4e-08 W=4e-07 
M19 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M20 Y 5 VDD VNW pch L=4e-08 W=2.8e-07 
M21 VDD 5 Y VNW pch L=4e-08 W=2.8e-07 
M22 Y 5 VDD VNW pch L=4e-08 W=2.8e-07 
M23 5 B0N VDD VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT OAI21B_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M6 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M7 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M8 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M9 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M10 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M11 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M12 Y 5 1 VPW nch L=4e-08 W=3.6e-07 
M13 1 5 Y VPW nch L=4e-08 W=3.6e-07 
M14 Y 5 1 VPW nch L=4e-08 W=3.6e-07 
M15 1 5 Y VPW nch L=4e-08 W=3.6e-07 
M16 5 B0N VSS VPW nch L=4e-08 W=3.5e-07 
M17 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M18 Y A0 9 VNW pch L=4e-08 W=4e-07 
M19 10 A0 Y VNW pch L=4e-08 W=4e-07 
M20 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M21 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M22 Y A0 11 VNW pch L=4e-08 W=4e-07 
M23 12 A0 Y VNW pch L=4e-08 W=4e-07 
M24 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M25 13 A1 VDD VNW pch L=4e-08 W=4e-07 
M26 Y A0 13 VNW pch L=4e-08 W=4e-07 
M27 14 A0 Y VNW pch L=4e-08 W=4e-07 
M28 VDD A1 14 VNW pch L=4e-08 W=4e-07 
M29 Y 5 VDD VNW pch L=4e-08 W=3.15e-07 
M30 VDD 5 Y VNW pch L=4e-08 W=3.15e-07 
M31 Y 5 VDD VNW pch L=4e-08 W=3.15e-07 
M32 VDD 5 Y VNW pch L=4e-08 W=3.15e-07 
M33 5 B0N VDD VNW pch L=4e-08 W=2.25e-07 
M34 VDD B0N 5 VNW pch L=4e-08 W=2.25e-07 
.ENDS


.SUBCKT OAI21B_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0N
M0 VSS A0 3 VPW nch L=4e-08 W=3.85e-07 
M1 3 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M2 VSS A1 3 VPW nch L=4e-08 W=3.85e-07 
M3 3 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M4 VSS A0 3 VPW nch L=4e-08 W=3.85e-07 
M5 3 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M6 VSS A1 3 VPW nch L=4e-08 W=3.85e-07 
M7 3 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M8 VSS A0 3 VPW nch L=4e-08 W=3.85e-07 
M9 3 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M10 Y 5 3 VPW nch L=4e-08 W=3.85e-07 
M11 3 5 Y VPW nch L=4e-08 W=3.85e-07 
M12 Y 5 3 VPW nch L=4e-08 W=3.85e-07 
M13 3 5 Y VPW nch L=4e-08 W=3.85e-07 
M14 Y 5 3 VPW nch L=4e-08 W=3.85e-07 
M15 5 B0N VSS VPW nch L=4e-08 W=2.3e-07 
M16 VSS B0N 5 VPW nch L=4e-08 W=2.3e-07 
M17 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M18 Y A0 9 VNW pch L=4e-08 W=4e-07 
M19 10 A0 Y VNW pch L=4e-08 W=4e-07 
M20 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M21 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M22 Y A0 11 VNW pch L=4e-08 W=4e-07 
M23 12 A0 Y VNW pch L=4e-08 W=4e-07 
M24 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M25 13 A1 VDD VNW pch L=4e-08 W=4e-07 
M26 Y A0 13 VNW pch L=4e-08 W=4e-07 
M27 14 A0 Y VNW pch L=4e-08 W=4e-07 
M28 VDD A1 14 VNW pch L=4e-08 W=4e-07 
M29 15 A1 VDD VNW pch L=4e-08 W=4e-07 
M30 Y A0 15 VNW pch L=4e-08 W=4e-07 
M31 16 A0 Y VNW pch L=4e-08 W=4e-07 
M32 VDD A1 16 VNW pch L=4e-08 W=4e-07 
M33 Y 5 VDD VNW pch L=4e-08 W=3.35e-07 
M34 VDD 5 Y VNW pch L=4e-08 W=3.35e-07 
M35 Y 5 VDD VNW pch L=4e-08 W=3.35e-07 
M36 VDD 5 Y VNW pch L=4e-08 W=3.35e-07 
M37 Y 5 VDD VNW pch L=4e-08 W=3.35e-07 
M38 5 B0N VDD VNW pch L=4e-08 W=3e-07 
M39 VDD B0N 5 VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT OAI21_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=1.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=1.4e-07 
M2 Y B0 1 VPW nch L=4e-08 W=1.4e-07 
M3 8 A1 VDD VNW pch L=4e-08 W=2.3e-07 
M4 Y A0 8 VNW pch L=4e-08 W=2.3e-07 
M5 VDD B0 Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT OAI21_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=1.7e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=1.7e-07 
M2 Y B0 1 VPW nch L=4e-08 W=1.7e-07 
M3 8 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M4 Y A0 8 VNW pch L=4e-08 W=2.85e-07 
M5 VDD B0 Y VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT OAI21_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 Y B0 1 VPW nch L=4e-08 W=2.4e-07 
M3 8 A1 VDD VNW pch L=4e-08 W=4e-07 
M4 Y A0 8 VNW pch L=4e-08 W=4e-07 
M5 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI21_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A0 2 VPW nch L=4e-08 W=4e-07 
M1 2 A1 VSS VPW nch L=4e-08 W=4e-07 
M2 Y B0 2 VPW nch L=4e-08 W=4e-07 
M3 8 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M4 Y A0 8 VNW pch L=4e-08 W=2.85e-07 
M5 9 A0 Y VNW pch L=4e-08 W=2.85e-07 
M6 VDD A1 9 VNW pch L=4e-08 W=2.85e-07 
M7 Y B0 VDD VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT OAI21_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M4 Y B0 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 B0 Y VPW nch L=4e-08 W=2.4e-07 
M6 8 A1 VDD VNW pch L=4e-08 W=4e-07 
M7 Y A0 8 VNW pch L=4e-08 W=4e-07 
M8 9 A0 Y VNW pch L=4e-08 W=4e-07 
M9 VDD A1 9 VNW pch L=4e-08 W=4e-07 
M10 Y B0 VDD VNW pch L=4e-08 W=2.1e-07 
M11 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI21_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M6 Y B0 1 VPW nch L=4e-08 W=3.6e-07 
M7 1 B0 Y VPW nch L=4e-08 W=3.6e-07 
M8 8 A1 VDD VNW pch L=4e-08 W=4e-07 
M9 Y A0 8 VNW pch L=4e-08 W=4e-07 
M10 9 A0 Y VNW pch L=4e-08 W=4e-07 
M11 VDD A1 9 VNW pch L=4e-08 W=4e-07 
M12 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y A0 10 VNW pch L=4e-08 W=4e-07 
M14 VDD B0 Y VNW pch L=4e-08 W=3.15e-07 
M15 Y B0 VDD VNW pch L=4e-08 W=3.15e-07 
.ENDS


.SUBCKT OAI21_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M6 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M7 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M8 Y B0 1 VPW nch L=4e-08 W=3.2e-07 
M9 1 B0 Y VPW nch L=4e-08 W=3.2e-07 
M10 Y B0 1 VPW nch L=4e-08 W=3.2e-07 
M11 8 A1 VDD VNW pch L=4e-08 W=4e-07 
M12 Y A0 8 VNW pch L=4e-08 W=4e-07 
M13 9 A0 Y VNW pch L=4e-08 W=4e-07 
M14 VDD A1 9 VNW pch L=4e-08 W=4e-07 
M15 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M16 Y A0 10 VNW pch L=4e-08 W=4e-07 
M17 11 A0 Y VNW pch L=4e-08 W=4e-07 
M18 VDD A1 11 VNW pch L=4e-08 W=4e-07 
M19 Y B0 VDD VNW pch L=4e-08 W=2.8e-07 
M20 VDD B0 Y VNW pch L=4e-08 W=2.8e-07 
M21 Y B0 VDD VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT OAI21_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M6 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M7 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M8 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M9 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M10 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M11 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M12 Y B0 1 VPW nch L=4e-08 W=3.6e-07 
M13 1 B0 Y VPW nch L=4e-08 W=3.6e-07 
M14 Y B0 1 VPW nch L=4e-08 W=3.6e-07 
M15 1 B0 Y VPW nch L=4e-08 W=3.6e-07 
M16 8 A1 VDD VNW pch L=4e-08 W=4e-07 
M17 Y A0 8 VNW pch L=4e-08 W=4e-07 
M18 9 A0 Y VNW pch L=4e-08 W=4e-07 
M19 VDD A1 9 VNW pch L=4e-08 W=4e-07 
M20 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M21 Y A0 10 VNW pch L=4e-08 W=4e-07 
M22 11 A0 Y VNW pch L=4e-08 W=4e-07 
M23 VDD A1 11 VNW pch L=4e-08 W=4e-07 
M24 12 A1 VDD VNW pch L=4e-08 W=4e-07 
M25 Y A0 12 VNW pch L=4e-08 W=4e-07 
M26 13 A0 Y VNW pch L=4e-08 W=4e-07 
M27 VDD A1 13 VNW pch L=4e-08 W=4e-07 
M28 Y B0 VDD VNW pch L=4e-08 W=3.15e-07 
M29 VDD B0 Y VNW pch L=4e-08 W=3.15e-07 
M30 Y B0 VDD VNW pch L=4e-08 W=3.15e-07 
M31 VDD B0 Y VNW pch L=4e-08 W=3.15e-07 
.ENDS


.SUBCKT OAI21_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0
M0 VSS A0 3 VPW nch L=4e-08 W=3.85e-07 
M1 3 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M2 VSS A1 3 VPW nch L=4e-08 W=3.85e-07 
M3 3 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M4 VSS A0 3 VPW nch L=4e-08 W=3.85e-07 
M5 3 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M6 VSS A1 3 VPW nch L=4e-08 W=3.85e-07 
M7 3 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M8 VSS A0 3 VPW nch L=4e-08 W=3.85e-07 
M9 3 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M10 Y B0 3 VPW nch L=4e-08 W=3.85e-07 
M11 3 B0 Y VPW nch L=4e-08 W=3.85e-07 
M12 Y B0 3 VPW nch L=4e-08 W=3.85e-07 
M13 3 B0 Y VPW nch L=4e-08 W=3.85e-07 
M14 Y B0 3 VPW nch L=4e-08 W=3.85e-07 
M15 8 A1 VDD VNW pch L=4e-08 W=4e-07 
M16 Y A0 8 VNW pch L=4e-08 W=4e-07 
M17 9 A0 Y VNW pch L=4e-08 W=4e-07 
M18 VDD A1 9 VNW pch L=4e-08 W=4e-07 
M19 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M20 Y A0 10 VNW pch L=4e-08 W=4e-07 
M21 11 A0 Y VNW pch L=4e-08 W=4e-07 
M22 VDD A1 11 VNW pch L=4e-08 W=4e-07 
M23 12 A1 VDD VNW pch L=4e-08 W=4e-07 
M24 Y A0 12 VNW pch L=4e-08 W=4e-07 
M25 13 A0 Y VNW pch L=4e-08 W=4e-07 
M26 VDD A1 13 VNW pch L=4e-08 W=4e-07 
M27 14 A1 VDD VNW pch L=4e-08 W=4e-07 
M28 Y A0 14 VNW pch L=4e-08 W=4e-07 
M29 15 A0 Y VNW pch L=4e-08 W=4e-07 
M30 VDD A1 15 VNW pch L=4e-08 W=4e-07 
M31 Y B0 VDD VNW pch L=4e-08 W=3.35e-07 
M32 VDD B0 Y VNW pch L=4e-08 W=3.35e-07 
M33 Y B0 VDD VNW pch L=4e-08 W=3.35e-07 
M34 VDD B0 Y VNW pch L=4e-08 W=3.35e-07 
M35 Y B0 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT OAI221_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 VSS A1 1 VPW nch L=4e-08 W=2.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.1e-07 
M2 5 B0 1 VPW nch L=4e-08 W=2.1e-07 
M3 1 B1 5 VPW nch L=4e-08 W=2.1e-07 
M4 Y C0 5 VPW nch L=4e-08 W=2.1e-07 
M5 11 A1 VDD VNW pch L=4e-08 W=2.3e-07 
M6 Y A0 11 VNW pch L=4e-08 W=2.3e-07 
M7 12 B0 Y VNW pch L=4e-08 W=2.3e-07 
M8 VDD B1 12 VNW pch L=4e-08 W=2.3e-07 
M9 Y C0 VDD VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT OAI221_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 VSS A1 1 VPW nch L=4e-08 W=2.2e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.2e-07 
M2 5 B0 1 VPW nch L=4e-08 W=2.2e-07 
M3 1 B1 5 VPW nch L=4e-08 W=2.2e-07 
M4 Y C0 5 VPW nch L=4e-08 W=2.2e-07 
M5 11 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M6 Y A0 11 VNW pch L=4e-08 W=2.85e-07 
M7 12 B0 Y VNW pch L=4e-08 W=2.85e-07 
M8 VDD B1 12 VNW pch L=4e-08 W=2.85e-07 
M9 Y C0 VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT OAI221_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M4 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M5 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M6 Y A0 11 VNW pch L=4e-08 W=4e-07 
M7 12 B0 Y VNW pch L=4e-08 W=4e-07 
M8 VDD B1 12 VNW pch L=4e-08 W=4e-07 
M9 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI221_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 VSS A1 1 VPW nch L=4e-08 W=2.2e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.2e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.2e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.2e-07 
M4 5 B1 1 VPW nch L=4e-08 W=2.2e-07 
M5 1 B0 5 VPW nch L=4e-08 W=2.2e-07 
M6 5 B0 1 VPW nch L=4e-08 W=2.2e-07 
M7 1 B1 5 VPW nch L=4e-08 W=2.2e-07 
M8 Y C0 5 VPW nch L=4e-08 W=2.2e-07 
M9 5 C0 Y VPW nch L=4e-08 W=2.2e-07 
M10 11 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M11 Y A0 11 VNW pch L=4e-08 W=2.85e-07 
M12 12 A0 Y VNW pch L=4e-08 W=2.85e-07 
M13 VDD A1 12 VNW pch L=4e-08 W=2.85e-07 
M14 13 B1 VDD VNW pch L=4e-08 W=2.85e-07 
M15 Y B0 13 VNW pch L=4e-08 W=2.85e-07 
M16 14 B0 Y VNW pch L=4e-08 W=2.85e-07 
M17 VDD B1 14 VNW pch L=4e-08 W=2.85e-07 
M18 Y C0 VDD VNW pch L=4e-08 W=1.5e-07 
M19 VDD C0 Y VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT OAI221_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 5 B1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 B0 5 VPW nch L=4e-08 W=3.1e-07 
M6 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M8 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M9 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M10 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M11 Y A0 11 VNW pch L=4e-08 W=4e-07 
M12 12 A0 Y VNW pch L=4e-08 W=4e-07 
M13 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M14 13 B1 VDD VNW pch L=4e-08 W=4e-07 
M15 Y B0 13 VNW pch L=4e-08 W=4e-07 
M16 14 B0 Y VNW pch L=4e-08 W=4e-07 
M17 VDD B1 14 VNW pch L=4e-08 W=4e-07 
M18 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
M19 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI221_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M8 5 B1 1 VPW nch L=4e-08 W=3.1e-07 
M9 1 B0 5 VPW nch L=4e-08 W=3.1e-07 
M10 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M11 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M12 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M13 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M14 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M15 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M16 Y A0 11 VNW pch L=4e-08 W=4e-07 
M17 12 A0 Y VNW pch L=4e-08 W=4e-07 
M18 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M19 13 A1 VDD VNW pch L=4e-08 W=4e-07 
M20 Y A0 13 VNW pch L=4e-08 W=4e-07 
M21 14 B0 Y VNW pch L=4e-08 W=4e-07 
M22 VDD B1 14 VNW pch L=4e-08 W=4e-07 
M23 15 B1 VDD VNW pch L=4e-08 W=4e-07 
M24 Y B0 15 VNW pch L=4e-08 W=4e-07 
M25 16 B0 Y VNW pch L=4e-08 W=4e-07 
M26 VDD B1 16 VNW pch L=4e-08 W=4e-07 
M27 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
M28 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
M29 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI221_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M8 5 B1 1 VPW nch L=4e-08 W=3.1e-07 
M9 1 B0 5 VPW nch L=4e-08 W=3.1e-07 
M10 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M11 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M12 5 B1 1 VPW nch L=4e-08 W=3.1e-07 
M13 1 B0 5 VPW nch L=4e-08 W=3.1e-07 
M14 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M15 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M16 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M17 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M18 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M19 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M20 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M21 Y A0 11 VNW pch L=4e-08 W=4e-07 
M22 12 A0 Y VNW pch L=4e-08 W=4e-07 
M23 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M24 13 A1 VDD VNW pch L=4e-08 W=4e-07 
M25 Y A0 13 VNW pch L=4e-08 W=4e-07 
M26 14 A0 Y VNW pch L=4e-08 W=4e-07 
M27 VDD A1 14 VNW pch L=4e-08 W=4e-07 
M28 15 B1 VDD VNW pch L=4e-08 W=4e-07 
M29 Y B0 15 VNW pch L=4e-08 W=4e-07 
M30 16 B0 Y VNW pch L=4e-08 W=4e-07 
M31 VDD B1 16 VNW pch L=4e-08 W=4e-07 
M32 17 B1 VDD VNW pch L=4e-08 W=4e-07 
M33 Y B0 17 VNW pch L=4e-08 W=4e-07 
M34 18 B0 Y VNW pch L=4e-08 W=4e-07 
M35 VDD B1 18 VNW pch L=4e-08 W=4e-07 
M36 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
M37 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
M38 Y C0 VDD VNW pch L=4e-08 W=2.1e-07 
M39 VDD C0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI222_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 VSS A1 1 VPW nch L=4e-08 W=2.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.1e-07 
M2 5 B0 1 VPW nch L=4e-08 W=2.1e-07 
M3 1 B1 5 VPW nch L=4e-08 W=2.1e-07 
M4 Y C1 5 VPW nch L=4e-08 W=2.1e-07 
M5 5 C0 Y VPW nch L=4e-08 W=2.1e-07 
M6 12 A1 VDD VNW pch L=4e-08 W=2e-07 
M7 Y A0 12 VNW pch L=4e-08 W=2e-07 
M8 13 B0 Y VNW pch L=4e-08 W=2e-07 
M9 VDD B1 13 VNW pch L=4e-08 W=2e-07 
M10 14 C1 VDD VNW pch L=4e-08 W=2e-07 
M11 Y C0 14 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OAI222_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 VSS A1 1 VPW nch L=4e-08 W=2.2e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.2e-07 
M2 5 B0 1 VPW nch L=4e-08 W=2.2e-07 
M3 1 B1 5 VPW nch L=4e-08 W=2.2e-07 
M4 Y C1 5 VPW nch L=4e-08 W=2.2e-07 
M5 5 C0 Y VPW nch L=4e-08 W=2.2e-07 
M6 12 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M7 Y A0 12 VNW pch L=4e-08 W=2.85e-07 
M8 13 B0 Y VNW pch L=4e-08 W=2.85e-07 
M9 VDD B1 13 VNW pch L=4e-08 W=2.85e-07 
M10 14 C1 VDD VNW pch L=4e-08 W=2.85e-07 
M11 Y C0 14 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OAI222_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M4 Y C1 5 VPW nch L=4e-08 W=3.1e-07 
M5 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M6 12 A1 VDD VNW pch L=4e-08 W=4e-07 
M7 Y A0 12 VNW pch L=4e-08 W=4e-07 
M8 13 B0 Y VNW pch L=4e-08 W=4e-07 
M9 VDD B1 13 VNW pch L=4e-08 W=4e-07 
M10 14 C1 VDD VNW pch L=4e-08 W=4e-07 
M11 Y C0 14 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI222_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 VSS A1 1 VPW nch L=4e-08 W=2.2e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.2e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.2e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.2e-07 
M4 5 B1 1 VPW nch L=4e-08 W=2.2e-07 
M5 1 B0 5 VPW nch L=4e-08 W=2.2e-07 
M6 5 B0 1 VPW nch L=4e-08 W=2.2e-07 
M7 1 B1 5 VPW nch L=4e-08 W=2.2e-07 
M8 Y C1 5 VPW nch L=4e-08 W=2.2e-07 
M9 5 C0 Y VPW nch L=4e-08 W=2.2e-07 
M10 Y C0 5 VPW nch L=4e-08 W=2.2e-07 
M11 5 C1 Y VPW nch L=4e-08 W=2.2e-07 
M12 12 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M13 Y A0 12 VNW pch L=4e-08 W=2.85e-07 
M14 13 A0 Y VNW pch L=4e-08 W=2.85e-07 
M15 VDD A1 13 VNW pch L=4e-08 W=2.85e-07 
M16 14 B1 VDD VNW pch L=4e-08 W=2.85e-07 
M17 Y B0 14 VNW pch L=4e-08 W=2.85e-07 
M18 15 B0 Y VNW pch L=4e-08 W=2.85e-07 
M19 VDD B1 15 VNW pch L=4e-08 W=2.85e-07 
M20 16 C1 VDD VNW pch L=4e-08 W=2.85e-07 
M21 Y C0 16 VNW pch L=4e-08 W=2.85e-07 
M22 17 C0 Y VNW pch L=4e-08 W=2.85e-07 
M23 VDD C1 17 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OAI222_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 5 B1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 B0 5 VPW nch L=4e-08 W=3.1e-07 
M6 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M8 Y C1 5 VPW nch L=4e-08 W=3.1e-07 
M9 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M10 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M11 5 C1 Y VPW nch L=4e-08 W=3.1e-07 
M12 12 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y A0 12 VNW pch L=4e-08 W=4e-07 
M14 13 A0 Y VNW pch L=4e-08 W=4e-07 
M15 VDD A1 13 VNW pch L=4e-08 W=4e-07 
M16 14 B1 VDD VNW pch L=4e-08 W=4e-07 
M17 Y B0 14 VNW pch L=4e-08 W=4e-07 
M18 15 B0 Y VNW pch L=4e-08 W=4e-07 
M19 VDD B1 15 VNW pch L=4e-08 W=4e-07 
M20 16 C1 VDD VNW pch L=4e-08 W=4e-07 
M21 Y C0 16 VNW pch L=4e-08 W=4e-07 
M22 17 C0 Y VNW pch L=4e-08 W=4e-07 
M23 VDD C1 17 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI222_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M8 5 B1 1 VPW nch L=4e-08 W=3.1e-07 
M9 1 B0 5 VPW nch L=4e-08 W=3.1e-07 
M10 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M11 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M12 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M13 5 C1 Y VPW nch L=4e-08 W=3.1e-07 
M14 Y C1 5 VPW nch L=4e-08 W=3.1e-07 
M15 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M16 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M17 5 C1 Y VPW nch L=4e-08 W=3.1e-07 
M18 12 A1 VDD VNW pch L=4e-08 W=4e-07 
M19 Y A0 12 VNW pch L=4e-08 W=4e-07 
M20 13 A0 Y VNW pch L=4e-08 W=4e-07 
M21 VDD A1 13 VNW pch L=4e-08 W=4e-07 
M22 14 A1 VDD VNW pch L=4e-08 W=4e-07 
M23 Y A0 14 VNW pch L=4e-08 W=4e-07 
M24 15 B0 Y VNW pch L=4e-08 W=4e-07 
M25 VDD B1 15 VNW pch L=4e-08 W=4e-07 
M26 16 B1 VDD VNW pch L=4e-08 W=4e-07 
M27 Y B0 16 VNW pch L=4e-08 W=4e-07 
M28 17 B0 Y VNW pch L=4e-08 W=4e-07 
M29 VDD B1 17 VNW pch L=4e-08 W=4e-07 
M30 18 C0 Y VNW pch L=4e-08 W=4e-07 
M31 VDD C1 18 VNW pch L=4e-08 W=4e-07 
M32 19 C1 VDD VNW pch L=4e-08 W=4e-07 
M33 Y C0 19 VNW pch L=4e-08 W=4e-07 
M34 20 C0 Y VNW pch L=4e-08 W=4e-07 
M35 VDD C1 20 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI222_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
M0 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS A1 1 VPW nch L=4e-08 W=3.1e-07 
M5 1 A0 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VSS A0 1 VPW nch L=4e-08 W=3.1e-07 
M7 1 A1 VSS VPW nch L=4e-08 W=3.1e-07 
M8 5 B1 1 VPW nch L=4e-08 W=3.1e-07 
M9 1 B0 5 VPW nch L=4e-08 W=3.1e-07 
M10 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M11 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M12 5 B1 1 VPW nch L=4e-08 W=3.1e-07 
M13 1 B0 5 VPW nch L=4e-08 W=3.1e-07 
M14 5 B0 1 VPW nch L=4e-08 W=3.1e-07 
M15 1 B1 5 VPW nch L=4e-08 W=3.1e-07 
M16 Y C1 5 VPW nch L=4e-08 W=3.1e-07 
M17 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M18 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M19 5 C1 Y VPW nch L=4e-08 W=3.1e-07 
M20 Y C1 5 VPW nch L=4e-08 W=3.1e-07 
M21 5 C0 Y VPW nch L=4e-08 W=3.1e-07 
M22 Y C0 5 VPW nch L=4e-08 W=3.1e-07 
M23 5 C1 Y VPW nch L=4e-08 W=3.1e-07 
M24 12 A1 VDD VNW pch L=4e-08 W=4e-07 
M25 Y A0 12 VNW pch L=4e-08 W=4e-07 
M26 13 A0 Y VNW pch L=4e-08 W=4e-07 
M27 VDD A1 13 VNW pch L=4e-08 W=4e-07 
M28 14 A1 VDD VNW pch L=4e-08 W=4e-07 
M29 Y A0 14 VNW pch L=4e-08 W=4e-07 
M30 15 A0 Y VNW pch L=4e-08 W=4e-07 
M31 VDD A1 15 VNW pch L=4e-08 W=4e-07 
M32 16 B1 VDD VNW pch L=4e-08 W=4e-07 
M33 Y B0 16 VNW pch L=4e-08 W=4e-07 
M34 17 B0 Y VNW pch L=4e-08 W=4e-07 
M35 VDD B1 17 VNW pch L=4e-08 W=4e-07 
M36 18 B1 VDD VNW pch L=4e-08 W=4e-07 
M37 Y B0 18 VNW pch L=4e-08 W=4e-07 
M38 19 B0 Y VNW pch L=4e-08 W=4e-07 
M39 VDD B1 19 VNW pch L=4e-08 W=4e-07 
M40 20 C1 VDD VNW pch L=4e-08 W=4e-07 
M41 Y C0 20 VNW pch L=4e-08 W=4e-07 
M42 21 C0 Y VNW pch L=4e-08 W=4e-07 
M43 VDD C1 21 VNW pch L=4e-08 W=4e-07 
M44 22 C1 VDD VNW pch L=4e-08 W=4e-07 
M45 Y C0 22 VNW pch L=4e-08 W=4e-07 
M46 23 C0 Y VNW pch L=4e-08 W=4e-07 
M47 VDD C1 23 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI22BB_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 11 B1N VSS VPW nch L=4e-08 W=1.2e-07 
M1 3 B0N 11 VPW nch L=4e-08 W=1.2e-07 
M2 VSS A1 4 VPW nch L=4e-08 W=1.4e-07 
M3 4 A0 VSS VPW nch L=4e-08 W=1.4e-07 
M4 Y 3 4 VPW nch L=4e-08 W=1.4e-07 
M5 3 B1N VDD VNW pch L=4e-08 W=1.2e-07 
M6 VDD B0N 3 VNW pch L=4e-08 W=1.2e-07 
M7 10 A1 VDD VNW pch L=4e-08 W=2.3e-07 
M8 Y A0 10 VNW pch L=4e-08 W=2.3e-07 
M9 VDD 3 Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT OAI22BB_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 11 B1N VSS VPW nch L=4e-08 W=1.3e-07 
M1 3 B0N 11 VPW nch L=4e-08 W=1.3e-07 
M2 VSS A1 4 VPW nch L=4e-08 W=1.7e-07 
M3 4 A0 VSS VPW nch L=4e-08 W=1.7e-07 
M4 Y 3 4 VPW nch L=4e-08 W=1.7e-07 
M5 3 B1N VDD VNW pch L=4e-08 W=1.2e-07 
M6 VDD B0N 3 VNW pch L=4e-08 W=1.2e-07 
M7 10 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M8 Y A0 10 VNW pch L=4e-08 W=2.85e-07 
M9 VDD 3 Y VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT OAI22BB_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 11 B1N VSS VPW nch L=4e-08 W=1.5e-07 
M1 3 B0N 11 VPW nch L=4e-08 W=1.5e-07 
M2 VSS A1 4 VPW nch L=4e-08 W=2.4e-07 
M3 4 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M4 Y 3 4 VPW nch L=4e-08 W=2.4e-07 
M5 3 B1N VDD VNW pch L=4e-08 W=1.3e-07 
M6 VDD B0N 3 VNW pch L=4e-08 W=1.3e-07 
M7 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M8 Y A0 10 VNW pch L=4e-08 W=4e-07 
M9 VDD 3 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI22BB_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 12 B1N VSS VPW nch L=4e-08 W=2e-07 
M1 3 B0N 12 VPW nch L=4e-08 W=2e-07 
M2 VSS A0 4 VPW nch L=4e-08 W=3.4e-07 
M3 4 A1 VSS VPW nch L=4e-08 W=3.4e-07 
M4 Y 3 4 VPW nch L=4e-08 W=3.4e-07 
M5 3 B1N VDD VNW pch L=4e-08 W=1.7e-07 
M6 VDD B0N 3 VNW pch L=4e-08 W=1.7e-07 
M7 10 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M8 Y A0 10 VNW pch L=4e-08 W=2.85e-07 
M9 11 A0 Y VNW pch L=4e-08 W=2.85e-07 
M10 VDD A1 11 VNW pch L=4e-08 W=2.85e-07 
M11 Y 3 VDD VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT OAI22BB_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 12 B1N VSS VPW nch L=4e-08 W=2.45e-07 
M1 3 B0N 12 VPW nch L=4e-08 W=2.45e-07 
M2 Y 3 4 VPW nch L=4e-08 W=2.4e-07 
M3 4 3 Y VPW nch L=4e-08 W=2.4e-07 
M4 VSS A1 4 VPW nch L=4e-08 W=2.4e-07 
M5 4 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M6 VSS A0 4 VPW nch L=4e-08 W=2.4e-07 
M7 4 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M8 3 B1N VDD VNW pch L=4e-08 W=2.1e-07 
M9 VDD B0N 3 VNW pch L=4e-08 W=2.1e-07 
M10 Y 3 VDD VNW pch L=4e-08 W=2.1e-07 
M11 VDD 3 Y VNW pch L=4e-08 W=2.1e-07 
M12 10 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y A0 10 VNW pch L=4e-08 W=4e-07 
M14 11 A0 Y VNW pch L=4e-08 W=4e-07 
M15 VDD A1 11 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI22BB_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 13 B1N VSS VPW nch L=4e-08 W=3.45e-07 
M1 3 B0N 13 VPW nch L=4e-08 W=3.45e-07 
M2 VSS A0 4 VPW nch L=4e-08 W=3.6e-07 
M3 4 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M4 VSS A1 4 VPW nch L=4e-08 W=3.6e-07 
M5 4 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M6 Y 3 4 VPW nch L=4e-08 W=3.6e-07 
M7 4 3 Y VPW nch L=4e-08 W=3.6e-07 
M8 3 B1N VDD VNW pch L=4e-08 W=3e-07 
M9 VDD B0N 3 VNW pch L=4e-08 W=3e-07 
M10 10 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M11 Y A0 10 VNW pch L=4e-08 W=3.8e-07 
M12 11 A0 Y VNW pch L=4e-08 W=3.8e-07 
M13 VDD A1 11 VNW pch L=4e-08 W=3.8e-07 
M14 12 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M15 Y A0 12 VNW pch L=4e-08 W=3.8e-07 
M16 VDD 3 Y VNW pch L=4e-08 W=3.15e-07 
M17 Y 3 VDD VNW pch L=4e-08 W=3.15e-07 
.ENDS


.SUBCKT OAI22BB_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 14 B1N VSS VPW nch L=4e-08 W=2.5e-07 
M1 3 B0N 14 VPW nch L=4e-08 W=2.5e-07 
M2 15 B0N 3 VPW nch L=4e-08 W=2.5e-07 
M3 VSS B1N 15 VPW nch L=4e-08 W=2.5e-07 
M4 5 3 Y VPW nch L=4e-08 W=3.2e-07 
M5 Y 3 5 VPW nch L=4e-08 W=3.2e-07 
M6 5 3 Y VPW nch L=4e-08 W=3.2e-07 
M7 VSS A1 5 VPW nch L=4e-08 W=3.2e-07 
M8 5 A0 VSS VPW nch L=4e-08 W=3.2e-07 
M9 VSS A0 5 VPW nch L=4e-08 W=3.2e-07 
M10 5 A1 VSS VPW nch L=4e-08 W=3.2e-07 
M11 VSS A1 5 VPW nch L=4e-08 W=3.2e-07 
M12 5 A0 VSS VPW nch L=4e-08 W=3.2e-07 
M13 3 B1N VDD VNW pch L=4e-08 W=2.2e-07 
M14 VDD B0N 3 VNW pch L=4e-08 W=2.2e-07 
M15 3 B0N VDD VNW pch L=4e-08 W=2.2e-07 
M16 VDD B1N 3 VNW pch L=4e-08 W=2.2e-07 
M17 VDD 3 Y VNW pch L=4e-08 W=2.8e-07 
M18 Y 3 VDD VNW pch L=4e-08 W=2.8e-07 
M19 VDD 3 Y VNW pch L=4e-08 W=2.8e-07 
M20 10 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M21 Y A0 10 VNW pch L=4e-08 W=3.8e-07 
M22 11 A0 Y VNW pch L=4e-08 W=3.8e-07 
M23 VDD A1 11 VNW pch L=4e-08 W=3.8e-07 
M24 12 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M25 Y A0 12 VNW pch L=4e-08 W=3.8e-07 
M26 13 A0 Y VNW pch L=4e-08 W=3.8e-07 
M27 VDD A1 13 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT OAI22BB_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 16 B1N VSS VPW nch L=4e-08 W=3.55e-07 
M1 3 B0N 16 VPW nch L=4e-08 W=3.55e-07 
M2 17 B0N 3 VPW nch L=4e-08 W=3.55e-07 
M3 VSS B1N 17 VPW nch L=4e-08 W=3.55e-07 
M4 Y 3 4 VPW nch L=4e-08 W=3.6e-07 
M5 4 3 Y VPW nch L=4e-08 W=3.6e-07 
M6 Y 3 4 VPW nch L=4e-08 W=3.6e-07 
M7 4 3 Y VPW nch L=4e-08 W=3.6e-07 
M8 VSS A1 4 VPW nch L=4e-08 W=3.6e-07 
M9 4 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M10 VSS A0 4 VPW nch L=4e-08 W=3.6e-07 
M11 4 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M12 VSS A1 4 VPW nch L=4e-08 W=3.6e-07 
M13 4 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M14 VSS A0 4 VPW nch L=4e-08 W=3.6e-07 
M15 4 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M16 3 B1N VDD VNW pch L=4e-08 W=3.05e-07 
M17 VDD B0N 3 VNW pch L=4e-08 W=3.05e-07 
M18 3 B0N VDD VNW pch L=4e-08 W=3.05e-07 
M19 VDD B1N 3 VNW pch L=4e-08 W=3.05e-07 
M20 Y 3 VDD VNW pch L=4e-08 W=3.15e-07 
M21 VDD 3 Y VNW pch L=4e-08 W=3.15e-07 
M22 Y 3 VDD VNW pch L=4e-08 W=3.15e-07 
M23 VDD 3 Y VNW pch L=4e-08 W=3.15e-07 
M24 10 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M25 Y A0 10 VNW pch L=4e-08 W=3.8e-07 
M26 11 A0 Y VNW pch L=4e-08 W=3.8e-07 
M27 VDD A1 11 VNW pch L=4e-08 W=3.8e-07 
M28 12 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M29 Y A0 12 VNW pch L=4e-08 W=3.8e-07 
M30 13 A0 Y VNW pch L=4e-08 W=3.8e-07 
M31 VDD A1 13 VNW pch L=4e-08 W=3.8e-07 
M32 14 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M33 Y A0 14 VNW pch L=4e-08 W=3.8e-07 
M34 15 A0 Y VNW pch L=4e-08 W=3.8e-07 
M35 VDD A1 15 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT OAI22BB_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0N B1N
M0 18 B0N 1 VPW nch L=4e-08 W=3.25e-07 
M1 VSS B1N 18 VPW nch L=4e-08 W=3.25e-07 
M2 19 B1N VSS VPW nch L=4e-08 W=3.25e-07 
M3 1 B0N 19 VPW nch L=4e-08 W=3.25e-07 
M4 20 B0N 1 VPW nch L=4e-08 W=3.25e-07 
M5 VSS B1N 20 VPW nch L=4e-08 W=3.25e-07 
M6 5 1 Y VPW nch L=4e-08 W=3.85e-07 
M7 Y 1 5 VPW nch L=4e-08 W=3.85e-07 
M8 5 1 Y VPW nch L=4e-08 W=3.85e-07 
M9 Y 1 5 VPW nch L=4e-08 W=3.85e-07 
M10 5 1 Y VPW nch L=4e-08 W=3.85e-07 
M11 VSS A1 5 VPW nch L=4e-08 W=3.85e-07 
M12 5 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M13 VSS A0 5 VPW nch L=4e-08 W=3.85e-07 
M14 5 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M15 VSS A1 5 VPW nch L=4e-08 W=3.85e-07 
M16 5 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M17 VSS A0 5 VPW nch L=4e-08 W=3.85e-07 
M18 5 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M19 VSS A1 5 VPW nch L=4e-08 W=3.85e-07 
M20 5 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M21 1 B0N VDD VNW pch L=4e-08 W=2.8e-07 
M22 VDD B1N 1 VNW pch L=4e-08 W=2.8e-07 
M23 1 B1N VDD VNW pch L=4e-08 W=2.8e-07 
M24 VDD B0N 1 VNW pch L=4e-08 W=2.8e-07 
M25 1 B0N VDD VNW pch L=4e-08 W=2.8e-07 
M26 VDD B1N 1 VNW pch L=4e-08 W=2.8e-07 
M27 VDD 1 Y VNW pch L=4e-08 W=3.35e-07 
M28 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
M29 VDD 1 Y VNW pch L=4e-08 W=3.35e-07 
M30 Y 1 VDD VNW pch L=4e-08 W=3.35e-07 
M31 VDD 1 Y VNW pch L=4e-08 W=3.35e-07 
M32 10 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M33 Y A0 10 VNW pch L=4e-08 W=3.8e-07 
M34 11 A0 Y VNW pch L=4e-08 W=3.8e-07 
M35 VDD A1 11 VNW pch L=4e-08 W=3.8e-07 
M36 12 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M37 Y A0 12 VNW pch L=4e-08 W=3.8e-07 
M38 13 A0 Y VNW pch L=4e-08 W=3.8e-07 
M39 VDD A1 13 VNW pch L=4e-08 W=3.8e-07 
M40 14 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M41 Y A0 14 VNW pch L=4e-08 W=3.8e-07 
M42 15 A0 Y VNW pch L=4e-08 W=3.8e-07 
M43 VDD A1 15 VNW pch L=4e-08 W=3.8e-07 
M44 16 A1 VDD VNW pch L=4e-08 W=3.8e-07 
M45 Y A0 16 VNW pch L=4e-08 W=3.8e-07 
M46 17 A0 Y VNW pch L=4e-08 W=3.8e-07 
M47 VDD A1 17 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT OAI22_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=2.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.1e-07 
M2 Y B0 1 VPW nch L=4e-08 W=2.1e-07 
M3 1 B1 Y VPW nch L=4e-08 W=2.1e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=2e-07 
M5 Y A0 9 VNW pch L=4e-08 W=2e-07 
M6 10 B0 Y VNW pch L=4e-08 W=2e-07 
M7 VDD B1 10 VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OAI22_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=2.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.1e-07 
M2 Y B0 1 VPW nch L=4e-08 W=2.1e-07 
M3 1 B1 Y VPW nch L=4e-08 W=2.1e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M5 Y A0 9 VNW pch L=4e-08 W=2.85e-07 
M6 10 B0 Y VNW pch L=4e-08 W=2.85e-07 
M7 VDD B1 10 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OAI22_X1M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 Y B0 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 B1 Y VPW nch L=4e-08 W=2.4e-07 
M4 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M5 Y A0 9 VNW pch L=4e-08 W=4e-07 
M6 10 B0 Y VNW pch L=4e-08 W=4e-07 
M7 VDD B1 10 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI22_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=2.1e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.1e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.1e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.1e-07 
M4 Y B1 1 VPW nch L=4e-08 W=2.1e-07 
M5 1 B0 Y VPW nch L=4e-08 W=2.1e-07 
M6 Y B0 1 VPW nch L=4e-08 W=2.1e-07 
M7 1 B1 Y VPW nch L=4e-08 W=2.1e-07 
M8 9 A1 VDD VNW pch L=4e-08 W=2.85e-07 
M9 Y A0 9 VNW pch L=4e-08 W=2.85e-07 
M10 10 A0 Y VNW pch L=4e-08 W=2.85e-07 
M11 VDD A1 10 VNW pch L=4e-08 W=2.85e-07 
M12 11 B1 VDD VNW pch L=4e-08 W=2.85e-07 
M13 Y B0 11 VNW pch L=4e-08 W=2.85e-07 
M14 12 B0 Y VNW pch L=4e-08 W=2.85e-07 
M15 VDD B1 12 VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OAI22_X2M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 1 VPW nch L=4e-08 W=2.4e-07 
M1 1 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A0 1 VPW nch L=4e-08 W=2.4e-07 
M3 1 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M4 Y B1 1 VPW nch L=4e-08 W=2.4e-07 
M5 1 B0 Y VPW nch L=4e-08 W=2.4e-07 
M6 Y B0 1 VPW nch L=4e-08 W=2.4e-07 
M7 1 B1 Y VPW nch L=4e-08 W=2.4e-07 
M8 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M9 Y A0 9 VNW pch L=4e-08 W=4e-07 
M10 10 A0 Y VNW pch L=4e-08 W=4e-07 
M11 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M12 11 B1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y B0 11 VNW pch L=4e-08 W=4e-07 
M14 12 B0 Y VNW pch L=4e-08 W=4e-07 
M15 VDD B1 12 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI22_X3M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A0 2 VPW nch L=4e-08 W=3.6e-07 
M1 2 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M2 VSS A1 2 VPW nch L=4e-08 W=3.6e-07 
M3 2 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M4 Y B0 2 VPW nch L=4e-08 W=3.6e-07 
M5 2 B1 Y VPW nch L=4e-08 W=3.6e-07 
M6 Y B1 2 VPW nch L=4e-08 W=3.6e-07 
M7 2 B0 Y VPW nch L=4e-08 W=3.6e-07 
M8 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M9 Y A0 9 VNW pch L=4e-08 W=4e-07 
M10 10 A0 Y VNW pch L=4e-08 W=4e-07 
M11 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M12 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y A0 11 VNW pch L=4e-08 W=4e-07 
M14 12 B0 Y VNW pch L=4e-08 W=4e-07 
M15 VDD B1 12 VNW pch L=4e-08 W=4e-07 
M16 13 B1 VDD VNW pch L=4e-08 W=4e-07 
M17 Y B0 13 VNW pch L=4e-08 W=4e-07 
M18 14 B0 Y VNW pch L=4e-08 W=4e-07 
M19 VDD B1 14 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI22_X4M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A0 2 VPW nch L=4e-08 W=3.2e-07 
M1 2 A1 VSS VPW nch L=4e-08 W=3.2e-07 
M2 VSS A1 2 VPW nch L=4e-08 W=3.2e-07 
M3 2 A0 VSS VPW nch L=4e-08 W=3.2e-07 
M4 VSS A0 2 VPW nch L=4e-08 W=3.2e-07 
M5 2 A1 VSS VPW nch L=4e-08 W=3.2e-07 
M6 Y B1 2 VPW nch L=4e-08 W=3.2e-07 
M7 2 B0 Y VPW nch L=4e-08 W=3.2e-07 
M8 Y B0 2 VPW nch L=4e-08 W=3.2e-07 
M9 2 B1 Y VPW nch L=4e-08 W=3.2e-07 
M10 Y B1 2 VPW nch L=4e-08 W=3.2e-07 
M11 2 B0 Y VPW nch L=4e-08 W=3.2e-07 
M12 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y A0 9 VNW pch L=4e-08 W=4e-07 
M14 10 A0 Y VNW pch L=4e-08 W=4e-07 
M15 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M16 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M17 Y A0 11 VNW pch L=4e-08 W=4e-07 
M18 12 A0 Y VNW pch L=4e-08 W=4e-07 
M19 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M20 13 B1 VDD VNW pch L=4e-08 W=4e-07 
M21 Y B0 13 VNW pch L=4e-08 W=4e-07 
M22 14 B0 Y VNW pch L=4e-08 W=4e-07 
M23 VDD B1 14 VNW pch L=4e-08 W=4e-07 
M24 15 B1 VDD VNW pch L=4e-08 W=4e-07 
M25 Y B0 15 VNW pch L=4e-08 W=4e-07 
M26 16 B0 Y VNW pch L=4e-08 W=4e-07 
M27 VDD B1 16 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI22_X6M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A1 3 VPW nch L=4e-08 W=3.6e-07 
M1 3 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M2 VSS A0 3 VPW nch L=4e-08 W=3.6e-07 
M3 3 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M4 VSS A1 3 VPW nch L=4e-08 W=3.6e-07 
M5 3 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M6 VSS A0 3 VPW nch L=4e-08 W=3.6e-07 
M7 3 A1 VSS VPW nch L=4e-08 W=3.6e-07 
M8 Y B1 3 VPW nch L=4e-08 W=3.6e-07 
M9 3 B0 Y VPW nch L=4e-08 W=3.6e-07 
M10 Y B0 3 VPW nch L=4e-08 W=3.6e-07 
M11 3 B1 Y VPW nch L=4e-08 W=3.6e-07 
M12 Y B1 3 VPW nch L=4e-08 W=3.6e-07 
M13 3 B0 Y VPW nch L=4e-08 W=3.6e-07 
M14 Y B0 3 VPW nch L=4e-08 W=3.6e-07 
M15 3 B1 Y VPW nch L=4e-08 W=3.6e-07 
M16 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M17 Y A0 9 VNW pch L=4e-08 W=4e-07 
M18 10 A0 Y VNW pch L=4e-08 W=4e-07 
M19 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M20 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M21 Y A0 11 VNW pch L=4e-08 W=4e-07 
M22 12 A0 Y VNW pch L=4e-08 W=4e-07 
M23 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M24 13 A1 VDD VNW pch L=4e-08 W=4e-07 
M25 Y A0 13 VNW pch L=4e-08 W=4e-07 
M26 14 A0 Y VNW pch L=4e-08 W=4e-07 
M27 VDD A1 14 VNW pch L=4e-08 W=4e-07 
M28 15 B1 VDD VNW pch L=4e-08 W=4e-07 
M29 Y B0 15 VNW pch L=4e-08 W=4e-07 
M30 16 B0 Y VNW pch L=4e-08 W=4e-07 
M31 VDD B1 16 VNW pch L=4e-08 W=4e-07 
M32 17 B1 VDD VNW pch L=4e-08 W=4e-07 
M33 Y B0 17 VNW pch L=4e-08 W=4e-07 
M34 18 B0 Y VNW pch L=4e-08 W=4e-07 
M35 VDD B1 18 VNW pch L=4e-08 W=4e-07 
M36 19 B1 VDD VNW pch L=4e-08 W=4e-07 
M37 Y B0 19 VNW pch L=4e-08 W=4e-07 
M38 20 B0 Y VNW pch L=4e-08 W=4e-07 
M39 VDD B1 20 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI22_X8M_A9TR Y VDD VNW VPW VSS A0 A1 B0 B1
M0 VSS A0 3 VPW nch L=4e-08 W=3.85e-07 
M1 3 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M2 VSS A1 3 VPW nch L=4e-08 W=3.85e-07 
M3 3 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M4 VSS A0 3 VPW nch L=4e-08 W=3.85e-07 
M5 3 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M6 VSS A1 3 VPW nch L=4e-08 W=3.85e-07 
M7 3 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M8 VSS A0 3 VPW nch L=4e-08 W=3.85e-07 
M9 3 A1 VSS VPW nch L=4e-08 W=3.85e-07 
M10 Y B1 3 VPW nch L=4e-08 W=3.85e-07 
M11 3 B0 Y VPW nch L=4e-08 W=3.85e-07 
M12 Y B0 3 VPW nch L=4e-08 W=3.85e-07 
M13 3 B1 Y VPW nch L=4e-08 W=3.85e-07 
M14 Y B1 3 VPW nch L=4e-08 W=3.85e-07 
M15 3 B0 Y VPW nch L=4e-08 W=3.85e-07 
M16 Y B0 3 VPW nch L=4e-08 W=3.85e-07 
M17 3 B1 Y VPW nch L=4e-08 W=3.85e-07 
M18 Y B1 3 VPW nch L=4e-08 W=3.85e-07 
M19 3 B0 Y VPW nch L=4e-08 W=3.85e-07 
M20 9 A1 VDD VNW pch L=4e-08 W=4e-07 
M21 Y A0 9 VNW pch L=4e-08 W=4e-07 
M22 10 A0 Y VNW pch L=4e-08 W=4e-07 
M23 VDD A1 10 VNW pch L=4e-08 W=4e-07 
M24 11 A1 VDD VNW pch L=4e-08 W=4e-07 
M25 Y A0 11 VNW pch L=4e-08 W=4e-07 
M26 12 A0 Y VNW pch L=4e-08 W=4e-07 
M27 VDD A1 12 VNW pch L=4e-08 W=4e-07 
M28 13 A1 VDD VNW pch L=4e-08 W=4e-07 
M29 Y A0 13 VNW pch L=4e-08 W=4e-07 
M30 14 A0 Y VNW pch L=4e-08 W=4e-07 
M31 VDD A1 14 VNW pch L=4e-08 W=4e-07 
M32 15 A1 VDD VNW pch L=4e-08 W=4e-07 
M33 Y A0 15 VNW pch L=4e-08 W=4e-07 
M34 16 A0 Y VNW pch L=4e-08 W=4e-07 
M35 VDD A1 16 VNW pch L=4e-08 W=4e-07 
M36 17 B1 VDD VNW pch L=4e-08 W=4e-07 
M37 Y B0 17 VNW pch L=4e-08 W=4e-07 
M38 18 B0 Y VNW pch L=4e-08 W=4e-07 
M39 VDD B1 18 VNW pch L=4e-08 W=4e-07 
M40 19 B1 VDD VNW pch L=4e-08 W=4e-07 
M41 Y B0 19 VNW pch L=4e-08 W=4e-07 
M42 20 B0 Y VNW pch L=4e-08 W=4e-07 
M43 VDD B1 20 VNW pch L=4e-08 W=4e-07 
M44 21 B1 VDD VNW pch L=4e-08 W=4e-07 
M45 Y B0 21 VNW pch L=4e-08 W=4e-07 
M46 22 B0 Y VNW pch L=4e-08 W=4e-07 
M47 VDD B1 22 VNW pch L=4e-08 W=4e-07 
M48 23 B1 VDD VNW pch L=4e-08 W=4e-07 
M49 Y B0 23 VNW pch L=4e-08 W=4e-07 
M50 24 B0 Y VNW pch L=4e-08 W=4e-07 
M51 VDD B1 24 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OAI2XB1_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 VSS A1N 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS 1 4 VPW nch L=4e-08 W=1.4e-07 
M2 4 A0 VSS VPW nch L=4e-08 W=1.4e-07 
M3 Y B0 4 VPW nch L=4e-08 W=1.4e-07 
M4 VDD A1N 1 VNW pch L=4e-08 W=1.55e-07 
M5 9 1 VDD VNW pch L=4e-08 W=2.3e-07 
M6 Y A0 9 VNW pch L=4e-08 W=2.3e-07 
M7 VDD B0 Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT OAI2XB1_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 VSS A1N 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS 1 4 VPW nch L=4e-08 W=1.7e-07 
M2 4 A0 VSS VPW nch L=4e-08 W=1.7e-07 
M3 Y B0 4 VPW nch L=4e-08 W=1.7e-07 
M4 VDD A1N 1 VNW pch L=4e-08 W=1.55e-07 
M5 9 1 VDD VNW pch L=4e-08 W=2.85e-07 
M6 Y A0 9 VNW pch L=4e-08 W=2.85e-07 
M7 VDD B0 Y VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT OAI2XB1_X1M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 VSS A1N 1 VPW nch L=4e-08 W=1.2e-07 
M1 VSS 1 4 VPW nch L=4e-08 W=2.4e-07 
M2 4 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M3 Y B0 4 VPW nch L=4e-08 W=2.4e-07 
M4 VDD A1N 1 VNW pch L=4e-08 W=1.55e-07 
M5 9 1 VDD VNW pch L=4e-08 W=4e-07 
M6 Y A0 9 VNW pch L=4e-08 W=4e-07 
M7 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI2XB1_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 VSS A1N 1 VPW nch L=4e-08 W=1.25e-07 
M1 VSS A0 4 VPW nch L=4e-08 W=3.4e-07 
M2 4 1 VSS VPW nch L=4e-08 W=3.4e-07 
M3 Y B0 4 VPW nch L=4e-08 W=3.4e-07 
M4 VDD A1N 1 VNW pch L=4e-08 W=1.6e-07 
M5 9 1 VDD VNW pch L=4e-08 W=2.85e-07 
M6 Y A0 9 VNW pch L=4e-08 W=2.85e-07 
M7 10 A0 Y VNW pch L=4e-08 W=2.85e-07 
M8 VDD 1 10 VNW pch L=4e-08 W=2.85e-07 
M9 Y B0 VDD VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT OAI2XB1_X2M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 VSS A1N 1 VPW nch L=4e-08 W=1.65e-07 
M1 VSS 1 4 VPW nch L=4e-08 W=2.4e-07 
M2 4 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M3 VSS A0 4 VPW nch L=4e-08 W=2.4e-07 
M4 4 1 VSS VPW nch L=4e-08 W=2.4e-07 
M5 Y B0 4 VPW nch L=4e-08 W=2.4e-07 
M6 4 B0 Y VPW nch L=4e-08 W=2.4e-07 
M7 VDD A1N 1 VNW pch L=4e-08 W=2.1e-07 
M8 9 1 VDD VNW pch L=4e-08 W=4e-07 
M9 Y A0 9 VNW pch L=4e-08 W=4e-07 
M10 10 A0 Y VNW pch L=4e-08 W=4e-07 
M11 VDD 1 10 VNW pch L=4e-08 W=4e-07 
M12 Y B0 VDD VNW pch L=4e-08 W=2.1e-07 
M13 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI2XB1_X3M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 VSS A1N 1 VPW nch L=4e-08 W=2.4e-07 
M1 VSS A0 4 VPW nch L=4e-08 W=3.6e-07 
M2 4 1 VSS VPW nch L=4e-08 W=3.6e-07 
M3 VSS 1 4 VPW nch L=4e-08 W=3.6e-07 
M4 4 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M5 Y B0 4 VPW nch L=4e-08 W=3.6e-07 
M6 4 B0 Y VPW nch L=4e-08 W=3.6e-07 
M7 VDD A1N 1 VNW pch L=4e-08 W=3.1e-07 
M8 9 1 VDD VNW pch L=4e-08 W=4e-07 
M9 Y A0 9 VNW pch L=4e-08 W=4e-07 
M10 10 A0 Y VNW pch L=4e-08 W=4e-07 
M11 VDD 1 10 VNW pch L=4e-08 W=4e-07 
M12 11 1 VDD VNW pch L=4e-08 W=4e-07 
M13 Y A0 11 VNW pch L=4e-08 W=4e-07 
M14 VDD B0 Y VNW pch L=4e-08 W=3.15e-07 
M15 Y B0 VDD VNW pch L=4e-08 W=3.15e-07 
.ENDS


.SUBCKT OAI2XB1_X4M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 VSS A1N 1 VPW nch L=4e-08 W=3.1e-07 
M1 VSS A0 4 VPW nch L=4e-08 W=3.2e-07 
M2 4 1 VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS 1 4 VPW nch L=4e-08 W=3.2e-07 
M4 4 A0 VSS VPW nch L=4e-08 W=3.2e-07 
M5 VSS A0 4 VPW nch L=4e-08 W=3.2e-07 
M6 4 1 VSS VPW nch L=4e-08 W=3.2e-07 
M7 Y B0 4 VPW nch L=4e-08 W=3.2e-07 
M8 4 B0 Y VPW nch L=4e-08 W=3.2e-07 
M9 Y B0 4 VPW nch L=4e-08 W=3.2e-07 
M10 VDD A1N 1 VNW pch L=4e-08 W=4e-07 
M11 9 1 VDD VNW pch L=4e-08 W=4e-07 
M12 Y A0 9 VNW pch L=4e-08 W=4e-07 
M13 10 A0 Y VNW pch L=4e-08 W=4e-07 
M14 VDD 1 10 VNW pch L=4e-08 W=4e-07 
M15 11 1 VDD VNW pch L=4e-08 W=4e-07 
M16 Y A0 11 VNW pch L=4e-08 W=4e-07 
M17 12 A0 Y VNW pch L=4e-08 W=4e-07 
M18 VDD 1 12 VNW pch L=4e-08 W=4e-07 
M19 Y B0 VDD VNW pch L=4e-08 W=2.8e-07 
M20 VDD B0 Y VNW pch L=4e-08 W=2.8e-07 
M21 Y B0 VDD VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT OAI2XB1_X6M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=2.4e-07 
M1 VSS A1N 3 VPW nch L=4e-08 W=2.4e-07 
M2 VSS 3 5 VPW nch L=4e-08 W=3.6e-07 
M3 5 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M4 VSS A0 5 VPW nch L=4e-08 W=3.6e-07 
M5 5 3 VSS VPW nch L=4e-08 W=3.6e-07 
M6 VSS 3 5 VPW nch L=4e-08 W=3.6e-07 
M7 5 A0 VSS VPW nch L=4e-08 W=3.6e-07 
M8 VSS A0 5 VPW nch L=4e-08 W=3.6e-07 
M9 5 3 VSS VPW nch L=4e-08 W=3.6e-07 
M10 Y B0 5 VPW nch L=4e-08 W=3.6e-07 
M11 5 B0 Y VPW nch L=4e-08 W=3.6e-07 
M12 Y B0 5 VPW nch L=4e-08 W=3.6e-07 
M13 5 B0 Y VPW nch L=4e-08 W=3.6e-07 
M14 3 A1N VDD VNW pch L=4e-08 W=3.05e-07 
M15 VDD A1N 3 VNW pch L=4e-08 W=3.05e-07 
M16 9 3 VDD VNW pch L=4e-08 W=4e-07 
M17 Y A0 9 VNW pch L=4e-08 W=4e-07 
M18 10 A0 Y VNW pch L=4e-08 W=4e-07 
M19 VDD 3 10 VNW pch L=4e-08 W=4e-07 
M20 11 3 VDD VNW pch L=4e-08 W=4e-07 
M21 Y A0 11 VNW pch L=4e-08 W=4e-07 
M22 12 A0 Y VNW pch L=4e-08 W=4e-07 
M23 VDD 3 12 VNW pch L=4e-08 W=4e-07 
M24 13 3 VDD VNW pch L=4e-08 W=4e-07 
M25 Y A0 13 VNW pch L=4e-08 W=4e-07 
M26 14 A0 Y VNW pch L=4e-08 W=4e-07 
M27 VDD 3 14 VNW pch L=4e-08 W=4e-07 
M28 Y B0 VDD VNW pch L=4e-08 W=3.15e-07 
M29 VDD B0 Y VNW pch L=4e-08 W=3.15e-07 
M30 Y B0 VDD VNW pch L=4e-08 W=3.15e-07 
M31 VDD B0 Y VNW pch L=4e-08 W=3.15e-07 
.ENDS


.SUBCKT OAI2XB1_X8M_A9TR Y VDD VNW VPW VSS A0 A1N B0
M0 3 A1N VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A1N 3 VPW nch L=4e-08 W=3.1e-07 
M2 VSS A0 5 VPW nch L=4e-08 W=3.85e-07 
M3 5 3 VSS VPW nch L=4e-08 W=3.85e-07 
M4 VSS 3 5 VPW nch L=4e-08 W=3.85e-07 
M5 5 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M6 VSS A0 5 VPW nch L=4e-08 W=3.85e-07 
M7 5 3 VSS VPW nch L=4e-08 W=3.85e-07 
M8 VSS 3 5 VPW nch L=4e-08 W=3.85e-07 
M9 5 A0 VSS VPW nch L=4e-08 W=3.85e-07 
M10 VSS A0 5 VPW nch L=4e-08 W=3.85e-07 
M11 5 3 VSS VPW nch L=4e-08 W=3.85e-07 
M12 Y B0 5 VPW nch L=4e-08 W=3.85e-07 
M13 5 B0 Y VPW nch L=4e-08 W=3.85e-07 
M14 Y B0 5 VPW nch L=4e-08 W=3.85e-07 
M15 5 B0 Y VPW nch L=4e-08 W=3.85e-07 
M16 Y B0 5 VPW nch L=4e-08 W=3.85e-07 
M17 3 A1N VDD VNW pch L=4e-08 W=4e-07 
M18 VDD A1N 3 VNW pch L=4e-08 W=4e-07 
M19 9 3 VDD VNW pch L=4e-08 W=4e-07 
M20 Y A0 9 VNW pch L=4e-08 W=4e-07 
M21 10 A0 Y VNW pch L=4e-08 W=4e-07 
M22 VDD 3 10 VNW pch L=4e-08 W=4e-07 
M23 11 3 VDD VNW pch L=4e-08 W=4e-07 
M24 Y A0 11 VNW pch L=4e-08 W=4e-07 
M25 12 A0 Y VNW pch L=4e-08 W=4e-07 
M26 VDD 3 12 VNW pch L=4e-08 W=4e-07 
M27 13 3 VDD VNW pch L=4e-08 W=4e-07 
M28 Y A0 13 VNW pch L=4e-08 W=4e-07 
M29 14 A0 Y VNW pch L=4e-08 W=4e-07 
M30 VDD 3 14 VNW pch L=4e-08 W=4e-07 
M31 15 3 VDD VNW pch L=4e-08 W=4e-07 
M32 Y A0 15 VNW pch L=4e-08 W=4e-07 
M33 16 A0 Y VNW pch L=4e-08 W=4e-07 
M34 VDD 3 16 VNW pch L=4e-08 W=4e-07 
M35 Y B0 VDD VNW pch L=4e-08 W=3.35e-07 
M36 VDD B0 Y VNW pch L=4e-08 W=3.35e-07 
M37 Y B0 VDD VNW pch L=4e-08 W=3.35e-07 
M38 VDD B0 Y VNW pch L=4e-08 W=3.35e-07 
M39 Y B0 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT OAI31_X0P5M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 3 A2 VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS A1 3 VPW nch L=4e-08 W=1.2e-07 
M2 3 A0 VSS VPW nch L=4e-08 W=1.2e-07 
M3 Y B0 3 VPW nch L=4e-08 W=1.2e-07 
M4 9 A2 VDD VNW pch L=4e-08 W=2e-07 
M5 10 A1 9 VNW pch L=4e-08 W=2e-07 
M6 Y A0 10 VNW pch L=4e-08 W=2e-07 
M7 VDD B0 Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT OAI31_X0P7M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 3 A2 VSS VPW nch L=4e-08 W=1.4e-07 
M1 VSS A1 3 VPW nch L=4e-08 W=1.4e-07 
M2 3 A0 VSS VPW nch L=4e-08 W=1.4e-07 
M3 Y B0 3 VPW nch L=4e-08 W=1.4e-07 
M4 9 A2 VDD VNW pch L=4e-08 W=3.45e-07 
M5 10 A1 9 VNW pch L=4e-08 W=3.45e-07 
M6 Y A0 10 VNW pch L=4e-08 W=3.45e-07 
M7 VDD B0 Y VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT OAI31_X1M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 3 A2 VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS A1 3 VPW nch L=4e-08 W=1.6e-07 
M2 3 A0 VSS VPW nch L=4e-08 W=1.6e-07 
M3 Y B0 3 VPW nch L=4e-08 W=1.6e-07 
M4 9 A2 VDD VNW pch L=4e-08 W=4e-07 
M5 10 A1 9 VNW pch L=4e-08 W=4e-07 
M6 Y A0 10 VNW pch L=4e-08 W=4e-07 
M7 VDD B0 Y VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT OAI31_X1P4M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 4 A2 VSS VPW nch L=4e-08 W=2.3e-07 
M1 VSS A1 4 VPW nch L=4e-08 W=2.3e-07 
M2 4 A0 VSS VPW nch L=4e-08 W=2.3e-07 
M3 Y B0 4 VPW nch L=4e-08 W=2.3e-07 
M4 VDD A2 1 VNW pch L=4e-08 W=2.85e-07 
M5 1 A2 VDD VNW pch L=4e-08 W=2.85e-07 
M6 10 A1 1 VNW pch L=4e-08 W=2.85e-07 
M7 Y A0 10 VNW pch L=4e-08 W=2.85e-07 
M8 11 A0 Y VNW pch L=4e-08 W=2.85e-07 
M9 1 A1 11 VNW pch L=4e-08 W=2.85e-07 
M10 Y B0 VDD VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT OAI31_X2M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 4 A2 VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS A1 4 VPW nch L=4e-08 W=3.2e-07 
M2 4 A0 VSS VPW nch L=4e-08 W=3.2e-07 
M3 Y B0 4 VPW nch L=4e-08 W=3.2e-07 
M4 VDD A2 1 VNW pch L=4e-08 W=4e-07 
M5 1 A2 VDD VNW pch L=4e-08 W=4e-07 
M6 10 A1 1 VNW pch L=4e-08 W=4e-07 
M7 Y A0 10 VNW pch L=4e-08 W=4e-07 
M8 11 A0 Y VNW pch L=4e-08 W=4e-07 
M9 1 A1 11 VNW pch L=4e-08 W=4e-07 
M10 Y B0 VDD VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT OAI31_X3M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 VSS A2 2 VPW nch L=4e-08 W=2.4e-07 
M1 2 A2 VSS VPW nch L=4e-08 W=2.4e-07 
M2 VSS A1 2 VPW nch L=4e-08 W=2.4e-07 
M3 2 A0 VSS VPW nch L=4e-08 W=2.4e-07 
M4 VSS A0 2 VPW nch L=4e-08 W=2.4e-07 
M5 2 A1 VSS VPW nch L=4e-08 W=2.4e-07 
M6 Y B0 2 VPW nch L=4e-08 W=2.4e-07 
M7 2 B0 Y VPW nch L=4e-08 W=2.4e-07 
M8 3 A2 VDD VNW pch L=4e-08 W=4e-07 
M9 VDD A2 3 VNW pch L=4e-08 W=4e-07 
M10 3 A2 VDD VNW pch L=4e-08 W=4e-07 
M11 10 A1 3 VNW pch L=4e-08 W=4e-07 
M12 Y A0 10 VNW pch L=4e-08 W=4e-07 
M13 11 A0 Y VNW pch L=4e-08 W=4e-07 
M14 3 A1 11 VNW pch L=4e-08 W=4e-07 
M15 12 A1 3 VNW pch L=4e-08 W=4e-07 
M16 Y A0 12 VNW pch L=4e-08 W=4e-07 
M17 VDD B0 Y VNW pch L=4e-08 W=2.1e-07 
M18 Y B0 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OAI31_X4M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 VSS A2 3 VPW nch L=4e-08 W=3.2e-07 
M1 3 A2 VSS VPW nch L=4e-08 W=3.2e-07 
M2 VSS A1 3 VPW nch L=4e-08 W=3.2e-07 
M3 3 A0 VSS VPW nch L=4e-08 W=3.2e-07 
M4 VSS A0 3 VPW nch L=4e-08 W=3.2e-07 
M5 3 A1 VSS VPW nch L=4e-08 W=3.2e-07 
M6 Y B0 3 VPW nch L=4e-08 W=3.2e-07 
M7 3 B0 Y VPW nch L=4e-08 W=3.2e-07 
M8 VDD A2 1 VNW pch L=4e-08 W=4e-07 
M9 1 A2 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD A2 1 VNW pch L=4e-08 W=4e-07 
M11 1 A2 VDD VNW pch L=4e-08 W=4e-07 
M12 10 A1 1 VNW pch L=4e-08 W=4e-07 
M13 Y A0 10 VNW pch L=4e-08 W=4e-07 
M14 11 A0 Y VNW pch L=4e-08 W=4e-07 
M15 1 A1 11 VNW pch L=4e-08 W=4e-07 
M16 12 A1 1 VNW pch L=4e-08 W=4e-07 
M17 Y A0 12 VNW pch L=4e-08 W=4e-07 
M18 13 A0 Y VNW pch L=4e-08 W=4e-07 
M19 1 A1 13 VNW pch L=4e-08 W=4e-07 
M20 Y B0 VDD VNW pch L=4e-08 W=2.8e-07 
M21 VDD B0 Y VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT OAI31_X6M_A9TR Y VDD VNW VPW VSS A0 A1 A2 B0
M0 4 A2 VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS A2 4 VPW nch L=4e-08 W=3.2e-07 
M2 4 A2 VSS VPW nch L=4e-08 W=3.2e-07 
M3 4 A0 VSS VPW nch L=4e-08 W=3.2e-07 
M4 VSS A1 4 VPW nch L=4e-08 W=3.2e-07 
M5 4 A1 VSS VPW nch L=4e-08 W=3.2e-07 
M6 VSS A0 4 VPW nch L=4e-08 W=3.2e-07 
M7 4 A0 VSS VPW nch L=4e-08 W=3.2e-07 
M8 VSS A1 4 VPW nch L=4e-08 W=3.2e-07 
M9 Y B0 4 VPW nch L=4e-08 W=3.2e-07 
M10 4 B0 Y VPW nch L=4e-08 W=3.2e-07 
M11 Y B0 4 VPW nch L=4e-08 W=3.2e-07 
M12 VDD A2 1 VNW pch L=4e-08 W=4e-07 
M13 1 A2 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD A2 1 VNW pch L=4e-08 W=4e-07 
M15 1 A2 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD A2 1 VNW pch L=4e-08 W=4e-07 
M17 1 A2 VDD VNW pch L=4e-08 W=4e-07 
M18 10 A1 1 VNW pch L=4e-08 W=4e-07 
M19 Y A0 10 VNW pch L=4e-08 W=4e-07 
M20 11 A0 Y VNW pch L=4e-08 W=4e-07 
M21 1 A1 11 VNW pch L=4e-08 W=4e-07 
M22 12 A1 1 VNW pch L=4e-08 W=4e-07 
M23 Y A0 12 VNW pch L=4e-08 W=4e-07 
M24 13 A0 Y VNW pch L=4e-08 W=4e-07 
M25 1 A1 13 VNW pch L=4e-08 W=4e-07 
M26 14 A1 1 VNW pch L=4e-08 W=4e-07 
M27 Y A0 14 VNW pch L=4e-08 W=4e-07 
M28 15 A0 Y VNW pch L=4e-08 W=4e-07 
M29 1 A1 15 VNW pch L=4e-08 W=4e-07 
M30 Y B0 VDD VNW pch L=4e-08 W=2.8e-07 
M31 VDD B0 Y VNW pch L=4e-08 W=2.8e-07 
M32 Y B0 VDD VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT OR2_X0P5B_A9TR Y VDD VNW VPW VSS A B
M0 2 A VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=1.2e-07 
M3 7 A 2 VNW pch L=4e-08 W=3.6e-07 
M4 VDD B 7 VNW pch L=4e-08 W=3.6e-07 
M5 Y 2 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT OR2_X0P5M_A9TR Y VDD VNW VPW VSS A B
M0 2 A VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=1.55e-07 
M3 7 A 2 VNW pch L=4e-08 W=2.95e-07 
M4 VDD B 7 VNW pch L=4e-08 W=2.95e-07 
M5 Y 2 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OR2_X0P7B_A9TR Y VDD VNW VPW VSS A B
M0 2 A VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=1.6e-07 
M3 7 A 2 VNW pch L=4e-08 W=3.6e-07 
M4 VDD B 7 VNW pch L=4e-08 W=3.6e-07 
M5 Y 2 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OR2_X0P7M_A9TR Y VDD VNW VPW VSS A B
M0 2 A VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=2.2e-07 
M3 7 A 2 VNW pch L=4e-08 W=2.95e-07 
M4 VDD B 7 VNW pch L=4e-08 W=2.95e-07 
M5 Y 2 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OR2_X11B_A9TR Y VDD VNW VPW VSS A B
M0 1 A VSS VPW nch L=4e-08 W=3.8e-07 
M1 VSS B 1 VPW nch L=4e-08 W=3.8e-07 
M2 1 B VSS VPW nch L=4e-08 W=3.8e-07 
M3 VSS A 1 VPW nch L=4e-08 W=3.8e-07 
M4 1 A VSS VPW nch L=4e-08 W=3.8e-07 
M5 VSS B 1 VPW nch L=4e-08 W=3.8e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.55e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M9 VSS 1 Y VPW nch L=4e-08 W=3.55e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M11 VSS 1 Y VPW nch L=4e-08 W=3.55e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M13 7 A 1 VNW pch L=4e-08 W=3.8e-07 
M14 VDD B 7 VNW pch L=4e-08 W=3.8e-07 
M15 8 B VDD VNW pch L=4e-08 W=3.8e-07 
M16 1 A 8 VNW pch L=4e-08 W=3.8e-07 
M17 9 A 1 VNW pch L=4e-08 W=3.8e-07 
M18 VDD B 9 VNW pch L=4e-08 W=3.8e-07 
M19 10 B VDD VNW pch L=4e-08 W=3.8e-07 
M20 1 A 10 VNW pch L=4e-08 W=3.8e-07 
M21 11 A 1 VNW pch L=4e-08 W=3.8e-07 
M22 VDD B 11 VNW pch L=4e-08 W=3.8e-07 
M23 12 B VDD VNW pch L=4e-08 W=3.8e-07 
M24 1 A 12 VNW pch L=4e-08 W=3.8e-07 
M25 13 A 1 VNW pch L=4e-08 W=3.8e-07 
M26 VDD B 13 VNW pch L=4e-08 W=3.8e-07 
M27 14 B VDD VNW pch L=4e-08 W=3.8e-07 
M28 1 A 14 VNW pch L=4e-08 W=3.8e-07 
M29 15 A 1 VNW pch L=4e-08 W=3.8e-07 
M30 VDD B 15 VNW pch L=4e-08 W=3.8e-07 
M31 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M33 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M35 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M37 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M39 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M41 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X11M_A9TR Y VDD VNW VPW VSS A B
M0 1 A VSS VPW nch L=4e-08 W=3.7e-07 
M1 VSS B 1 VPW nch L=4e-08 W=3.7e-07 
M2 1 B VSS VPW nch L=4e-08 W=3.7e-07 
M3 VSS A 1 VPW nch L=4e-08 W=3.7e-07 
M4 1 A VSS VPW nch L=4e-08 W=3.7e-07 
M5 VSS B 1 VPW nch L=4e-08 W=3.7e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=3.8e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.8e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.8e-07 
M9 VSS 1 Y VPW nch L=4e-08 W=3.8e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=3.8e-07 
M11 VSS 1 Y VPW nch L=4e-08 W=3.8e-07 
M12 Y 1 VSS VPW nch L=4e-08 W=3.8e-07 
M13 VSS 1 Y VPW nch L=4e-08 W=3.8e-07 
M14 Y 1 VSS VPW nch L=4e-08 W=3.8e-07 
M15 7 A 1 VNW pch L=4e-08 W=4e-07 
M16 VDD B 7 VNW pch L=4e-08 W=4e-07 
M17 8 B VDD VNW pch L=4e-08 W=4e-07 
M18 1 A 8 VNW pch L=4e-08 W=4e-07 
M19 9 A 1 VNW pch L=4e-08 W=4e-07 
M20 VDD B 9 VNW pch L=4e-08 W=4e-07 
M21 10 B VDD VNW pch L=4e-08 W=4e-07 
M22 1 A 10 VNW pch L=4e-08 W=4e-07 
M23 11 A 1 VNW pch L=4e-08 W=4e-07 
M24 VDD B 11 VNW pch L=4e-08 W=4e-07 
M25 12 B VDD VNW pch L=4e-08 W=4e-07 
M26 1 A 12 VNW pch L=4e-08 W=4e-07 
M27 13 A 1 VNW pch L=4e-08 W=4e-07 
M28 VDD B 13 VNW pch L=4e-08 W=4e-07 
M29 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M31 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M33 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M35 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M37 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M39 Y 1 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X1B_A9TR Y VDD VNW VPW VSS A B
M0 2 A VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=2.25e-07 
M3 7 A 2 VNW pch L=4e-08 W=3.6e-07 
M4 VDD B 7 VNW pch L=4e-08 W=3.6e-07 
M5 Y 2 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X1M_A9TR Y VDD VNW VPW VSS A B
M0 2 A VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS B 2 VPW nch L=4e-08 W=1.2e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=3.1e-07 
M3 7 A 2 VNW pch L=4e-08 W=2.95e-07 
M4 VDD B 7 VNW pch L=4e-08 W=2.95e-07 
M5 Y 2 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X1P4B_A9TR Y VDD VNW VPW VSS A B
M0 2 A VSS VPW nch L=4e-08 W=1.35e-07 
M1 VSS B 2 VPW nch L=4e-08 W=1.35e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS 2 Y VPW nch L=4e-08 W=1.6e-07 
M4 7 A 2 VNW pch L=4e-08 W=4e-07 
M5 VDD B 7 VNW pch L=4e-08 W=4e-07 
M6 Y 2 VDD VNW pch L=4e-08 W=2.85e-07 
M7 VDD 2 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OR2_X1P4M_A9TR Y VDD VNW VPW VSS A B
M0 2 A VSS VPW nch L=4e-08 W=1.5e-07 
M1 VSS B 2 VPW nch L=4e-08 W=1.5e-07 
M2 Y 2 VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS 2 Y VPW nch L=4e-08 W=2.2e-07 
M4 7 A 2 VNW pch L=4e-08 W=3.7e-07 
M5 VDD B 7 VNW pch L=4e-08 W=3.7e-07 
M6 Y 2 VDD VNW pch L=4e-08 W=2.85e-07 
M7 VDD 2 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OR2_X2B_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=2.15e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.15e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=2.25e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=2.25e-07 
M4 7 B VDD VNW pch L=4e-08 W=3.25e-07 
M5 3 A 7 VNW pch L=4e-08 W=3.25e-07 
M6 8 A 3 VNW pch L=4e-08 W=3.25e-07 
M7 VDD B 8 VNW pch L=4e-08 W=3.25e-07 
M8 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M9 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X2M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.2e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M4 7 B VDD VNW pch L=4e-08 W=2.7e-07 
M5 3 A 7 VNW pch L=4e-08 W=2.7e-07 
M6 8 A 3 VNW pch L=4e-08 W=2.7e-07 
M7 VDD B 8 VNW pch L=4e-08 W=2.7e-07 
M8 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M9 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X3B_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=2.95e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.95e-07 
M2 VSS 3 Y VPW nch L=4e-08 W=3.4e-07 
M3 Y 3 VSS VPW nch L=4e-08 W=3.4e-07 
M4 7 B VDD VNW pch L=4e-08 W=4e-07 
M5 3 A 7 VNW pch L=4e-08 W=4e-07 
M6 8 A 3 VNW pch L=4e-08 W=4e-07 
M7 VDD B 8 VNW pch L=4e-08 W=4e-07 
M8 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M9 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M10 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X3M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS B 3 VPW nch L=4e-08 W=3.1e-07 
M2 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M4 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M5 7 B VDD VNW pch L=4e-08 W=3.8e-07 
M6 3 A 7 VNW pch L=4e-08 W=3.8e-07 
M7 8 A 3 VNW pch L=4e-08 W=3.8e-07 
M8 VDD B 8 VNW pch L=4e-08 W=3.8e-07 
M9 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M10 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M11 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X4B_A9TR Y VDD VNW VPW VSS A B
M0 1 B VSS VPW nch L=4e-08 W=2e-07 
M1 VSS A 1 VPW nch L=4e-08 W=2e-07 
M2 1 A VSS VPW nch L=4e-08 W=2e-07 
M3 VSS B 1 VPW nch L=4e-08 W=2e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=3e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=3e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=3e-07 
M7 7 A 1 VNW pch L=4e-08 W=4e-07 
M8 VDD B 7 VNW pch L=4e-08 W=4e-07 
M9 8 B VDD VNW pch L=4e-08 W=4e-07 
M10 1 A 8 VNW pch L=4e-08 W=4e-07 
M11 9 A 1 VNW pch L=4e-08 W=4e-07 
M12 VDD B 9 VNW pch L=4e-08 W=4e-07 
M13 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M14 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M15 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M16 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X4M_A9TR Y VDD VNW VPW VSS A B
M0 1 B VSS VPW nch L=4e-08 W=2.1e-07 
M1 VSS A 1 VPW nch L=4e-08 W=2.1e-07 
M2 1 A VSS VPW nch L=4e-08 W=2.1e-07 
M3 VSS B 1 VPW nch L=4e-08 W=2.1e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M5 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M8 7 A 1 VNW pch L=4e-08 W=3.5e-07 
M9 VDD B 7 VNW pch L=4e-08 W=3.5e-07 
M10 8 B VDD VNW pch L=4e-08 W=3.5e-07 
M11 1 A 8 VNW pch L=4e-08 W=3.5e-07 
M12 9 A 1 VNW pch L=4e-08 W=3.5e-07 
M13 VDD B 9 VNW pch L=4e-08 W=3.5e-07 
M14 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M16 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M17 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X6B_A9TR Y VDD VNW VPW VSS A B
M0 1 B VSS VPW nch L=4e-08 W=3e-07 
M1 VSS A 1 VPW nch L=4e-08 W=3e-07 
M2 1 A VSS VPW nch L=4e-08 W=3e-07 
M3 VSS B 1 VPW nch L=4e-08 W=3e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=3.35e-07 
M5 Y 1 VSS VPW nch L=4e-08 W=3.35e-07 
M6 VSS 1 Y VPW nch L=4e-08 W=3.35e-07 
M7 Y 1 VSS VPW nch L=4e-08 W=3.35e-07 
M8 7 A 1 VNW pch L=4e-08 W=3.6e-07 
M9 VDD B 7 VNW pch L=4e-08 W=3.6e-07 
M10 8 B VDD VNW pch L=4e-08 W=3.6e-07 
M11 1 A 8 VNW pch L=4e-08 W=3.6e-07 
M12 9 A 1 VNW pch L=4e-08 W=3.6e-07 
M13 VDD B 9 VNW pch L=4e-08 W=3.6e-07 
M14 10 B VDD VNW pch L=4e-08 W=3.6e-07 
M15 1 A 10 VNW pch L=4e-08 W=3.6e-07 
M16 11 A 1 VNW pch L=4e-08 W=3.6e-07 
M17 VDD B 11 VNW pch L=4e-08 W=3.6e-07 
M18 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M20 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M22 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X6M_A9TR Y VDD VNW VPW VSS A B
M0 2 B VSS VPW nch L=4e-08 W=3.1e-07 
M1 VSS A 2 VPW nch L=4e-08 W=3.1e-07 
M2 2 A VSS VPW nch L=4e-08 W=3.1e-07 
M3 VSS B 2 VPW nch L=4e-08 W=3.1e-07 
M4 Y 2 VSS VPW nch L=4e-08 W=3.75e-07 
M5 VSS 2 Y VPW nch L=4e-08 W=3.75e-07 
M6 Y 2 VSS VPW nch L=4e-08 W=3.75e-07 
M7 VSS 2 Y VPW nch L=4e-08 W=3.75e-07 
M8 Y 2 VSS VPW nch L=4e-08 W=3.75e-07 
M9 7 B VDD VNW pch L=4e-08 W=3.85e-07 
M10 2 A 7 VNW pch L=4e-08 W=3.85e-07 
M11 8 A 2 VNW pch L=4e-08 W=3.85e-07 
M12 VDD B 8 VNW pch L=4e-08 W=3.85e-07 
M13 9 B VDD VNW pch L=4e-08 W=3.85e-07 
M14 2 A 9 VNW pch L=4e-08 W=3.85e-07 
M15 10 A 2 VNW pch L=4e-08 W=3.85e-07 
M16 VDD B 10 VNW pch L=4e-08 W=3.85e-07 
M17 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M19 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M21 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 2 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X8B_A9TR Y VDD VNW VPW VSS A B
M0 2 B VSS VPW nch L=4e-08 W=4e-07 
M1 VSS A 2 VPW nch L=4e-08 W=4e-07 
M2 2 A VSS VPW nch L=4e-08 W=4e-07 
M3 VSS B 2 VPW nch L=4e-08 W=4e-07 
M4 Y 2 VSS VPW nch L=4e-08 W=4e-07 
M5 VSS 2 Y VPW nch L=4e-08 W=4e-07 
M6 Y 2 VSS VPW nch L=4e-08 W=4e-07 
M7 7 B VDD VNW pch L=4e-08 W=4e-07 
M8 2 A 7 VNW pch L=4e-08 W=4e-07 
M9 8 A 2 VNW pch L=4e-08 W=4e-07 
M10 VDD B 8 VNW pch L=4e-08 W=4e-07 
M11 9 B VDD VNW pch L=4e-08 W=4e-07 
M12 2 A 9 VNW pch L=4e-08 W=4e-07 
M13 10 A 2 VNW pch L=4e-08 W=4e-07 
M14 VDD B 10 VNW pch L=4e-08 W=4e-07 
M15 11 B VDD VNW pch L=4e-08 W=4e-07 
M16 2 A 11 VNW pch L=4e-08 W=4e-07 
M17 12 A 2 VNW pch L=4e-08 W=4e-07 
M18 VDD B 12 VNW pch L=4e-08 W=4e-07 
M19 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M20 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M21 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M23 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD 2 Y VNW pch L=4e-08 W=4e-07 
M25 Y 2 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 2 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR2_X8M_A9TR Y VDD VNW VPW VSS A B
M0 1 B VSS VPW nch L=4e-08 W=4e-07 
M1 VSS A 1 VPW nch L=4e-08 W=4e-07 
M2 1 A VSS VPW nch L=4e-08 W=4e-07 
M3 VSS B 1 VPW nch L=4e-08 W=4e-07 
M4 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M5 VSS 1 Y VPW nch L=4e-08 W=3.55e-07 
M6 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M7 VSS 1 Y VPW nch L=4e-08 W=3.55e-07 
M8 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M9 VSS 1 Y VPW nch L=4e-08 W=3.55e-07 
M10 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M11 7 A 1 VNW pch L=4e-08 W=4e-07 
M12 VDD B 7 VNW pch L=4e-08 W=4e-07 
M13 8 B VDD VNW pch L=4e-08 W=4e-07 
M14 1 A 8 VNW pch L=4e-08 W=4e-07 
M15 9 A 1 VNW pch L=4e-08 W=4e-07 
M16 VDD B 9 VNW pch L=4e-08 W=4e-07 
M17 10 B VDD VNW pch L=4e-08 W=4e-07 
M18 1 A 10 VNW pch L=4e-08 W=4e-07 
M19 11 A 1 VNW pch L=4e-08 W=4e-07 
M20 VDD B 11 VNW pch L=4e-08 W=4e-07 
M21 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M22 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M23 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M24 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M25 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M27 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR3_X0P5M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 1 B VSS VPW nch L=4e-08 W=1.2e-07 
M2 VSS C 1 VPW nch L=4e-08 W=1.2e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=1.55e-07 
M4 8 A 1 VNW pch L=4e-08 W=4e-07 
M5 9 B 8 VNW pch L=4e-08 W=4e-07 
M6 VDD C 9 VNW pch L=4e-08 W=4e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=2e-07 
.ENDS


.SUBCKT OR3_X0P7M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS A 1 VPW nch L=4e-08 W=1.2e-07 
M1 1 B VSS VPW nch L=4e-08 W=1.2e-07 
M2 VSS C 1 VPW nch L=4e-08 W=1.2e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=2.2e-07 
M4 8 A 1 VNW pch L=4e-08 W=4e-07 
M5 9 B 8 VNW pch L=4e-08 W=4e-07 
M6 VDD C 9 VNW pch L=4e-08 W=4e-07 
M7 Y 1 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OR3_X1M_A9TR Y VDD VNW VPW VSS A B C
M0 4 C VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS B 4 VPW nch L=4e-08 W=1.6e-07 
M2 4 A VSS VPW nch L=4e-08 W=1.6e-07 
M3 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VDD C 1 VNW pch L=4e-08 W=2.9e-07 
M5 1 C VDD VNW pch L=4e-08 W=2.9e-07 
M6 9 B 1 VNW pch L=4e-08 W=2.9e-07 
M7 4 A 9 VNW pch L=4e-08 W=2.9e-07 
M8 10 A 4 VNW pch L=4e-08 W=2.9e-07 
M9 1 B 10 VNW pch L=4e-08 W=2.9e-07 
M10 Y 4 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR3_X1P4M_A9TR Y VDD VNW VPW VSS A B C
M0 4 C VSS VPW nch L=4e-08 W=2e-07 
M1 VSS B 4 VPW nch L=4e-08 W=2e-07 
M2 4 A VSS VPW nch L=4e-08 W=2e-07 
M3 Y 4 VSS VPW nch L=4e-08 W=2.2e-07 
M4 VSS 4 Y VPW nch L=4e-08 W=2.2e-07 
M5 VDD C 1 VNW pch L=4e-08 W=3.75e-07 
M6 1 C VDD VNW pch L=4e-08 W=3.75e-07 
M7 9 B 1 VNW pch L=4e-08 W=3.75e-07 
M8 4 A 9 VNW pch L=4e-08 W=3.75e-07 
M9 10 A 4 VNW pch L=4e-08 W=3.75e-07 
M10 1 B 10 VNW pch L=4e-08 W=3.75e-07 
M11 Y 4 VDD VNW pch L=4e-08 W=2.85e-07 
M12 VDD 4 Y VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT OR3_X2M_A9TR Y VDD VNW VPW VSS A B C
M0 1 A VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS B 1 VPW nch L=4e-08 W=2.85e-07 
M2 1 C VSS VPW nch L=4e-08 W=2.85e-07 
M3 Y 1 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS 1 Y VPW nch L=4e-08 W=3.1e-07 
M5 9 A 1 VNW pch L=4e-08 W=3.45e-07 
M6 2 B 9 VNW pch L=4e-08 W=3.45e-07 
M7 10 B 2 VNW pch L=4e-08 W=3.45e-07 
M8 1 A 10 VNW pch L=4e-08 W=3.45e-07 
M9 11 A 1 VNW pch L=4e-08 W=3.45e-07 
M10 2 B 11 VNW pch L=4e-08 W=3.45e-07 
M11 VDD C 2 VNW pch L=4e-08 W=3.45e-07 
M12 2 C VDD VNW pch L=4e-08 W=3.45e-07 
M13 VDD C 2 VNW pch L=4e-08 W=3.45e-07 
M14 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M15 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR3_X3M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 3 VPW nch L=4e-08 W=4e-07 
M1 3 B VSS VPW nch L=4e-08 W=4e-07 
M2 VSS A 3 VPW nch L=4e-08 W=4e-07 
M3 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M5 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M6 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M7 1 C VDD VNW pch L=4e-08 W=3.8e-07 
M8 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M9 1 C VDD VNW pch L=4e-08 W=3.8e-07 
M10 9 B 1 VNW pch L=4e-08 W=3.8e-07 
M11 3 A 9 VNW pch L=4e-08 W=3.8e-07 
M12 10 A 3 VNW pch L=4e-08 W=3.8e-07 
M13 1 B 10 VNW pch L=4e-08 W=3.8e-07 
M14 11 B 1 VNW pch L=4e-08 W=3.8e-07 
M15 3 A 11 VNW pch L=4e-08 W=3.8e-07 
M16 12 A 3 VNW pch L=4e-08 W=3.8e-07 
M17 1 B 12 VNW pch L=4e-08 W=3.8e-07 
M18 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M19 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M20 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR3_X4M_A9TR Y VDD VNW VPW VSS A B C
M0 4 C VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS C 4 VPW nch L=4e-08 W=2.85e-07 
M2 4 B VSS VPW nch L=4e-08 W=2.85e-07 
M3 VSS A 4 VPW nch L=4e-08 W=2.85e-07 
M4 4 A VSS VPW nch L=4e-08 W=2.85e-07 
M5 VSS B 4 VPW nch L=4e-08 W=2.85e-07 
M6 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M8 Y 4 VSS VPW nch L=4e-08 W=3.1e-07 
M9 VSS 4 Y VPW nch L=4e-08 W=3.1e-07 
M10 VDD C 1 VNW pch L=4e-08 W=3.6e-07 
M11 1 C VDD VNW pch L=4e-08 W=3.6e-07 
M12 VDD C 1 VNW pch L=4e-08 W=3.6e-07 
M13 1 C VDD VNW pch L=4e-08 W=3.6e-07 
M14 VDD C 1 VNW pch L=4e-08 W=3.6e-07 
M15 1 C VDD VNW pch L=4e-08 W=3.6e-07 
M16 9 B 1 VNW pch L=4e-08 W=3.6e-07 
M17 4 A 9 VNW pch L=4e-08 W=3.6e-07 
M18 10 A 4 VNW pch L=4e-08 W=3.6e-07 
M19 1 B 10 VNW pch L=4e-08 W=3.6e-07 
M20 11 B 1 VNW pch L=4e-08 W=3.6e-07 
M21 4 A 11 VNW pch L=4e-08 W=3.6e-07 
M22 12 A 4 VNW pch L=4e-08 W=3.6e-07 
M23 1 B 12 VNW pch L=4e-08 W=3.6e-07 
M24 13 B 1 VNW pch L=4e-08 W=3.6e-07 
M25 4 A 13 VNW pch L=4e-08 W=3.6e-07 
M26 14 A 4 VNW pch L=4e-08 W=3.6e-07 
M27 1 B 14 VNW pch L=4e-08 W=3.6e-07 
M28 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 4 Y VNW pch L=4e-08 W=4e-07 
M30 Y 4 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 4 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR3_X6M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 3 VPW nch L=4e-08 W=2.8e-07 
M1 3 C VSS VPW nch L=4e-08 W=2.8e-07 
M2 VSS C 3 VPW nch L=4e-08 W=2.8e-07 
M3 3 B VSS VPW nch L=4e-08 W=2.8e-07 
M4 VSS A 3 VPW nch L=4e-08 W=2.8e-07 
M5 3 A VSS VPW nch L=4e-08 W=2.8e-07 
M6 VSS B 3 VPW nch L=4e-08 W=2.8e-07 
M7 3 B VSS VPW nch L=4e-08 W=2.8e-07 
M8 VSS A 3 VPW nch L=4e-08 W=2.8e-07 
M9 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M11 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M13 Y 3 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 3 Y VPW nch L=4e-08 W=3.1e-07 
M15 VDD C 1 VNW pch L=4e-08 W=3.95e-07 
M16 1 C VDD VNW pch L=4e-08 W=3.95e-07 
M17 VDD C 1 VNW pch L=4e-08 W=3.95e-07 
M18 1 C VDD VNW pch L=4e-08 W=3.95e-07 
M19 VDD C 1 VNW pch L=4e-08 W=3.95e-07 
M20 1 C VDD VNW pch L=4e-08 W=3.95e-07 
M21 VDD C 1 VNW pch L=4e-08 W=3.95e-07 
M22 1 C VDD VNW pch L=4e-08 W=3.95e-07 
M23 9 B 1 VNW pch L=4e-08 W=3.95e-07 
M24 3 A 9 VNW pch L=4e-08 W=3.95e-07 
M25 10 A 3 VNW pch L=4e-08 W=3.95e-07 
M26 1 B 10 VNW pch L=4e-08 W=3.95e-07 
M27 11 B 1 VNW pch L=4e-08 W=3.95e-07 
M28 3 A 11 VNW pch L=4e-08 W=3.95e-07 
M29 12 A 3 VNW pch L=4e-08 W=3.95e-07 
M30 1 B 12 VNW pch L=4e-08 W=3.95e-07 
M31 13 B 1 VNW pch L=4e-08 W=3.95e-07 
M32 3 A 13 VNW pch L=4e-08 W=3.95e-07 
M33 14 A 3 VNW pch L=4e-08 W=3.95e-07 
M34 1 B 14 VNW pch L=4e-08 W=3.95e-07 
M35 15 B 1 VNW pch L=4e-08 W=3.95e-07 
M36 3 A 15 VNW pch L=4e-08 W=3.95e-07 
M37 16 A 3 VNW pch L=4e-08 W=3.95e-07 
M38 1 B 16 VNW pch L=4e-08 W=3.95e-07 
M39 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M41 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M42 VDD 3 Y VNW pch L=4e-08 W=4e-07 
M43 Y 3 VDD VNW pch L=4e-08 W=4e-07 
M44 VDD 3 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR3_X8M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS A 1 VPW nch L=4e-08 W=3.85e-07 
M1 1 B VSS VPW nch L=4e-08 W=3.85e-07 
M2 VSS B 1 VPW nch L=4e-08 W=3.85e-07 
M3 1 A VSS VPW nch L=4e-08 W=3.85e-07 
M4 VSS A 1 VPW nch L=4e-08 W=3.85e-07 
M5 1 B VSS VPW nch L=4e-08 W=3.85e-07 
M6 VSS C 1 VPW nch L=4e-08 W=3.85e-07 
M7 1 C VSS VPW nch L=4e-08 W=3.85e-07 
M8 VSS C 1 VPW nch L=4e-08 W=3.85e-07 
M9 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M10 VSS 1 Y VPW nch L=4e-08 W=3.55e-07 
M11 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M12 VSS 1 Y VPW nch L=4e-08 W=3.55e-07 
M13 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M14 VSS 1 Y VPW nch L=4e-08 W=3.55e-07 
M15 Y 1 VSS VPW nch L=4e-08 W=3.55e-07 
M16 9 A 1 VNW pch L=4e-08 W=3.9e-07 
M17 2 B 9 VNW pch L=4e-08 W=3.9e-07 
M18 10 B 2 VNW pch L=4e-08 W=3.9e-07 
M19 1 A 10 VNW pch L=4e-08 W=3.9e-07 
M20 11 A 1 VNW pch L=4e-08 W=3.9e-07 
M21 2 B 11 VNW pch L=4e-08 W=3.9e-07 
M22 12 B 2 VNW pch L=4e-08 W=3.9e-07 
M23 1 A 12 VNW pch L=4e-08 W=3.9e-07 
M24 13 A 1 VNW pch L=4e-08 W=3.9e-07 
M25 2 B 13 VNW pch L=4e-08 W=3.9e-07 
M26 14 B 2 VNW pch L=4e-08 W=3.9e-07 
M27 1 A 14 VNW pch L=4e-08 W=3.9e-07 
M28 15 A 1 VNW pch L=4e-08 W=3.9e-07 
M29 2 B 15 VNW pch L=4e-08 W=3.9e-07 
M30 16 B 2 VNW pch L=4e-08 W=3.9e-07 
M31 1 A 16 VNW pch L=4e-08 W=3.9e-07 
M32 17 A 1 VNW pch L=4e-08 W=3.9e-07 
M33 2 B 17 VNW pch L=4e-08 W=3.9e-07 
M34 18 B 2 VNW pch L=4e-08 W=3.9e-07 
M35 1 A 18 VNW pch L=4e-08 W=3.9e-07 
M36 19 A 1 VNW pch L=4e-08 W=3.9e-07 
M37 2 B 19 VNW pch L=4e-08 W=3.9e-07 
M38 VDD C 2 VNW pch L=4e-08 W=3.9e-07 
M39 2 C VDD VNW pch L=4e-08 W=3.9e-07 
M40 VDD C 2 VNW pch L=4e-08 W=3.9e-07 
M41 2 C VDD VNW pch L=4e-08 W=3.9e-07 
M42 VDD C 2 VNW pch L=4e-08 W=3.9e-07 
M43 2 C VDD VNW pch L=4e-08 W=3.9e-07 
M44 VDD C 2 VNW pch L=4e-08 W=3.9e-07 
M45 2 C VDD VNW pch L=4e-08 W=3.9e-07 
M46 VDD C 2 VNW pch L=4e-08 W=3.9e-07 
M47 2 C VDD VNW pch L=4e-08 W=3.9e-07 
M48 VDD C 2 VNW pch L=4e-08 W=3.9e-07 
M49 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M50 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M51 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M52 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M53 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M54 VDD 1 Y VNW pch L=4e-08 W=4e-07 
M55 Y 1 VDD VNW pch L=4e-08 W=4e-07 
M56 VDD 1 Y VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR4_X0P5M_A9TR Y VDD VNW VPW VSS A B C D
M0 2 C VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS D 2 VPW nch L=4e-08 W=1.2e-07 
M2 12 2 VSS VPW nch L=4e-08 W=2e-07 
M3 Y 5 12 VPW nch L=4e-08 W=2e-07 
M4 5 A VSS VPW nch L=4e-08 W=1.2e-07 
M5 VSS B 5 VPW nch L=4e-08 W=1.2e-07 
M6 10 C 2 VNW pch L=4e-08 W=2.95e-07 
M7 VDD D 10 VNW pch L=4e-08 W=2.95e-07 
M8 Y 2 VDD VNW pch L=4e-08 W=1.7e-07 
M9 VDD 5 Y VNW pch L=4e-08 W=1.7e-07 
M10 11 A 5 VNW pch L=4e-08 W=2.95e-07 
M11 VDD B 11 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT OR4_X0P7M_A9TR Y VDD VNW VPW VSS A B C D
M0 2 C VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS D 2 VPW nch L=4e-08 W=1.2e-07 
M2 12 2 VSS VPW nch L=4e-08 W=2.85e-07 
M3 Y 5 12 VPW nch L=4e-08 W=2.85e-07 
M4 5 A VSS VPW nch L=4e-08 W=1.2e-07 
M5 VSS B 5 VPW nch L=4e-08 W=1.2e-07 
M6 10 C 2 VNW pch L=4e-08 W=2.95e-07 
M7 VDD D 10 VNW pch L=4e-08 W=2.95e-07 
M8 Y 2 VDD VNW pch L=4e-08 W=2.45e-07 
M9 VDD 5 Y VNW pch L=4e-08 W=2.45e-07 
M10 11 A 5 VNW pch L=4e-08 W=2.95e-07 
M11 VDD B 11 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT OR4_X1M_A9TR Y VDD VNW VPW VSS A B C D
M0 2 C VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS D 2 VPW nch L=4e-08 W=1.2e-07 
M2 12 2 VSS VPW nch L=4e-08 W=4e-07 
M3 Y 5 12 VPW nch L=4e-08 W=4e-07 
M4 5 A VSS VPW nch L=4e-08 W=1.2e-07 
M5 VSS B 5 VPW nch L=4e-08 W=1.2e-07 
M6 10 C 2 VNW pch L=4e-08 W=2.95e-07 
M7 VDD D 10 VNW pch L=4e-08 W=2.95e-07 
M8 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M9 VDD 5 Y VNW pch L=4e-08 W=3.45e-07 
M10 11 A 5 VNW pch L=4e-08 W=2.95e-07 
M11 VDD B 11 VNW pch L=4e-08 W=2.95e-07 
.ENDS


.SUBCKT OR4_X1P4M_A9TR Y VDD VNW VPW VSS A B C D
M0 2 A VSS VPW nch L=4e-08 W=1.55e-07 
M1 VSS B 2 VPW nch L=4e-08 W=1.55e-07 
M2 12 5 VSS VPW nch L=4e-08 W=2.85e-07 
M3 Y 2 12 VPW nch L=4e-08 W=2.85e-07 
M4 13 2 Y VPW nch L=4e-08 W=2.85e-07 
M5 VSS 5 13 VPW nch L=4e-08 W=2.85e-07 
M6 5 D VSS VPW nch L=4e-08 W=1.55e-07 
M7 VSS C 5 VPW nch L=4e-08 W=1.55e-07 
M8 10 A 2 VNW pch L=4e-08 W=3.85e-07 
M9 VDD B 10 VNW pch L=4e-08 W=3.85e-07 
M10 Y 5 VDD VNW pch L=4e-08 W=2.45e-07 
M11 VDD 2 Y VNW pch L=4e-08 W=2.45e-07 
M12 Y 2 VDD VNW pch L=4e-08 W=2.45e-07 
M13 VDD 5 Y VNW pch L=4e-08 W=2.45e-07 
M14 11 D VDD VNW pch L=4e-08 W=3.85e-07 
M15 5 C 11 VNW pch L=4e-08 W=3.85e-07 
.ENDS


.SUBCKT OR4_X2M_A9TR Y VDD VNW VPW VSS A B C D
M0 3 C VSS VPW nch L=4e-08 W=2.3e-07 
M1 VSS D 3 VPW nch L=4e-08 W=2.3e-07 
M2 VSS 3 4 VPW nch L=4e-08 W=4e-07 
M3 4 3 VSS VPW nch L=4e-08 W=4e-07 
M4 Y 6 4 VPW nch L=4e-08 W=4e-07 
M5 4 6 Y VPW nch L=4e-08 W=4e-07 
M6 6 B VSS VPW nch L=4e-08 W=2.3e-07 
M7 VSS A 6 VPW nch L=4e-08 W=2.3e-07 
M8 11 D VDD VNW pch L=4e-08 W=2.8e-07 
M9 3 C 11 VNW pch L=4e-08 W=2.8e-07 
M10 12 C 3 VNW pch L=4e-08 W=2.8e-07 
M11 VDD D 12 VNW pch L=4e-08 W=2.8e-07 
M12 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M13 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M14 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M15 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M16 13 B VDD VNW pch L=4e-08 W=2.8e-07 
M17 6 A 13 VNW pch L=4e-08 W=2.8e-07 
M18 14 A 6 VNW pch L=4e-08 W=2.8e-07 
M19 VDD B 14 VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT OR4_X3M_A9TR Y VDD VNW VPW VSS A B C D
M0 3 C VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS D 3 VPW nch L=4e-08 W=3.2e-07 
M2 4 3 VSS VPW nch L=4e-08 W=4e-07 
M3 VSS 3 4 VPW nch L=4e-08 W=4e-07 
M4 4 3 VSS VPW nch L=4e-08 W=4e-07 
M5 Y 6 4 VPW nch L=4e-08 W=4e-07 
M6 4 6 Y VPW nch L=4e-08 W=4e-07 
M7 Y 6 4 VPW nch L=4e-08 W=4e-07 
M8 6 B VSS VPW nch L=4e-08 W=3.2e-07 
M9 VSS A 6 VPW nch L=4e-08 W=3.2e-07 
M10 11 D VDD VNW pch L=4e-08 W=3.95e-07 
M11 3 C 11 VNW pch L=4e-08 W=3.95e-07 
M12 12 C 3 VNW pch L=4e-08 W=3.95e-07 
M13 VDD D 12 VNW pch L=4e-08 W=3.95e-07 
M14 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M15 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M16 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M17 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M18 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M19 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M20 13 B VDD VNW pch L=4e-08 W=3.95e-07 
M21 6 A 13 VNW pch L=4e-08 W=3.95e-07 
M22 14 A 6 VNW pch L=4e-08 W=3.95e-07 
M23 VDD B 14 VNW pch L=4e-08 W=3.95e-07 
.ENDS


.SUBCKT OR4_X4M_A9TR Y VDD VNW VPW VSS A B C D
M0 3 C VSS VPW nch L=4e-08 W=2.2e-07 
M1 VSS D 3 VPW nch L=4e-08 W=2.2e-07 
M2 3 D VSS VPW nch L=4e-08 W=2.2e-07 
M3 VSS C 3 VPW nch L=4e-08 W=2.2e-07 
M4 VSS 3 4 VPW nch L=4e-08 W=4e-07 
M5 4 3 VSS VPW nch L=4e-08 W=4e-07 
M6 VSS 3 4 VPW nch L=4e-08 W=4e-07 
M7 4 3 VSS VPW nch L=4e-08 W=4e-07 
M8 Y 6 4 VPW nch L=4e-08 W=4e-07 
M9 4 6 Y VPW nch L=4e-08 W=4e-07 
M10 Y 6 4 VPW nch L=4e-08 W=4e-07 
M11 4 6 Y VPW nch L=4e-08 W=4e-07 
M12 6 A VSS VPW nch L=4e-08 W=2.2e-07 
M13 VSS B 6 VPW nch L=4e-08 W=2.2e-07 
M14 6 B VSS VPW nch L=4e-08 W=2.2e-07 
M15 VSS A 6 VPW nch L=4e-08 W=2.2e-07 
M16 11 D VDD VNW pch L=4e-08 W=3.65e-07 
M17 3 C 11 VNW pch L=4e-08 W=3.65e-07 
M18 12 C 3 VNW pch L=4e-08 W=3.65e-07 
M19 VDD D 12 VNW pch L=4e-08 W=3.65e-07 
M20 13 D VDD VNW pch L=4e-08 W=3.65e-07 
M21 3 C 13 VNW pch L=4e-08 W=3.65e-07 
M22 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M23 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M24 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M25 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M26 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M27 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M28 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M29 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M30 14 A 6 VNW pch L=4e-08 W=3.65e-07 
M31 VDD B 14 VNW pch L=4e-08 W=3.65e-07 
M32 15 B VDD VNW pch L=4e-08 W=3.65e-07 
M33 6 A 15 VNW pch L=4e-08 W=3.65e-07 
M34 16 A 6 VNW pch L=4e-08 W=3.65e-07 
M35 VDD B 16 VNW pch L=4e-08 W=3.65e-07 
.ENDS


.SUBCKT OR4_X6M_A9TR Y VDD VNW VPW VSS A B C D
M0 2 D VSS VPW nch L=4e-08 W=3.2e-07 
M1 VSS C 2 VPW nch L=4e-08 W=3.2e-07 
M2 2 C VSS VPW nch L=4e-08 W=3.2e-07 
M3 VSS D 2 VPW nch L=4e-08 W=3.2e-07 
M4 VSS 2 4 VPW nch L=4e-08 W=4e-07 
M5 4 2 VSS VPW nch L=4e-08 W=4e-07 
M6 VSS 2 4 VPW nch L=4e-08 W=4e-07 
M7 4 2 VSS VPW nch L=4e-08 W=4e-07 
M8 VSS 2 4 VPW nch L=4e-08 W=4e-07 
M9 4 2 VSS VPW nch L=4e-08 W=4e-07 
M10 Y 6 4 VPW nch L=4e-08 W=4e-07 
M11 4 6 Y VPW nch L=4e-08 W=4e-07 
M12 Y 6 4 VPW nch L=4e-08 W=4e-07 
M13 4 6 Y VPW nch L=4e-08 W=4e-07 
M14 Y 6 4 VPW nch L=4e-08 W=4e-07 
M15 4 6 Y VPW nch L=4e-08 W=4e-07 
M16 6 B VSS VPW nch L=4e-08 W=3.2e-07 
M17 VSS A 6 VPW nch L=4e-08 W=3.2e-07 
M18 6 A VSS VPW nch L=4e-08 W=3.2e-07 
M19 VSS B 6 VPW nch L=4e-08 W=3.2e-07 
M20 11 D VDD VNW pch L=4e-08 W=4e-07 
M21 2 C 11 VNW pch L=4e-08 W=4e-07 
M22 12 C 2 VNW pch L=4e-08 W=4e-07 
M23 VDD D 12 VNW pch L=4e-08 W=4e-07 
M24 13 D VDD VNW pch L=4e-08 W=4e-07 
M25 2 C 13 VNW pch L=4e-08 W=4e-07 
M26 14 C 2 VNW pch L=4e-08 W=4e-07 
M27 VDD D 14 VNW pch L=4e-08 W=4e-07 
M28 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M29 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M30 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M31 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M32 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M33 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M34 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M35 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M36 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M37 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M38 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M39 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M40 15 B VDD VNW pch L=4e-08 W=4e-07 
M41 6 A 15 VNW pch L=4e-08 W=4e-07 
M42 16 A 6 VNW pch L=4e-08 W=4e-07 
M43 VDD B 16 VNW pch L=4e-08 W=4e-07 
M44 17 B VDD VNW pch L=4e-08 W=4e-07 
M45 6 A 17 VNW pch L=4e-08 W=4e-07 
M46 18 A 6 VNW pch L=4e-08 W=4e-07 
M47 VDD B 18 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR4_X8M_A9TR Y VDD VNW VPW VSS A B C D
M0 2 C VSS VPW nch L=4e-08 W=3e-07 
M1 VSS D 2 VPW nch L=4e-08 W=3e-07 
M2 2 D VSS VPW nch L=4e-08 W=3e-07 
M3 VSS C 2 VPW nch L=4e-08 W=3e-07 
M4 2 C VSS VPW nch L=4e-08 W=3e-07 
M5 VSS D 2 VPW nch L=4e-08 W=3e-07 
M6 VSS 2 4 VPW nch L=4e-08 W=4e-07 
M7 4 2 VSS VPW nch L=4e-08 W=4e-07 
M8 VSS 2 4 VPW nch L=4e-08 W=4e-07 
M9 4 2 VSS VPW nch L=4e-08 W=4e-07 
M10 VSS 2 4 VPW nch L=4e-08 W=4e-07 
M11 4 2 VSS VPW nch L=4e-08 W=4e-07 
M12 VSS 2 4 VPW nch L=4e-08 W=4e-07 
M13 4 2 VSS VPW nch L=4e-08 W=4e-07 
M14 Y 6 4 VPW nch L=4e-08 W=4e-07 
M15 4 6 Y VPW nch L=4e-08 W=4e-07 
M16 Y 6 4 VPW nch L=4e-08 W=4e-07 
M17 4 6 Y VPW nch L=4e-08 W=4e-07 
M18 Y 6 4 VPW nch L=4e-08 W=4e-07 
M19 4 6 Y VPW nch L=4e-08 W=4e-07 
M20 Y 6 4 VPW nch L=4e-08 W=4e-07 
M21 4 6 Y VPW nch L=4e-08 W=4e-07 
M22 6 B VSS VPW nch L=4e-08 W=3e-07 
M23 VSS A 6 VPW nch L=4e-08 W=3e-07 
M24 6 A VSS VPW nch L=4e-08 W=3e-07 
M25 VSS B 6 VPW nch L=4e-08 W=3e-07 
M26 6 B VSS VPW nch L=4e-08 W=3e-07 
M27 VSS A 6 VPW nch L=4e-08 W=3e-07 
M28 11 D VDD VNW pch L=4e-08 W=3.65e-07 
M29 2 C 11 VNW pch L=4e-08 W=3.65e-07 
M30 12 C 2 VNW pch L=4e-08 W=3.65e-07 
M31 VDD D 12 VNW pch L=4e-08 W=3.65e-07 
M32 13 D VDD VNW pch L=4e-08 W=3.65e-07 
M33 2 C 13 VNW pch L=4e-08 W=3.65e-07 
M34 14 C 2 VNW pch L=4e-08 W=3.65e-07 
M35 VDD D 14 VNW pch L=4e-08 W=3.65e-07 
M36 15 D VDD VNW pch L=4e-08 W=3.65e-07 
M37 2 C 15 VNW pch L=4e-08 W=3.65e-07 
M38 16 C 2 VNW pch L=4e-08 W=3.65e-07 
M39 VDD D 16 VNW pch L=4e-08 W=3.65e-07 
M40 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M41 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M42 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M43 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M44 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M45 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M46 Y 2 VDD VNW pch L=4e-08 W=3.45e-07 
M47 VDD 2 Y VNW pch L=4e-08 W=3.45e-07 
M48 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M49 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M50 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M51 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M52 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M53 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M54 Y 6 VDD VNW pch L=4e-08 W=3.45e-07 
M55 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M56 17 B VDD VNW pch L=4e-08 W=3.65e-07 
M57 6 A 17 VNW pch L=4e-08 W=3.65e-07 
M58 18 A 6 VNW pch L=4e-08 W=3.65e-07 
M59 VDD B 18 VNW pch L=4e-08 W=3.65e-07 
M60 19 B VDD VNW pch L=4e-08 W=3.65e-07 
M61 6 A 19 VNW pch L=4e-08 W=3.65e-07 
M62 20 A 6 VNW pch L=4e-08 W=3.65e-07 
M63 VDD B 20 VNW pch L=4e-08 W=3.65e-07 
M64 21 B VDD VNW pch L=4e-08 W=3.65e-07 
M65 6 A 21 VNW pch L=4e-08 W=3.65e-07 
M66 22 A 6 VNW pch L=4e-08 W=3.65e-07 
M67 VDD B 22 VNW pch L=4e-08 W=3.65e-07 
.ENDS


.SUBCKT OR6_X0P5M_A9TR Y VDD VNW VPW VSS A B C D E F
M0 VSS D 1 VPW nch L=4e-08 W=1.2e-07 
M1 1 E VSS VPW nch L=4e-08 W=1.2e-07 
M2 VSS F 1 VPW nch L=4e-08 W=1.2e-07 
M3 16 1 VSS VPW nch L=4e-08 W=2e-07 
M4 Y 5 16 VPW nch L=4e-08 W=2e-07 
M5 VSS A 5 VPW nch L=4e-08 W=1.2e-07 
M6 5 B VSS VPW nch L=4e-08 W=1.2e-07 
M7 VSS C 5 VPW nch L=4e-08 W=1.2e-07 
M8 12 D 1 VNW pch L=4e-08 W=4e-07 
M9 13 E 12 VNW pch L=4e-08 W=4e-07 
M10 VDD F 13 VNW pch L=4e-08 W=4e-07 
M11 Y 1 VDD VNW pch L=4e-08 W=1.7e-07 
M12 VDD 5 Y VNW pch L=4e-08 W=1.7e-07 
M13 14 A 5 VNW pch L=4e-08 W=4e-07 
M14 15 B 14 VNW pch L=4e-08 W=4e-07 
M15 VDD C 15 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR6_X0P7M_A9TR Y VDD VNW VPW VSS A B C D E F
M0 VSS D 1 VPW nch L=4e-08 W=1.2e-07 
M1 1 E VSS VPW nch L=4e-08 W=1.2e-07 
M2 VSS F 1 VPW nch L=4e-08 W=1.2e-07 
M3 16 1 VSS VPW nch L=4e-08 W=2.85e-07 
M4 Y 5 16 VPW nch L=4e-08 W=2.85e-07 
M5 VSS A 5 VPW nch L=4e-08 W=1.2e-07 
M6 5 B VSS VPW nch L=4e-08 W=1.2e-07 
M7 VSS C 5 VPW nch L=4e-08 W=1.2e-07 
M8 12 D 1 VNW pch L=4e-08 W=4e-07 
M9 13 E 12 VNW pch L=4e-08 W=4e-07 
M10 VDD F 13 VNW pch L=4e-08 W=4e-07 
M11 Y 1 VDD VNW pch L=4e-08 W=2.45e-07 
M12 VDD 5 Y VNW pch L=4e-08 W=2.45e-07 
M13 14 A 5 VNW pch L=4e-08 W=4e-07 
M14 15 B 14 VNW pch L=4e-08 W=4e-07 
M15 VDD C 15 VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT OR6_X1M_A9TR Y VDD VNW VPW VSS A B C D E F
M0 3 F VSS VPW nch L=4e-08 W=1.6e-07 
M1 VSS E 3 VPW nch L=4e-08 W=1.6e-07 
M2 3 D VSS VPW nch L=4e-08 W=1.6e-07 
M3 VSS 3 4 VPW nch L=4e-08 W=2e-07 
M4 4 3 VSS VPW nch L=4e-08 W=2e-07 
M5 Y 6 4 VPW nch L=4e-08 W=2e-07 
M6 4 6 Y VPW nch L=4e-08 W=2e-07 
M7 VSS A 6 VPW nch L=4e-08 W=1.6e-07 
M8 6 B VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS C 6 VPW nch L=4e-08 W=1.6e-07 
M10 13 F VDD VNW pch L=4e-08 W=3e-07 
M11 14 E 13 VNW pch L=4e-08 W=3e-07 
M12 3 D 14 VNW pch L=4e-08 W=3e-07 
M13 15 D 3 VNW pch L=4e-08 W=3e-07 
M14 16 E 15 VNW pch L=4e-08 W=3e-07 
M15 VDD F 16 VNW pch L=4e-08 W=3e-07 
M16 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M17 VDD 6 Y VNW pch L=4e-08 W=3.45e-07 
M18 17 C VDD VNW pch L=4e-08 W=3e-07 
M19 18 B 17 VNW pch L=4e-08 W=3e-07 
M20 6 A 18 VNW pch L=4e-08 W=3e-07 
M21 19 A 6 VNW pch L=4e-08 W=3e-07 
M22 20 B 19 VNW pch L=4e-08 W=3e-07 
M23 VDD C 20 VNW pch L=4e-08 W=3e-07 
.ENDS


.SUBCKT OR6_X1P4M_A9TR Y VDD VNW VPW VSS A B C D E F
M0 3 F VSS VPW nch L=4e-08 W=2.1e-07 
M1 VSS E 3 VPW nch L=4e-08 W=2.1e-07 
M2 3 D VSS VPW nch L=4e-08 W=2.1e-07 
M3 VSS 3 4 VPW nch L=4e-08 W=2.85e-07 
M4 4 3 VSS VPW nch L=4e-08 W=2.85e-07 
M5 Y 6 4 VPW nch L=4e-08 W=2.85e-07 
M6 4 6 Y VPW nch L=4e-08 W=2.85e-07 
M7 VSS A 6 VPW nch L=4e-08 W=2.1e-07 
M8 6 B VSS VPW nch L=4e-08 W=2.1e-07 
M9 VSS C 6 VPW nch L=4e-08 W=2.1e-07 
M10 13 F VDD VNW pch L=4e-08 W=3.9e-07 
M11 14 E 13 VNW pch L=4e-08 W=3.9e-07 
M12 3 D 14 VNW pch L=4e-08 W=3.9e-07 
M13 15 D 3 VNW pch L=4e-08 W=3.9e-07 
M14 16 E 15 VNW pch L=4e-08 W=3.9e-07 
M15 VDD F 16 VNW pch L=4e-08 W=3.9e-07 
M16 Y 3 VDD VNW pch L=4e-08 W=2.45e-07 
M17 VDD 3 Y VNW pch L=4e-08 W=2.45e-07 
M18 Y 6 VDD VNW pch L=4e-08 W=2.45e-07 
M19 VDD 6 Y VNW pch L=4e-08 W=2.45e-07 
M20 17 C VDD VNW pch L=4e-08 W=3.9e-07 
M21 18 B 17 VNW pch L=4e-08 W=3.9e-07 
M22 6 A 18 VNW pch L=4e-08 W=3.9e-07 
M23 19 A 6 VNW pch L=4e-08 W=3.9e-07 
M24 20 B 19 VNW pch L=4e-08 W=3.9e-07 
M25 VDD C 20 VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT OR6_X2M_A9TR Y VDD VNW VPW VSS A B C D E F
M0 1 D VSS VPW nch L=4e-08 W=2.85e-07 
M1 VSS E 1 VPW nch L=4e-08 W=2.85e-07 
M2 1 F VSS VPW nch L=4e-08 W=2.85e-07 
M3 VSS 1 5 VPW nch L=4e-08 W=4e-07 
M4 5 1 VSS VPW nch L=4e-08 W=4e-07 
M5 Y 8 5 VPW nch L=4e-08 W=4e-07 
M6 5 8 Y VPW nch L=4e-08 W=4e-07 
M7 VSS C 8 VPW nch L=4e-08 W=2.85e-07 
M8 8 B VSS VPW nch L=4e-08 W=2.85e-07 
M9 VSS A 8 VPW nch L=4e-08 W=2.85e-07 
M10 15 D 1 VNW pch L=4e-08 W=3.55e-07 
M11 2 E 15 VNW pch L=4e-08 W=3.55e-07 
M12 16 E 2 VNW pch L=4e-08 W=3.55e-07 
M13 1 D 16 VNW pch L=4e-08 W=3.55e-07 
M14 17 D 1 VNW pch L=4e-08 W=3.55e-07 
M15 2 E 17 VNW pch L=4e-08 W=3.55e-07 
M16 VDD F 2 VNW pch L=4e-08 W=3.55e-07 
M17 2 F VDD VNW pch L=4e-08 W=3.55e-07 
M18 VDD F 2 VNW pch L=4e-08 W=3.55e-07 
M19 Y 1 VDD VNW pch L=4e-08 W=3.45e-07 
M20 VDD 1 Y VNW pch L=4e-08 W=3.45e-07 
M21 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M22 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M23 7 C VDD VNW pch L=4e-08 W=3.55e-07 
M24 VDD C 7 VNW pch L=4e-08 W=3.55e-07 
M25 7 C VDD VNW pch L=4e-08 W=3.55e-07 
M26 18 B 7 VNW pch L=4e-08 W=3.55e-07 
M27 8 A 18 VNW pch L=4e-08 W=3.55e-07 
M28 19 A 8 VNW pch L=4e-08 W=3.55e-07 
M29 7 B 19 VNW pch L=4e-08 W=3.55e-07 
M30 20 B 7 VNW pch L=4e-08 W=3.55e-07 
M31 8 A 20 VNW pch L=4e-08 W=3.55e-07 
.ENDS


.SUBCKT OR6_X3M_A9TR Y VDD VNW VPW VSS A B C D E F
M0 4 F VSS VPW nch L=4e-08 W=2.1e-07 
M1 VSS F 4 VPW nch L=4e-08 W=2.1e-07 
M2 4 E VSS VPW nch L=4e-08 W=2.1e-07 
M3 VSS D 4 VPW nch L=4e-08 W=2.1e-07 
M4 4 D VSS VPW nch L=4e-08 W=2.1e-07 
M5 VSS E 4 VPW nch L=4e-08 W=2.1e-07 
M6 6 4 VSS VPW nch L=4e-08 W=4e-07 
M7 VSS 4 6 VPW nch L=4e-08 W=4e-07 
M8 6 4 VSS VPW nch L=4e-08 W=4e-07 
M9 Y 8 6 VPW nch L=4e-08 W=4e-07 
M10 6 8 Y VPW nch L=4e-08 W=4e-07 
M11 Y 8 6 VPW nch L=4e-08 W=4e-07 
M12 8 B VSS VPW nch L=4e-08 W=2.1e-07 
M13 VSS A 8 VPW nch L=4e-08 W=2.1e-07 
M14 8 A VSS VPW nch L=4e-08 W=2.1e-07 
M15 VSS B 8 VPW nch L=4e-08 W=2.1e-07 
M16 8 C VSS VPW nch L=4e-08 W=2.1e-07 
M17 VSS C 8 VPW nch L=4e-08 W=2.1e-07 
M18 VDD F 1 VNW pch L=4e-08 W=3.9e-07 
M19 1 F VDD VNW pch L=4e-08 W=3.9e-07 
M20 VDD F 1 VNW pch L=4e-08 W=3.9e-07 
M21 1 F VDD VNW pch L=4e-08 W=3.9e-07 
M22 15 E 1 VNW pch L=4e-08 W=3.9e-07 
M23 4 D 15 VNW pch L=4e-08 W=3.9e-07 
M24 16 D 4 VNW pch L=4e-08 W=3.9e-07 
M25 1 E 16 VNW pch L=4e-08 W=3.9e-07 
M26 17 E 1 VNW pch L=4e-08 W=3.9e-07 
M27 4 D 17 VNW pch L=4e-08 W=3.9e-07 
M28 18 D 4 VNW pch L=4e-08 W=3.9e-07 
M29 1 E 18 VNW pch L=4e-08 W=3.9e-07 
M30 VDD 4 Y VNW pch L=4e-08 W=3.45e-07 
M31 Y 4 VDD VNW pch L=4e-08 W=3.45e-07 
M32 VDD 4 Y VNW pch L=4e-08 W=3.45e-07 
M33 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M34 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M35 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M36 19 B 7 VNW pch L=4e-08 W=3.9e-07 
M37 8 A 19 VNW pch L=4e-08 W=3.9e-07 
M38 20 A 8 VNW pch L=4e-08 W=3.9e-07 
M39 7 B 20 VNW pch L=4e-08 W=3.9e-07 
M40 21 B 7 VNW pch L=4e-08 W=3.9e-07 
M41 8 A 21 VNW pch L=4e-08 W=3.9e-07 
M42 22 A 8 VNW pch L=4e-08 W=3.9e-07 
M43 7 B 22 VNW pch L=4e-08 W=3.9e-07 
M44 VDD C 7 VNW pch L=4e-08 W=3.9e-07 
M45 7 C VDD VNW pch L=4e-08 W=3.9e-07 
M46 VDD C 7 VNW pch L=4e-08 W=3.9e-07 
M47 7 C VDD VNW pch L=4e-08 W=3.9e-07 
.ENDS


.SUBCKT OR6_X4M_A9TR Y VDD VNW VPW VSS A B C D E F
M0 4 F VSS VPW nch L=4e-08 W=3e-07 
M1 VSS F 4 VPW nch L=4e-08 W=3e-07 
M2 4 E VSS VPW nch L=4e-08 W=3e-07 
M3 VSS D 4 VPW nch L=4e-08 W=3e-07 
M4 4 D VSS VPW nch L=4e-08 W=3e-07 
M5 VSS E 4 VPW nch L=4e-08 W=3e-07 
M6 VSS 4 5 VPW nch L=4e-08 W=4e-07 
M7 5 4 VSS VPW nch L=4e-08 W=4e-07 
M8 VSS 4 5 VPW nch L=4e-08 W=4e-07 
M9 5 4 VSS VPW nch L=4e-08 W=4e-07 
M10 Y 8 5 VPW nch L=4e-08 W=4e-07 
M11 5 8 Y VPW nch L=4e-08 W=4e-07 
M12 Y 8 5 VPW nch L=4e-08 W=4e-07 
M13 5 8 Y VPW nch L=4e-08 W=4e-07 
M14 8 B VSS VPW nch L=4e-08 W=3e-07 
M15 VSS A 8 VPW nch L=4e-08 W=3e-07 
M16 8 A VSS VPW nch L=4e-08 W=3e-07 
M17 VSS B 8 VPW nch L=4e-08 W=3e-07 
M18 8 C VSS VPW nch L=4e-08 W=3e-07 
M19 VSS C 8 VPW nch L=4e-08 W=3e-07 
M20 VDD F 1 VNW pch L=4e-08 W=3.7e-07 
M21 1 F VDD VNW pch L=4e-08 W=3.7e-07 
M22 VDD F 1 VNW pch L=4e-08 W=3.7e-07 
M23 1 F VDD VNW pch L=4e-08 W=3.7e-07 
M24 VDD F 1 VNW pch L=4e-08 W=3.7e-07 
M25 1 F VDD VNW pch L=4e-08 W=3.7e-07 
M26 15 E 1 VNW pch L=4e-08 W=3.7e-07 
M27 4 D 15 VNW pch L=4e-08 W=3.7e-07 
M28 16 D 4 VNW pch L=4e-08 W=3.7e-07 
M29 1 E 16 VNW pch L=4e-08 W=3.7e-07 
M30 17 E 1 VNW pch L=4e-08 W=3.7e-07 
M31 4 D 17 VNW pch L=4e-08 W=3.7e-07 
M32 18 D 4 VNW pch L=4e-08 W=3.7e-07 
M33 1 E 18 VNW pch L=4e-08 W=3.7e-07 
M34 19 E 1 VNW pch L=4e-08 W=3.7e-07 
M35 4 D 19 VNW pch L=4e-08 W=3.7e-07 
M36 20 D 4 VNW pch L=4e-08 W=3.7e-07 
M37 1 E 20 VNW pch L=4e-08 W=3.7e-07 
M38 Y 4 VDD VNW pch L=4e-08 W=3.45e-07 
M39 VDD 4 Y VNW pch L=4e-08 W=3.45e-07 
M40 Y 4 VDD VNW pch L=4e-08 W=3.45e-07 
M41 VDD 4 Y VNW pch L=4e-08 W=3.45e-07 
M42 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M43 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M44 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M45 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M46 21 B 7 VNW pch L=4e-08 W=3.7e-07 
M47 8 A 21 VNW pch L=4e-08 W=3.7e-07 
M48 22 A 8 VNW pch L=4e-08 W=3.7e-07 
M49 7 B 22 VNW pch L=4e-08 W=3.7e-07 
M50 23 B 7 VNW pch L=4e-08 W=3.7e-07 
M51 8 A 23 VNW pch L=4e-08 W=3.7e-07 
M52 24 A 8 VNW pch L=4e-08 W=3.7e-07 
M53 7 B 24 VNW pch L=4e-08 W=3.7e-07 
M54 25 B 7 VNW pch L=4e-08 W=3.7e-07 
M55 8 A 25 VNW pch L=4e-08 W=3.7e-07 
M56 26 A 8 VNW pch L=4e-08 W=3.7e-07 
M57 7 B 26 VNW pch L=4e-08 W=3.7e-07 
M58 VDD C 7 VNW pch L=4e-08 W=3.7e-07 
M59 7 C VDD VNW pch L=4e-08 W=3.7e-07 
M60 VDD C 7 VNW pch L=4e-08 W=3.7e-07 
M61 7 C VDD VNW pch L=4e-08 W=3.7e-07 
M62 VDD C 7 VNW pch L=4e-08 W=3.7e-07 
M63 7 C VDD VNW pch L=4e-08 W=3.7e-07 
.ENDS


.SUBCKT OR6_X6M_A9TR Y VDD VNW VPW VSS A B C D E F
M0 VSS F 3 VPW nch L=4e-08 W=2.95e-07 
M1 3 F VSS VPW nch L=4e-08 W=2.95e-07 
M2 VSS F 3 VPW nch L=4e-08 W=2.95e-07 
M3 3 E VSS VPW nch L=4e-08 W=2.95e-07 
M4 VSS D 3 VPW nch L=4e-08 W=2.95e-07 
M5 3 D VSS VPW nch L=4e-08 W=2.95e-07 
M6 VSS E 3 VPW nch L=4e-08 W=2.95e-07 
M7 3 E VSS VPW nch L=4e-08 W=2.95e-07 
M8 VSS D 3 VPW nch L=4e-08 W=2.95e-07 
M9 VSS 3 5 VPW nch L=4e-08 W=4e-07 
M10 5 3 VSS VPW nch L=4e-08 W=4e-07 
M11 VSS 3 5 VPW nch L=4e-08 W=4e-07 
M12 5 3 VSS VPW nch L=4e-08 W=4e-07 
M13 VSS 3 5 VPW nch L=4e-08 W=4e-07 
M14 5 3 VSS VPW nch L=4e-08 W=4e-07 
M15 Y 8 5 VPW nch L=4e-08 W=4e-07 
M16 5 8 Y VPW nch L=4e-08 W=4e-07 
M17 Y 8 5 VPW nch L=4e-08 W=4e-07 
M18 5 8 Y VPW nch L=4e-08 W=4e-07 
M19 Y 8 5 VPW nch L=4e-08 W=4e-07 
M20 5 8 Y VPW nch L=4e-08 W=4e-07 
M21 8 A VSS VPW nch L=4e-08 W=2.95e-07 
M22 VSS B 8 VPW nch L=4e-08 W=2.95e-07 
M23 8 B VSS VPW nch L=4e-08 W=2.95e-07 
M24 VSS A 8 VPW nch L=4e-08 W=2.95e-07 
M25 8 A VSS VPW nch L=4e-08 W=2.95e-07 
M26 VSS B 8 VPW nch L=4e-08 W=2.95e-07 
M27 8 C VSS VPW nch L=4e-08 W=2.95e-07 
M28 VSS C 8 VPW nch L=4e-08 W=2.95e-07 
M29 8 C VSS VPW nch L=4e-08 W=2.95e-07 
M30 VDD F 1 VNW pch L=4e-08 W=4e-07 
M31 1 F VDD VNW pch L=4e-08 W=4e-07 
M32 VDD F 1 VNW pch L=4e-08 W=4e-07 
M33 1 F VDD VNW pch L=4e-08 W=4e-07 
M34 VDD F 1 VNW pch L=4e-08 W=4e-07 
M35 1 F VDD VNW pch L=4e-08 W=4e-07 
M36 VDD F 1 VNW pch L=4e-08 W=4e-07 
M37 1 F VDD VNW pch L=4e-08 W=4e-07 
M38 15 E 1 VNW pch L=4e-08 W=4e-07 
M39 3 D 15 VNW pch L=4e-08 W=4e-07 
M40 16 D 3 VNW pch L=4e-08 W=4e-07 
M41 1 E 16 VNW pch L=4e-08 W=4e-07 
M42 17 E 1 VNW pch L=4e-08 W=4e-07 
M43 3 D 17 VNW pch L=4e-08 W=4e-07 
M44 18 D 3 VNW pch L=4e-08 W=4e-07 
M45 1 E 18 VNW pch L=4e-08 W=4e-07 
M46 19 E 1 VNW pch L=4e-08 W=4e-07 
M47 3 D 19 VNW pch L=4e-08 W=4e-07 
M48 20 D 3 VNW pch L=4e-08 W=4e-07 
M49 1 E 20 VNW pch L=4e-08 W=4e-07 
M50 21 E 1 VNW pch L=4e-08 W=4e-07 
M51 3 D 21 VNW pch L=4e-08 W=4e-07 
M52 22 D 3 VNW pch L=4e-08 W=4e-07 
M53 1 E 22 VNW pch L=4e-08 W=4e-07 
M54 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M55 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M56 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M57 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M58 Y 3 VDD VNW pch L=4e-08 W=3.45e-07 
M59 VDD 3 Y VNW pch L=4e-08 W=3.45e-07 
M60 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M61 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M62 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M63 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M64 Y 8 VDD VNW pch L=4e-08 W=3.45e-07 
M65 VDD 8 Y VNW pch L=4e-08 W=3.45e-07 
M66 23 B 7 VNW pch L=4e-08 W=4e-07 
M67 8 A 23 VNW pch L=4e-08 W=4e-07 
M68 24 A 8 VNW pch L=4e-08 W=4e-07 
M69 7 B 24 VNW pch L=4e-08 W=4e-07 
M70 25 B 7 VNW pch L=4e-08 W=4e-07 
M71 8 A 25 VNW pch L=4e-08 W=4e-07 
M72 26 A 8 VNW pch L=4e-08 W=4e-07 
M73 7 B 26 VNW pch L=4e-08 W=4e-07 
M74 27 B 7 VNW pch L=4e-08 W=4e-07 
M75 8 A 27 VNW pch L=4e-08 W=4e-07 
M76 28 A 8 VNW pch L=4e-08 W=4e-07 
M77 7 B 28 VNW pch L=4e-08 W=4e-07 
M78 29 B 7 VNW pch L=4e-08 W=4e-07 
M79 8 A 29 VNW pch L=4e-08 W=4e-07 
M80 30 A 8 VNW pch L=4e-08 W=4e-07 
M81 7 B 30 VNW pch L=4e-08 W=4e-07 
M82 VDD C 7 VNW pch L=4e-08 W=4e-07 
M83 7 C VDD VNW pch L=4e-08 W=4e-07 
M84 VDD C 7 VNW pch L=4e-08 W=4e-07 
M85 7 C VDD VNW pch L=4e-08 W=4e-07 
M86 VDD C 7 VNW pch L=4e-08 W=4e-07 
M87 7 C VDD VNW pch L=4e-08 W=4e-07 
M88 VDD C 7 VNW pch L=4e-08 W=4e-07 
M89 7 C VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X0P5B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=1.9e-07 
M6 6 5 14 VPW nch L=4e-08 W=1.9e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=1.2e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M12 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M13 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M15 6 SEN VDD VNW pch L=4e-08 W=1.6e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.6e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.4e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT POSTICG_X0P6B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=1.9e-07 
M6 6 5 14 VPW nch L=4e-08 W=1.9e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=1.35e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M12 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M13 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M15 6 SEN VDD VNW pch L=4e-08 W=1.6e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.6e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.4e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT POSTICG_X0P7B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=1.9e-07 
M6 6 5 14 VPW nch L=4e-08 W=1.9e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=1.6e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M12 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M13 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M15 6 SEN VDD VNW pch L=4e-08 W=1.6e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.6e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.4e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT POSTICG_X0P8B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=1.9e-07 
M6 6 5 14 VPW nch L=4e-08 W=1.9e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=1.9e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M12 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M13 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M15 6 SEN VDD VNW pch L=4e-08 W=1.6e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.6e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.4e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT POSTICG_X11B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=2.6e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.6e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=3.8e-07 
M6 6 5 14 VPW nch L=4e-08 W=3.8e-07 
M7 15 6 VSS VPW nch L=4e-08 W=3.4e-07 
M8 7 CK 15 VPW nch L=4e-08 W=3.4e-07 
M9 16 CK 7 VPW nch L=4e-08 W=3.4e-07 
M10 VSS 6 16 VPW nch L=4e-08 W=3.4e-07 
M11 17 6 VSS VPW nch L=4e-08 W=3.4e-07 
M12 7 CK 17 VPW nch L=4e-08 W=3.4e-07 
M13 ECK 7 VSS VPW nch L=4e-08 W=3.55e-07 
M14 VSS 7 ECK VPW nch L=4e-08 W=3.55e-07 
M15 ECK 7 VSS VPW nch L=4e-08 W=3.55e-07 
M16 VSS 7 ECK VPW nch L=4e-08 W=3.55e-07 
M17 ECK 7 VSS VPW nch L=4e-08 W=3.55e-07 
M18 VSS 7 ECK VPW nch L=4e-08 W=3.55e-07 
M19 ECK 7 VSS VPW nch L=4e-08 W=3.55e-07 
M20 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M21 4 E VDD VNW pch L=4e-08 W=3.3e-07 
M22 5 CK 4 VNW pch L=4e-08 W=2.6e-07 
M23 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M25 6 SEN VDD VNW pch L=4e-08 W=3.2e-07 
M26 VDD 5 6 VNW pch L=4e-08 W=3.2e-07 
M27 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M28 VDD CK 7 VNW pch L=4e-08 W=2.25e-07 
M29 7 CK VDD VNW pch L=4e-08 W=2.25e-07 
M30 VDD CK 7 VNW pch L=4e-08 W=2.25e-07 
M31 7 CK VDD VNW pch L=4e-08 W=2.25e-07 
M32 VDD CK 7 VNW pch L=4e-08 W=2.25e-07 
M33 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M35 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M37 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M39 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M41 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M42 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M43 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X13B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=2.8e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.8e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2e-07 
M6 6 5 14 VPW nch L=4e-08 W=2e-07 
M7 15 5 6 VPW nch L=4e-08 W=2e-07 
M8 VSS SEN 15 VPW nch L=4e-08 W=2e-07 
M9 16 6 VSS VPW nch L=4e-08 W=3e-07 
M10 7 CK 16 VPW nch L=4e-08 W=3e-07 
M11 17 CK 7 VPW nch L=4e-08 W=3e-07 
M12 VSS 6 17 VPW nch L=4e-08 W=3e-07 
M13 18 6 VSS VPW nch L=4e-08 W=3e-07 
M14 7 CK 18 VPW nch L=4e-08 W=3e-07 
M15 19 CK 7 VPW nch L=4e-08 W=3e-07 
M16 VSS 6 19 VPW nch L=4e-08 W=3e-07 
M17 VSS 7 ECK VPW nch L=4e-08 W=3.25e-07 
M18 ECK 7 VSS VPW nch L=4e-08 W=3.25e-07 
M19 VSS 7 ECK VPW nch L=4e-08 W=3.25e-07 
M20 ECK 7 VSS VPW nch L=4e-08 W=3.25e-07 
M21 VSS 7 ECK VPW nch L=4e-08 W=3.25e-07 
M22 ECK 7 VSS VPW nch L=4e-08 W=3.25e-07 
M23 VSS 7 ECK VPW nch L=4e-08 W=3.25e-07 
M24 ECK 7 VSS VPW nch L=4e-08 W=3.25e-07 
M25 VSS 7 ECK VPW nch L=4e-08 W=3.25e-07 
M26 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M27 4 E VDD VNW pch L=4e-08 W=3.65e-07 
M28 5 CK 4 VNW pch L=4e-08 W=2.8e-07 
M29 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M31 6 SEN VDD VNW pch L=4e-08 W=1.75e-07 
M32 VDD 5 6 VNW pch L=4e-08 W=1.75e-07 
M33 6 5 VDD VNW pch L=4e-08 W=1.75e-07 
M34 VDD SEN 6 VNW pch L=4e-08 W=1.75e-07 
M35 7 CK VDD VNW pch L=4e-08 W=2.3e-07 
M36 VDD CK 7 VNW pch L=4e-08 W=2.3e-07 
M37 7 CK VDD VNW pch L=4e-08 W=2.3e-07 
M38 VDD CK 7 VNW pch L=4e-08 W=2.3e-07 
M39 7 CK VDD VNW pch L=4e-08 W=2.3e-07 
M40 VDD CK 7 VNW pch L=4e-08 W=2.3e-07 
M41 7 6 VDD VNW pch L=4e-08 W=1.4e-07 
M42 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M43 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M44 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M45 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M46 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M47 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M48 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M49 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M50 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M51 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M52 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M53 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M54 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X16B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=3.1e-07 
M2 5 1 4 VPW nch L=4e-08 W=3.1e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2.5e-07 
M6 6 5 14 VPW nch L=4e-08 W=2.5e-07 
M7 15 5 6 VPW nch L=4e-08 W=2.5e-07 
M8 VSS SEN 15 VPW nch L=4e-08 W=2.5e-07 
M9 16 6 VSS VPW nch L=4e-08 W=3.5e-07 
M10 7 CK 16 VPW nch L=4e-08 W=3.5e-07 
M11 17 CK 7 VPW nch L=4e-08 W=3.5e-07 
M12 VSS 6 17 VPW nch L=4e-08 W=3.5e-07 
M13 18 6 VSS VPW nch L=4e-08 W=3.5e-07 
M14 7 CK 18 VPW nch L=4e-08 W=3.5e-07 
M15 19 CK 7 VPW nch L=4e-08 W=3.5e-07 
M16 VSS 6 19 VPW nch L=4e-08 W=3.5e-07 
M17 ECK 7 VSS VPW nch L=4e-08 W=3.6e-07 
M18 VSS 7 ECK VPW nch L=4e-08 W=3.6e-07 
M19 ECK 7 VSS VPW nch L=4e-08 W=3.6e-07 
M20 VSS 7 ECK VPW nch L=4e-08 W=3.6e-07 
M21 ECK 7 VSS VPW nch L=4e-08 W=3.6e-07 
M22 VSS 7 ECK VPW nch L=4e-08 W=3.6e-07 
M23 ECK 7 VSS VPW nch L=4e-08 W=3.6e-07 
M24 VSS 7 ECK VPW nch L=4e-08 W=3.6e-07 
M25 ECK 7 VSS VPW nch L=4e-08 W=3.6e-07 
M26 VSS 7 ECK VPW nch L=4e-08 W=3.6e-07 
M27 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M28 4 E VDD VNW pch L=4e-08 W=3.8e-07 
M29 5 CK 4 VNW pch L=4e-08 W=3.1e-07 
M30 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M32 6 SEN VDD VNW pch L=4e-08 W=2.15e-07 
M33 VDD 5 6 VNW pch L=4e-08 W=2.15e-07 
M34 6 5 VDD VNW pch L=4e-08 W=2.15e-07 
M35 VDD SEN 6 VNW pch L=4e-08 W=2.15e-07 
M36 7 6 VDD VNW pch L=4e-08 W=1.65e-07 
M37 VDD CK 7 VNW pch L=4e-08 W=2.35e-07 
M38 7 CK VDD VNW pch L=4e-08 W=2.35e-07 
M39 VDD CK 7 VNW pch L=4e-08 W=2.35e-07 
M40 7 CK VDD VNW pch L=4e-08 W=2.35e-07 
M41 VDD CK 7 VNW pch L=4e-08 W=2.35e-07 
M42 7 CK VDD VNW pch L=4e-08 W=2.35e-07 
M43 VDD CK 7 VNW pch L=4e-08 W=2.35e-07 
M44 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M45 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M46 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M47 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M48 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M49 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M50 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M51 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M52 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M53 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M54 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M55 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M56 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M57 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M58 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M59 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X1B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=1.9e-07 
M6 6 5 14 VPW nch L=4e-08 W=1.9e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=2.25e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M12 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M13 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M15 6 SEN VDD VNW pch L=4e-08 W=1.6e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.6e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.3e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.3e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X1P2B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=1.9e-07 
M6 6 5 14 VPW nch L=4e-08 W=1.9e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.45e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.45e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=2.7e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M12 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M13 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M15 6 SEN VDD VNW pch L=4e-08 W=1.65e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.65e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.7e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.4e-07 
M20 VDD 7 ECK VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT POSTICG_X1P4B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=1.95e-07 
M6 6 5 14 VPW nch L=4e-08 W=1.95e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.6e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.6e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=3.2e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M12 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M13 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M15 6 SEN VDD VNW pch L=4e-08 W=1.65e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.65e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.9e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.85e-07 
M20 VDD 7 ECK VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT POSTICG_X1P7B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2e-07 
M6 6 5 14 VPW nch L=4e-08 W=2e-07 
M7 15 6 VSS VPW nch L=4e-08 W=1.8e-07 
M8 7 CK 15 VPW nch L=4e-08 W=1.8e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=3.8e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M12 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M13 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M15 6 SEN VDD VNW pch L=4e-08 W=1.7e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.7e-07 
M17 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M18 VDD CK 7 VNW pch L=4e-08 W=2.1e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=3.35e-07 
M20 VDD 7 ECK VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT POSTICG_X2B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2e-07 
M6 6 5 14 VPW nch L=4e-08 W=2e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.1e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.1e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=2.25e-07 
M10 VSS 7 ECK VPW nch L=4e-08 W=2.25e-07 
M11 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M12 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M16 6 SEN VDD VNW pch L=4e-08 W=1.7e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.7e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M19 VDD CK 7 VNW pch L=4e-08 W=2.4e-07 
M20 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X2P5B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2.1e-07 
M6 6 5 14 VPW nch L=4e-08 W=2.1e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.55e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.55e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=2.85e-07 
M10 VSS 7 ECK VPW nch L=4e-08 W=2.85e-07 
M11 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M12 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M16 6 SEN VDD VNW pch L=4e-08 W=1.8e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.8e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M19 VDD CK 7 VNW pch L=4e-08 W=2.95e-07 
M20 ECK 7 VDD VNW pch L=4e-08 W=3.35e-07 
M21 VDD 7 ECK VNW pch L=4e-08 W=3.35e-07 
M22 ECK 7 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT POSTICG_X3B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2.1e-07 
M6 6 5 14 VPW nch L=4e-08 W=2.1e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.9e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.9e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=3.4e-07 
M10 VSS 7 ECK VPW nch L=4e-08 W=3.4e-07 
M11 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M12 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M16 6 SEN VDD VNW pch L=4e-08 W=1.8e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.8e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M19 VDD CK 7 VNW pch L=4e-08 W=3.4e-07 
M20 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M22 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X3P5B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2.2e-07 
M6 6 5 14 VPW nch L=4e-08 W=2.2e-07 
M7 15 6 VSS VPW nch L=4e-08 W=3.2e-07 
M8 7 CK 15 VPW nch L=4e-08 W=3.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=4e-07 
M10 VSS 7 ECK VPW nch L=4e-08 W=4e-07 
M11 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M12 4 E VDD VNW pch L=4e-08 W=1.9e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M16 6 SEN VDD VNW pch L=4e-08 W=2e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=2e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M19 VDD CK 7 VNW pch L=4e-08 W=3.65e-07 
M20 ECK 7 VDD VNW pch L=4e-08 W=3.5e-07 
M21 VDD 7 ECK VNW pch L=4e-08 W=3.5e-07 
M22 ECK 7 VDD VNW pch L=4e-08 W=3.5e-07 
M23 VDD 7 ECK VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT POSTICG_X4B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.7e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.7e-07 
M3 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 15 SEN VSS VPW nch L=4e-08 W=2.5e-07 
M6 6 5 15 VPW nch L=4e-08 W=2.5e-07 
M7 16 6 VSS VPW nch L=4e-08 W=2.05e-07 
M8 7 CK 16 VPW nch L=4e-08 W=2.05e-07 
M9 17 CK 7 VPW nch L=4e-08 W=2.05e-07 
M10 VSS 6 17 VPW nch L=4e-08 W=2.05e-07 
M11 VSS 7 ECK VPW nch L=4e-08 W=3e-07 
M12 ECK 7 VSS VPW nch L=4e-08 W=3e-07 
M13 VSS 7 ECK VPW nch L=4e-08 W=3e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M15 4 E VDD VNW pch L=4e-08 W=2.2e-07 
M16 5 CK 4 VNW pch L=4e-08 W=1.7e-07 
M17 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M18 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M19 6 SEN VDD VNW pch L=4e-08 W=2.1e-07 
M20 VDD 5 6 VNW pch L=4e-08 W=2.1e-07 
M21 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M22 7 CK VDD VNW pch L=4e-08 W=2.4e-07 
M23 VDD CK 7 VNW pch L=4e-08 W=2.4e-07 
M24 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M26 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X5B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.8e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.8e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2.6e-07 
M6 6 5 14 VPW nch L=4e-08 W=2.6e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.5e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.5e-07 
M9 16 CK 7 VPW nch L=4e-08 W=2.5e-07 
M10 VSS 6 16 VPW nch L=4e-08 W=2.5e-07 
M11 VSS 7 ECK VPW nch L=4e-08 W=3.75e-07 
M12 ECK 7 VSS VPW nch L=4e-08 W=3.75e-07 
M13 VSS 7 ECK VPW nch L=4e-08 W=3.75e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M15 4 E VDD VNW pch L=4e-08 W=2.3e-07 
M16 5 CK 4 VNW pch L=4e-08 W=1.8e-07 
M17 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M18 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M19 6 SEN VDD VNW pch L=4e-08 W=2.2e-07 
M20 VDD 5 6 VNW pch L=4e-08 W=2.2e-07 
M21 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M22 VDD CK 7 VNW pch L=4e-08 W=2e-07 
M23 7 CK VDD VNW pch L=4e-08 W=2e-07 
M24 VDD CK 7 VNW pch L=4e-08 W=2e-07 
M25 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M27 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M29 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X6B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=1.95e-07 
M2 5 1 4 VPW nch L=4e-08 W=1.95e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2.7e-07 
M6 6 5 14 VPW nch L=4e-08 W=2.7e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.9e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.9e-07 
M9 16 CK 7 VPW nch L=4e-08 W=2.9e-07 
M10 VSS 6 16 VPW nch L=4e-08 W=2.9e-07 
M11 ECK 7 VSS VPW nch L=4e-08 W=3.35e-07 
M12 VSS 7 ECK VPW nch L=4e-08 W=3.35e-07 
M13 ECK 7 VSS VPW nch L=4e-08 W=3.35e-07 
M14 VSS 7 ECK VPW nch L=4e-08 W=3.35e-07 
M15 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M16 4 E VDD VNW pch L=4e-08 W=2.5e-07 
M17 5 CK 4 VNW pch L=4e-08 W=1.95e-07 
M18 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M20 6 SEN VDD VNW pch L=4e-08 W=2.3e-07 
M21 VDD 5 6 VNW pch L=4e-08 W=2.3e-07 
M22 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M23 VDD CK 7 VNW pch L=4e-08 W=2.25e-07 
M24 7 CK VDD VNW pch L=4e-08 W=2.25e-07 
M25 VDD CK 7 VNW pch L=4e-08 W=2.25e-07 
M26 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M28 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M29 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M30 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT POSTICG_X7P5B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=2.1e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.1e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=2.9e-07 
M6 6 5 14 VPW nch L=4e-08 W=2.9e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.45e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.45e-07 
M9 16 CK 7 VPW nch L=4e-08 W=2.45e-07 
M10 VSS 6 16 VPW nch L=4e-08 W=2.45e-07 
M11 17 6 VSS VPW nch L=4e-08 W=2.45e-07 
M12 7 CK 17 VPW nch L=4e-08 W=2.45e-07 
M13 ECK 7 VSS VPW nch L=4e-08 W=2.85e-07 
M14 VSS 7 ECK VPW nch L=4e-08 W=2.85e-07 
M15 ECK 7 VSS VPW nch L=4e-08 W=2.85e-07 
M16 VSS 7 ECK VPW nch L=4e-08 W=2.85e-07 
M17 ECK 7 VSS VPW nch L=4e-08 W=2.85e-07 
M18 VSS 7 ECK VPW nch L=4e-08 W=2.85e-07 
M19 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M20 4 E VDD VNW pch L=4e-08 W=2.7e-07 
M21 5 CK 4 VNW pch L=4e-08 W=2.1e-07 
M22 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M24 6 SEN VDD VNW pch L=4e-08 W=2.5e-07 
M25 VDD 5 6 VNW pch L=4e-08 W=2.5e-07 
M26 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M27 7 CK VDD VNW pch L=4e-08 W=2.15e-07 
M28 VDD CK 7 VNW pch L=4e-08 W=2.15e-07 
M29 7 CK VDD VNW pch L=4e-08 W=2.15e-07 
M30 VDD CK 7 VNW pch L=4e-08 W=2.15e-07 
M31 ECK 7 VDD VNW pch L=4e-08 W=3.75e-07 
M32 VDD 7 ECK VNW pch L=4e-08 W=3.75e-07 
M33 ECK 7 VDD VNW pch L=4e-08 W=3.75e-07 
M34 VDD 7 ECK VNW pch L=4e-08 W=3.75e-07 
M35 ECK 7 VDD VNW pch L=4e-08 W=3.75e-07 
M36 VDD 7 ECK VNW pch L=4e-08 W=3.75e-07 
M37 ECK 7 VDD VNW pch L=4e-08 W=3.75e-07 
M38 VDD 7 ECK VNW pch L=4e-08 W=3.75e-07 
.ENDS


.SUBCKT POSTICG_X9B_A9TR ECK VDD VNW VPW VSS CK E SEN
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 E VSS VPW nch L=4e-08 W=2.3e-07 
M2 5 1 4 VPW nch L=4e-08 W=2.3e-07 
M3 13 CK 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 13 VPW nch L=4e-08 W=1.2e-07 
M5 14 SEN VSS VPW nch L=4e-08 W=3.5e-07 
M6 6 5 14 VPW nch L=4e-08 W=3.5e-07 
M7 15 CK 7 VPW nch L=4e-08 W=2.75e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=2.75e-07 
M9 16 6 VSS VPW nch L=4e-08 W=2.75e-07 
M10 7 CK 16 VPW nch L=4e-08 W=2.75e-07 
M11 17 CK 7 VPW nch L=4e-08 W=2.75e-07 
M12 VSS 6 17 VPW nch L=4e-08 W=2.75e-07 
M13 VSS 7 ECK VPW nch L=4e-08 W=2.9e-07 
M14 ECK 7 VSS VPW nch L=4e-08 W=2.9e-07 
M15 VSS 7 ECK VPW nch L=4e-08 W=2.9e-07 
M16 ECK 7 VSS VPW nch L=4e-08 W=2.9e-07 
M17 VSS 7 ECK VPW nch L=4e-08 W=2.9e-07 
M18 ECK 7 VSS VPW nch L=4e-08 W=2.9e-07 
M19 VSS 7 ECK VPW nch L=4e-08 W=2.9e-07 
M20 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M21 4 E VDD VNW pch L=4e-08 W=3e-07 
M22 5 CK 4 VNW pch L=4e-08 W=2.3e-07 
M23 12 1 5 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 6 12 VNW pch L=4e-08 W=1.2e-07 
M25 6 SEN VDD VNW pch L=4e-08 W=3e-07 
M26 VDD 5 6 VNW pch L=4e-08 W=3e-07 
M27 7 CK VDD VNW pch L=4e-08 W=2.4e-07 
M28 VDD CK 7 VNW pch L=4e-08 W=2.4e-07 
M29 7 CK VDD VNW pch L=4e-08 W=2.4e-07 
M30 VDD CK 7 VNW pch L=4e-08 W=2.4e-07 
M31 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M32 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M33 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M34 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M35 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M37 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M39 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X0P5B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 VSS E 4 VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=1.2e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M12 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.4e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT PREICG_X0P6B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 VSS E 4 VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=1.35e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M12 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.4e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT PREICG_X0P7B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 VSS E 4 VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=1.6e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M12 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.4e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT PREICG_X0P8B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 VSS E 4 VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=1.9e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M12 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.4e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT PREICG_X11B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=2.6e-07 
M2 4 E VSS VPW nch L=4e-08 W=2.6e-07 
M3 6 1 4 VPW nch L=4e-08 W=2.6e-07 
M4 14 CK 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 14 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2.4e-07 
M7 15 CK 8 VPW nch L=4e-08 W=3.4e-07 
M8 VSS 7 15 VPW nch L=4e-08 W=3.4e-07 
M9 16 7 VSS VPW nch L=4e-08 W=3.4e-07 
M10 8 CK 16 VPW nch L=4e-08 W=3.4e-07 
M11 17 CK 8 VPW nch L=4e-08 W=3.4e-07 
M12 VSS 7 17 VPW nch L=4e-08 W=3.4e-07 
M13 VSS 8 ECK VPW nch L=4e-08 W=3.55e-07 
M14 ECK 8 VSS VPW nch L=4e-08 W=3.55e-07 
M15 VSS 8 ECK VPW nch L=4e-08 W=3.55e-07 
M16 ECK 8 VSS VPW nch L=4e-08 W=3.55e-07 
M17 VSS 8 ECK VPW nch L=4e-08 W=3.55e-07 
M18 ECK 8 VSS VPW nch L=4e-08 W=3.55e-07 
M19 VSS 8 ECK VPW nch L=4e-08 W=3.55e-07 
M20 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M21 5 SE VDD VNW pch L=4e-08 W=3.2e-07 
M22 VDD SE 5 VNW pch L=4e-08 W=3.2e-07 
M23 4 E 5 VNW pch L=4e-08 W=3.35e-07 
M24 6 CK 4 VNW pch L=4e-08 W=2.6e-07 
M25 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M27 7 6 VDD VNW pch L=4e-08 W=3.1e-07 
M28 8 CK VDD VNW pch L=4e-08 W=2.25e-07 
M29 VDD CK 8 VNW pch L=4e-08 W=2.25e-07 
M30 8 CK VDD VNW pch L=4e-08 W=2.25e-07 
M31 VDD CK 8 VNW pch L=4e-08 W=2.25e-07 
M32 8 CK VDD VNW pch L=4e-08 W=2.25e-07 
M33 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M34 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M35 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M37 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M38 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M39 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M40 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M41 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M42 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M43 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M44 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X13B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=2.8e-07 
M2 4 E VSS VPW nch L=4e-08 W=2.8e-07 
M3 6 1 4 VPW nch L=4e-08 W=2.8e-07 
M4 15 CK 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2.6e-07 
M7 16 7 VSS VPW nch L=4e-08 W=3e-07 
M8 8 CK 16 VPW nch L=4e-08 W=3e-07 
M9 17 CK 8 VPW nch L=4e-08 W=3e-07 
M10 VSS 7 17 VPW nch L=4e-08 W=3e-07 
M11 18 7 VSS VPW nch L=4e-08 W=3e-07 
M12 8 CK 18 VPW nch L=4e-08 W=3e-07 
M13 19 CK 8 VPW nch L=4e-08 W=3e-07 
M14 VSS 7 19 VPW nch L=4e-08 W=3e-07 
M15 VSS 8 ECK VPW nch L=4e-08 W=3.25e-07 
M16 ECK 8 VSS VPW nch L=4e-08 W=3.25e-07 
M17 VSS 8 ECK VPW nch L=4e-08 W=3.25e-07 
M18 ECK 8 VSS VPW nch L=4e-08 W=3.25e-07 
M19 VSS 8 ECK VPW nch L=4e-08 W=3.25e-07 
M20 ECK 8 VSS VPW nch L=4e-08 W=3.25e-07 
M21 VSS 8 ECK VPW nch L=4e-08 W=3.25e-07 
M22 ECK 8 VSS VPW nch L=4e-08 W=3.25e-07 
M23 VSS 8 ECK VPW nch L=4e-08 W=3.25e-07 
M24 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M25 5 SE VDD VNW pch L=4e-08 W=3.4e-07 
M26 VDD SE 5 VNW pch L=4e-08 W=3.4e-07 
M27 4 E 5 VNW pch L=4e-08 W=3.6e-07 
M28 6 CK 4 VNW pch L=4e-08 W=2.8e-07 
M29 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M31 7 6 VDD VNW pch L=4e-08 W=3.4e-07 
M32 8 CK VDD VNW pch L=4e-08 W=2.3e-07 
M33 VDD CK 8 VNW pch L=4e-08 W=2.3e-07 
M34 8 CK VDD VNW pch L=4e-08 W=2.3e-07 
M35 VDD CK 8 VNW pch L=4e-08 W=2.3e-07 
M36 8 CK VDD VNW pch L=4e-08 W=2.3e-07 
M37 VDD CK 8 VNW pch L=4e-08 W=2.3e-07 
M38 8 7 VDD VNW pch L=4e-08 W=1.4e-07 
M39 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M40 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M41 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M42 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M43 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M44 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M45 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M46 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M47 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M48 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M49 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M50 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M51 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X16B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=3.1e-07 
M2 4 E VSS VPW nch L=4e-08 W=3.1e-07 
M3 6 1 4 VPW nch L=4e-08 W=3.1e-07 
M4 14 CK 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 14 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2.8e-07 
M7 15 7 VSS VPW nch L=4e-08 W=3.5e-07 
M8 8 CK 15 VPW nch L=4e-08 W=3.5e-07 
M9 16 CK 8 VPW nch L=4e-08 W=3.5e-07 
M10 VSS 7 16 VPW nch L=4e-08 W=3.5e-07 
M11 17 7 VSS VPW nch L=4e-08 W=3.5e-07 
M12 8 CK 17 VPW nch L=4e-08 W=3.5e-07 
M13 18 CK 8 VPW nch L=4e-08 W=3.5e-07 
M14 VSS 7 18 VPW nch L=4e-08 W=3.5e-07 
M15 ECK 8 VSS VPW nch L=4e-08 W=3.6e-07 
M16 VSS 8 ECK VPW nch L=4e-08 W=3.6e-07 
M17 ECK 8 VSS VPW nch L=4e-08 W=3.6e-07 
M18 VSS 8 ECK VPW nch L=4e-08 W=3.6e-07 
M19 ECK 8 VSS VPW nch L=4e-08 W=3.6e-07 
M20 VSS 8 ECK VPW nch L=4e-08 W=3.6e-07 
M21 ECK 8 VSS VPW nch L=4e-08 W=3.6e-07 
M22 VSS 8 ECK VPW nch L=4e-08 W=3.6e-07 
M23 ECK 8 VSS VPW nch L=4e-08 W=3.6e-07 
M24 VSS 8 ECK VPW nch L=4e-08 W=3.6e-07 
M25 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M26 5 SE VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD SE 5 VNW pch L=4e-08 W=3.8e-07 
M28 4 E 5 VNW pch L=4e-08 W=4e-07 
M29 6 CK 4 VNW pch L=4e-08 W=3.1e-07 
M30 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M32 7 6 VDD VNW pch L=4e-08 W=3.6e-07 
M33 8 7 VDD VNW pch L=4e-08 W=1.65e-07 
M34 VDD CK 8 VNW pch L=4e-08 W=2.35e-07 
M35 8 CK VDD VNW pch L=4e-08 W=2.35e-07 
M36 VDD CK 8 VNW pch L=4e-08 W=2.35e-07 
M37 8 CK VDD VNW pch L=4e-08 W=2.35e-07 
M38 VDD CK 8 VNW pch L=4e-08 W=2.35e-07 
M39 8 CK VDD VNW pch L=4e-08 W=2.35e-07 
M40 VDD CK 8 VNW pch L=4e-08 W=2.35e-07 
M41 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M42 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M43 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M44 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M45 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M46 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M47 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M48 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M49 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M50 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M51 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M52 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M53 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M54 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M55 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M56 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X1B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 VSS E 4 VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.2e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=2.25e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M12 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.4e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.4e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X1P2B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 VSS E 4 VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.45e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.45e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=2.7e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M12 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.7e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.4e-07 
M20 VDD 7 ECK VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT PREICG_X1P4B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 VSS E 4 VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 CK 7 VPW nch L=4e-08 W=1.6e-07 
M8 VSS 6 15 VPW nch L=4e-08 W=1.6e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=3.2e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M12 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M17 7 CK VDD VNW pch L=4e-08 W=1.9e-07 
M18 VDD 6 7 VNW pch L=4e-08 W=1.2e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=2.85e-07 
M20 VDD 7 ECK VNW pch L=4e-08 W=2.85e-07 
.ENDS


.SUBCKT PREICG_X1P7B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 VSS E 4 VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 6 VSS VPW nch L=4e-08 W=1.8e-07 
M8 7 CK 15 VPW nch L=4e-08 W=1.8e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=3.8e-07 
M10 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M11 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M12 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M13 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M14 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M17 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M18 VDD CK 7 VNW pch L=4e-08 W=2.1e-07 
M19 ECK 7 VDD VNW pch L=4e-08 W=3.35e-07 
M20 VDD 7 ECK VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT PREICG_X2B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 VSS E 4 VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.1e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.1e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=2.25e-07 
M10 VSS 7 ECK VPW nch L=4e-08 W=2.25e-07 
M11 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M12 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M13 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M14 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M15 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M16 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M17 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M19 VDD CK 7 VNW pch L=4e-08 W=2.4e-07 
M20 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X2P5B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.55e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.55e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=2.85e-07 
M10 VSS 7 ECK VPW nch L=4e-08 W=2.85e-07 
M11 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M12 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M13 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M14 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M15 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M16 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M17 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M19 VDD CK 7 VNW pch L=4e-08 W=2.95e-07 
M20 ECK 7 VDD VNW pch L=4e-08 W=3.35e-07 
M21 VDD 7 ECK VNW pch L=4e-08 W=3.35e-07 
M22 ECK 7 VDD VNW pch L=4e-08 W=3.35e-07 
.ENDS


.SUBCKT PREICG_X3B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.5e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.5e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.9e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.9e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=3.4e-07 
M10 VSS 7 ECK VPW nch L=4e-08 W=3.4e-07 
M11 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M12 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M13 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M14 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M15 13 1 5 VNW pch L=4e-08 W=1.5e-07 
M16 VDD 6 13 VNW pch L=4e-08 W=1.5e-07 
M17 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M19 VDD CK 7 VNW pch L=4e-08 W=3.4e-07 
M20 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M21 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M22 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X3P5B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.5e-07 
M2 4 E VSS VPW nch L=4e-08 W=1.5e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.5e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M7 15 6 VSS VPW nch L=4e-08 W=3.2e-07 
M8 7 CK 15 VPW nch L=4e-08 W=3.2e-07 
M9 ECK 7 VSS VPW nch L=4e-08 W=4e-07 
M10 VSS 7 ECK VPW nch L=4e-08 W=4e-07 
M11 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M12 12 SE VDD VNW pch L=4e-08 W=3.6e-07 
M13 4 E 12 VNW pch L=4e-08 W=1.95e-07 
M14 5 CK 4 VNW pch L=4e-08 W=1.5e-07 
M15 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M16 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M17 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M18 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M19 VDD CK 7 VNW pch L=4e-08 W=3.65e-07 
M20 ECK 7 VDD VNW pch L=4e-08 W=3.5e-07 
M21 VDD 7 ECK VNW pch L=4e-08 W=3.5e-07 
M22 ECK 7 VDD VNW pch L=4e-08 W=3.5e-07 
M23 VDD 7 ECK VNW pch L=4e-08 W=3.5e-07 
.ENDS


.SUBCKT PREICG_X4B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.7e-07 
M2 4 E VSS VPW nch L=4e-08 W=1.7e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.7e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.3e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.05e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.05e-07 
M9 16 CK 7 VPW nch L=4e-08 W=2.05e-07 
M10 VSS 6 16 VPW nch L=4e-08 W=2.05e-07 
M11 VSS 7 ECK VPW nch L=4e-08 W=3e-07 
M12 ECK 7 VSS VPW nch L=4e-08 W=3e-07 
M13 VSS 7 ECK VPW nch L=4e-08 W=3e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M15 12 SE VDD VNW pch L=4e-08 W=4e-07 
M16 4 E 12 VNW pch L=4e-08 W=2.7e-07 
M17 5 CK 4 VNW pch L=4e-08 W=1.7e-07 
M18 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M20 6 5 VDD VNW pch L=4e-08 W=1.7e-07 
M21 7 CK VDD VNW pch L=4e-08 W=2.4e-07 
M22 VDD CK 7 VNW pch L=4e-08 W=2.4e-07 
M23 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M24 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M25 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M26 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M27 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X5B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.8e-07 
M2 4 E VSS VPW nch L=4e-08 W=1.8e-07 
M3 5 1 4 VPW nch L=4e-08 W=1.8e-07 
M4 14 CK 5 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M6 6 5 VSS VPW nch L=4e-08 W=1.45e-07 
M7 15 6 VSS VPW nch L=4e-08 W=2.5e-07 
M8 7 CK 15 VPW nch L=4e-08 W=2.5e-07 
M9 16 CK 7 VPW nch L=4e-08 W=2.5e-07 
M10 VSS 6 16 VPW nch L=4e-08 W=2.5e-07 
M11 VSS 7 ECK VPW nch L=4e-08 W=3.75e-07 
M12 ECK 7 VSS VPW nch L=4e-08 W=3.75e-07 
M13 VSS 7 ECK VPW nch L=4e-08 W=3.75e-07 
M14 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M15 12 SE VDD VNW pch L=4e-08 W=4e-07 
M16 4 E 12 VNW pch L=4e-08 W=2.3e-07 
M17 5 CK 4 VNW pch L=4e-08 W=1.8e-07 
M18 13 1 5 VNW pch L=4e-08 W=1.2e-07 
M19 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M20 6 5 VDD VNW pch L=4e-08 W=1.9e-07 
M21 7 6 VDD VNW pch L=4e-08 W=1.2e-07 
M22 VDD CK 7 VNW pch L=4e-08 W=2e-07 
M23 7 CK VDD VNW pch L=4e-08 W=2e-07 
M24 VDD CK 7 VNW pch L=4e-08 W=2e-07 
M25 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M27 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 7 ECK VNW pch L=4e-08 W=4e-07 
M29 ECK 7 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X6B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=1.95e-07 
M2 4 E VSS VPW nch L=4e-08 W=1.95e-07 
M3 6 1 4 VPW nch L=4e-08 W=1.95e-07 
M4 14 CK 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 14 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.5e-07 
M7 15 7 VSS VPW nch L=4e-08 W=2.9e-07 
M8 8 CK 15 VPW nch L=4e-08 W=2.9e-07 
M9 16 CK 8 VPW nch L=4e-08 W=2.9e-07 
M10 VSS 7 16 VPW nch L=4e-08 W=2.9e-07 
M11 ECK 8 VSS VPW nch L=4e-08 W=3.35e-07 
M12 VSS 8 ECK VPW nch L=4e-08 W=3.35e-07 
M13 ECK 8 VSS VPW nch L=4e-08 W=3.35e-07 
M14 VSS 8 ECK VPW nch L=4e-08 W=3.35e-07 
M15 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M16 5 SE VDD VNW pch L=4e-08 W=2.3e-07 
M17 VDD SE 5 VNW pch L=4e-08 W=2.3e-07 
M18 4 E 5 VNW pch L=4e-08 W=2.8e-07 
M19 6 CK 4 VNW pch L=4e-08 W=1.95e-07 
M20 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M22 7 6 VDD VNW pch L=4e-08 W=2e-07 
M23 8 7 VDD VNW pch L=4e-08 W=1.2e-07 
M24 VDD CK 8 VNW pch L=4e-08 W=2.25e-07 
M25 8 CK VDD VNW pch L=4e-08 W=2.25e-07 
M26 VDD CK 8 VNW pch L=4e-08 W=2.25e-07 
M27 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M29 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M30 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M31 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M32 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT PREICG_X7P5B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=2.1e-07 
M2 4 E VSS VPW nch L=4e-08 W=2.1e-07 
M3 6 1 4 VPW nch L=4e-08 W=2.1e-07 
M4 15 CK 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 15 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=1.65e-07 
M7 16 7 VSS VPW nch L=4e-08 W=2.45e-07 
M8 8 CK 16 VPW nch L=4e-08 W=2.45e-07 
M9 17 CK 8 VPW nch L=4e-08 W=2.45e-07 
M10 VSS 7 17 VPW nch L=4e-08 W=2.45e-07 
M11 18 7 VSS VPW nch L=4e-08 W=2.45e-07 
M12 8 CK 18 VPW nch L=4e-08 W=2.45e-07 
M13 ECK 8 VSS VPW nch L=4e-08 W=2.85e-07 
M14 VSS 8 ECK VPW nch L=4e-08 W=2.85e-07 
M15 ECK 8 VSS VPW nch L=4e-08 W=2.85e-07 
M16 VSS 8 ECK VPW nch L=4e-08 W=2.85e-07 
M17 ECK 8 VSS VPW nch L=4e-08 W=2.85e-07 
M18 VSS 8 ECK VPW nch L=4e-08 W=2.85e-07 
M19 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M20 5 SE VDD VNW pch L=4e-08 W=2.55e-07 
M21 VDD SE 5 VNW pch L=4e-08 W=2.55e-07 
M22 4 E 5 VNW pch L=4e-08 W=2.7e-07 
M23 6 CK 4 VNW pch L=4e-08 W=2.1e-07 
M24 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M26 7 6 VDD VNW pch L=4e-08 W=2.15e-07 
M27 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M28 8 CK VDD VNW pch L=4e-08 W=2.15e-07 
M29 VDD CK 8 VNW pch L=4e-08 W=2.15e-07 
M30 8 CK VDD VNW pch L=4e-08 W=2.15e-07 
M31 VDD CK 8 VNW pch L=4e-08 W=2.15e-07 
M32 ECK 8 VDD VNW pch L=4e-08 W=3.75e-07 
M33 VDD 8 ECK VNW pch L=4e-08 W=3.75e-07 
M34 ECK 8 VDD VNW pch L=4e-08 W=3.75e-07 
M35 VDD 8 ECK VNW pch L=4e-08 W=3.75e-07 
M36 ECK 8 VDD VNW pch L=4e-08 W=3.75e-07 
M37 VDD 8 ECK VNW pch L=4e-08 W=3.75e-07 
M38 ECK 8 VDD VNW pch L=4e-08 W=3.75e-07 
M39 VDD 8 ECK VNW pch L=4e-08 W=3.75e-07 
.ENDS


.SUBCKT PREICG_X9B_A9TR ECK VDD VNW VPW VSS CK E SE
M0 VSS CK 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 SE VSS VPW nch L=4e-08 W=2.3e-07 
M2 4 E VSS VPW nch L=4e-08 W=2.3e-07 
M3 6 1 4 VPW nch L=4e-08 W=2.3e-07 
M4 14 CK 6 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 7 14 VPW nch L=4e-08 W=1.2e-07 
M6 7 6 VSS VPW nch L=4e-08 W=2e-07 
M7 15 CK 8 VPW nch L=4e-08 W=2.75e-07 
M8 VSS 7 15 VPW nch L=4e-08 W=2.75e-07 
M9 16 7 VSS VPW nch L=4e-08 W=2.75e-07 
M10 8 CK 16 VPW nch L=4e-08 W=2.75e-07 
M11 17 CK 8 VPW nch L=4e-08 W=2.75e-07 
M12 VSS 7 17 VPW nch L=4e-08 W=2.75e-07 
M13 VSS 8 ECK VPW nch L=4e-08 W=2.9e-07 
M14 ECK 8 VSS VPW nch L=4e-08 W=2.9e-07 
M15 VSS 8 ECK VPW nch L=4e-08 W=2.9e-07 
M16 ECK 8 VSS VPW nch L=4e-08 W=2.9e-07 
M17 VSS 8 ECK VPW nch L=4e-08 W=2.9e-07 
M18 ECK 8 VSS VPW nch L=4e-08 W=2.9e-07 
M19 VSS 8 ECK VPW nch L=4e-08 W=2.9e-07 
M20 VDD CK 1 VNW pch L=4e-08 W=1.55e-07 
M21 5 SE VDD VNW pch L=4e-08 W=2.7e-07 
M22 VDD SE 5 VNW pch L=4e-08 W=2.7e-07 
M23 4 E 5 VNW pch L=4e-08 W=3e-07 
M24 6 CK 4 VNW pch L=4e-08 W=2.3e-07 
M25 13 1 6 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 7 13 VNW pch L=4e-08 W=1.2e-07 
M27 7 6 VDD VNW pch L=4e-08 W=2.6e-07 
M28 8 CK VDD VNW pch L=4e-08 W=2.4e-07 
M29 VDD CK 8 VNW pch L=4e-08 W=2.4e-07 
M30 8 CK VDD VNW pch L=4e-08 W=2.4e-07 
M31 VDD CK 8 VNW pch L=4e-08 W=2.4e-07 
M32 8 7 VDD VNW pch L=4e-08 W=1.2e-07 
M33 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M34 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M35 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M36 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M37 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M38 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M39 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
M40 ECK 8 VDD VNW pch L=4e-08 W=4e-07 
M41 VDD 8 ECK VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT RF1R1WS_X1M_A9TR RBL VDD VNW VPW VSS RWL WBL WWL
M0 VSS WWL 1 VPW nch L=4e-08 W=1.8e-07 
M1 4 WBL VSS VPW nch L=4e-08 W=1.6e-07 
M2 5 WWL 4 VPW nch L=4e-08 W=1.6e-07 
M3 14 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 7 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 RBL RWL 7 VPW nch L=4e-08 W=3.1e-07 
M8 9 RWL VSS VPW nch L=4e-08 W=1.6e-07 
M9 VDD WWL 1 VNW pch L=4e-08 W=2.4e-07 
M10 4 WBL VDD VNW pch L=4e-08 W=2.3e-07 
M11 5 1 4 VNW pch L=4e-08 W=1.6e-07 
M12 13 WWL 5 VNW pch L=4e-08 W=1.2e-07 
M13 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M14 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M15 7 5 VDD VNW pch L=4e-08 W=4e-07 
M16 RBL 9 7 VNW pch L=4e-08 W=3.1e-07 
M17 9 RWL VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT RF1R1WS_X1P4M_A9TR RBL VDD VNW VPW VSS RWL WBL WWL
M0 VSS WWL 1 VPW nch L=4e-08 W=1.9e-07 
M1 4 WBL VSS VPW nch L=4e-08 W=2e-07 
M2 5 WWL 4 VPW nch L=4e-08 W=2e-07 
M3 14 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 7 5 VSS VPW nch L=4e-08 W=2.2e-07 
M7 VSS 5 7 VPW nch L=4e-08 W=2.2e-07 
M8 RBL RWL 7 VPW nch L=4e-08 W=2.2e-07 
M9 7 RWL RBL VPW nch L=4e-08 W=2.2e-07 
M10 9 RWL VSS VPW nch L=4e-08 W=2.1e-07 
M11 VDD WWL 1 VNW pch L=4e-08 W=2.4e-07 
M12 4 WBL VDD VNW pch L=4e-08 W=2.9e-07 
M13 5 1 4 VNW pch L=4e-08 W=2e-07 
M14 13 WWL 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M17 7 5 VDD VNW pch L=4e-08 W=2.85e-07 
M18 VDD 5 7 VNW pch L=4e-08 W=2.85e-07 
M19 RBL 9 7 VNW pch L=4e-08 W=2.2e-07 
M20 7 9 RBL VNW pch L=4e-08 W=2.2e-07 
M21 9 RWL VDD VNW pch L=4e-08 W=2.7e-07 
.ENDS


.SUBCKT RF1R1WS_X2M_A9TR RBL VDD VNW VPW VSS RWL WBL WWL
M0 VSS WWL 1 VPW nch L=4e-08 W=2e-07 
M1 4 WBL VSS VPW nch L=4e-08 W=2.5e-07 
M2 5 WWL 4 VPW nch L=4e-08 W=2.5e-07 
M3 14 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 14 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 7 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 5 7 VPW nch L=4e-08 W=3.1e-07 
M8 RBL RWL 7 VPW nch L=4e-08 W=3.1e-07 
M9 7 RWL RBL VPW nch L=4e-08 W=3.1e-07 
M10 9 RWL VSS VPW nch L=4e-08 W=2.65e-07 
M11 VDD WWL 1 VNW pch L=4e-08 W=2.6e-07 
M12 4 WBL VDD VNW pch L=4e-08 W=3.3e-07 
M13 5 1 4 VNW pch L=4e-08 W=2.5e-07 
M14 13 WWL 5 VNW pch L=4e-08 W=1.2e-07 
M15 VDD 6 13 VNW pch L=4e-08 W=1.2e-07 
M16 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M17 7 5 VDD VNW pch L=4e-08 W=4e-07 
M18 VDD 5 7 VNW pch L=4e-08 W=4e-07 
M19 RBL 9 7 VNW pch L=4e-08 W=3.1e-07 
M20 7 9 RBL VNW pch L=4e-08 W=3.1e-07 
M21 9 RWL VDD VNW pch L=4e-08 W=3.4e-07 
.ENDS


.SUBCKT RF1R2WS_X1M_A9TR RBL VDD VNW VPW VSS RWL WBL1 WBL2 WWL1 WWL2
M0 VSS WWL1 1 VPW nch L=4e-08 W=1.9e-07 
M1 4 WBL1 VSS VPW nch L=4e-08 W=2e-07 
M2 5 WWL1 4 VPW nch L=4e-08 W=2e-07 
M3 19 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 20 6 19 VPW nch L=4e-08 W=1.6e-07 
M5 VSS 8 20 VPW nch L=4e-08 W=1.6e-07 
M6 6 WWL2 VSS VPW nch L=4e-08 W=1.9e-07 
M7 7 WWL2 5 VPW nch L=4e-08 W=2e-07 
M8 VSS WBL2 7 VPW nch L=4e-08 W=2e-07 
M9 VSS 5 8 VPW nch L=4e-08 W=1.2e-07 
M10 9 5 VSS VPW nch L=4e-08 W=3.1e-07 
M11 RBL RWL 9 VPW nch L=4e-08 W=3.1e-07 
M12 11 RWL VSS VPW nch L=4e-08 W=1.6e-07 
M13 VDD WWL1 1 VNW pch L=4e-08 W=2.5e-07 
M14 4 WBL1 VDD VNW pch L=4e-08 W=2.6e-07 
M15 5 1 4 VNW pch L=4e-08 W=2e-07 
M16 17 WWL1 5 VNW pch L=4e-08 W=1.6e-07 
M17 18 WWL2 17 VNW pch L=4e-08 W=1.6e-07 
M18 VDD 8 18 VNW pch L=4e-08 W=1.6e-07 
M19 6 WWL2 VDD VNW pch L=4e-08 W=2.5e-07 
M20 7 6 5 VNW pch L=4e-08 W=2e-07 
M21 VDD WBL2 7 VNW pch L=4e-08 W=2.6e-07 
M22 VDD 5 8 VNW pch L=4e-08 W=1.2e-07 
M23 9 5 VDD VNW pch L=4e-08 W=4e-07 
M24 RBL 11 9 VNW pch L=4e-08 W=3.1e-07 
M25 11 RWL VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT RF1R2WS_X1P4M_A9TR RBL VDD VNW VPW VSS RWL WBL1 WBL2 WWL1 WWL2
M0 VSS WWL1 1 VPW nch L=4e-08 W=1.9e-07 
M1 4 WBL1 VSS VPW nch L=4e-08 W=2.2e-07 
M2 5 WWL1 4 VPW nch L=4e-08 W=2.2e-07 
M3 19 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 20 6 19 VPW nch L=4e-08 W=1.6e-07 
M5 VSS 8 20 VPW nch L=4e-08 W=1.6e-07 
M6 6 WWL2 VSS VPW nch L=4e-08 W=1.9e-07 
M7 7 WWL2 5 VPW nch L=4e-08 W=2.2e-07 
M8 VSS WBL2 7 VPW nch L=4e-08 W=2.2e-07 
M9 VSS 5 8 VPW nch L=4e-08 W=1.2e-07 
M10 9 5 VSS VPW nch L=4e-08 W=2.2e-07 
M11 VSS 5 9 VPW nch L=4e-08 W=2.2e-07 
M12 RBL RWL 9 VPW nch L=4e-08 W=2.2e-07 
M13 9 RWL RBL VPW nch L=4e-08 W=2.2e-07 
M14 11 RWL VSS VPW nch L=4e-08 W=2.1e-07 
M15 VDD WWL1 1 VNW pch L=4e-08 W=2.5e-07 
M16 4 WBL1 VDD VNW pch L=4e-08 W=2.8e-07 
M17 5 1 4 VNW pch L=4e-08 W=2.2e-07 
M18 17 WWL1 5 VNW pch L=4e-08 W=1.6e-07 
M19 18 WWL2 17 VNW pch L=4e-08 W=1.6e-07 
M20 VDD 8 18 VNW pch L=4e-08 W=1.6e-07 
M21 6 WWL2 VDD VNW pch L=4e-08 W=2.5e-07 
M22 7 6 5 VNW pch L=4e-08 W=2.2e-07 
M23 VDD WBL2 7 VNW pch L=4e-08 W=2.8e-07 
M24 VDD 5 8 VNW pch L=4e-08 W=1.2e-07 
M25 9 5 VDD VNW pch L=4e-08 W=2.85e-07 
M26 VDD 5 9 VNW pch L=4e-08 W=2.85e-07 
M27 RBL 11 9 VNW pch L=4e-08 W=2.2e-07 
M28 9 11 RBL VNW pch L=4e-08 W=2.2e-07 
M29 11 RWL VDD VNW pch L=4e-08 W=2.7e-07 
.ENDS


.SUBCKT RF1R2WS_X2M_A9TR RBL VDD VNW VPW VSS RWL WBL1 WBL2 WWL1 WWL2
M0 VSS WWL1 1 VPW nch L=4e-08 W=2.1e-07 
M1 4 WBL1 VSS VPW nch L=4e-08 W=2.8e-07 
M2 5 WWL1 4 VPW nch L=4e-08 W=2.8e-07 
M3 19 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 20 6 19 VPW nch L=4e-08 W=1.6e-07 
M5 VSS 8 20 VPW nch L=4e-08 W=1.6e-07 
M6 6 WWL2 VSS VPW nch L=4e-08 W=2.1e-07 
M7 7 WWL2 5 VPW nch L=4e-08 W=2.8e-07 
M8 VSS WBL2 7 VPW nch L=4e-08 W=2.8e-07 
M9 VSS 5 8 VPW nch L=4e-08 W=1.2e-07 
M10 9 5 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 5 9 VPW nch L=4e-08 W=3.1e-07 
M12 RBL RWL 9 VPW nch L=4e-08 W=3.1e-07 
M13 9 RWL RBL VPW nch L=4e-08 W=3.1e-07 
M14 11 RWL VSS VPW nch L=4e-08 W=2.65e-07 
M15 VDD WWL1 1 VNW pch L=4e-08 W=2.7e-07 
M16 4 WBL1 VDD VNW pch L=4e-08 W=3.6e-07 
M17 5 1 4 VNW pch L=4e-08 W=2.8e-07 
M18 17 WWL1 5 VNW pch L=4e-08 W=1.6e-07 
M19 18 WWL2 17 VNW pch L=4e-08 W=1.6e-07 
M20 VDD 8 18 VNW pch L=4e-08 W=1.6e-07 
M21 6 WWL2 VDD VNW pch L=4e-08 W=2.7e-07 
M22 7 6 5 VNW pch L=4e-08 W=2.8e-07 
M23 VDD WBL2 7 VNW pch L=4e-08 W=3.6e-07 
M24 VDD 5 8 VNW pch L=4e-08 W=1.2e-07 
M25 9 5 VDD VNW pch L=4e-08 W=4e-07 
M26 VDD 5 9 VNW pch L=4e-08 W=4e-07 
M27 RBL 11 9 VNW pch L=4e-08 W=3.1e-07 
M28 9 11 RBL VNW pch L=4e-08 W=3.1e-07 
M29 11 RWL VDD VNW pch L=4e-08 W=3.4e-07 
.ENDS


.SUBCKT RF2R1WS_X1M_A9TR RBL1 RBL2 VDD VNW VPW VSS RWL1 RWL2 WBL WWL
M0 VSS WWL 1 VPW nch L=4e-08 W=2.2e-07 
M1 4 WBL VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 WWL 4 VPW nch L=4e-08 W=2.9e-07 
M3 18 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 18 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 7 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 RBL1 RWL1 7 VPW nch L=4e-08 W=3.1e-07 
M8 9 RWL1 VSS VPW nch L=4e-08 W=1.6e-07 
M9 10 5 VSS VPW nch L=4e-08 W=3.1e-07 
M10 RBL2 RWL2 10 VPW nch L=4e-08 W=3.1e-07 
M11 12 RWL2 VSS VPW nch L=4e-08 W=1.6e-07 
M12 VDD WWL 1 VNW pch L=4e-08 W=2.8e-07 
M13 4 WBL VDD VNW pch L=4e-08 W=3.8e-07 
M14 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M15 17 WWL 5 VNW pch L=4e-08 W=1.2e-07 
M16 VDD 6 17 VNW pch L=4e-08 W=1.2e-07 
M17 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M18 7 5 VDD VNW pch L=4e-08 W=4e-07 
M19 RBL1 9 7 VNW pch L=4e-08 W=3.1e-07 
M20 9 RWL1 VDD VNW pch L=4e-08 W=2.1e-07 
M21 10 5 VDD VNW pch L=4e-08 W=4e-07 
M22 RBL2 12 10 VNW pch L=4e-08 W=3.1e-07 
M23 12 RWL2 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT RF2R1WS_X1P4M_A9TR RBL1 RBL2 VDD VNW VPW VSS RWL1 RWL2 WBL WWL
M0 VSS WWL 1 VPW nch L=4e-08 W=2.2e-07 
M1 4 WBL VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 WWL 4 VPW nch L=4e-08 W=2.9e-07 
M3 18 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 18 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 7 5 VSS VPW nch L=4e-08 W=2.2e-07 
M7 VSS 5 7 VPW nch L=4e-08 W=2.2e-07 
M8 RBL1 RWL1 7 VPW nch L=4e-08 W=2.2e-07 
M9 7 RWL1 RBL1 VPW nch L=4e-08 W=2.2e-07 
M10 9 RWL1 VSS VPW nch L=4e-08 W=2.1e-07 
M11 10 5 VSS VPW nch L=4e-08 W=2.2e-07 
M12 VSS 5 10 VPW nch L=4e-08 W=2.2e-07 
M13 RBL2 RWL2 10 VPW nch L=4e-08 W=2.2e-07 
M14 10 RWL2 RBL2 VPW nch L=4e-08 W=2.2e-07 
M15 12 RWL2 VSS VPW nch L=4e-08 W=2.1e-07 
M16 VDD WWL 1 VNW pch L=4e-08 W=2.8e-07 
M17 4 WBL VDD VNW pch L=4e-08 W=3.8e-07 
M18 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M19 17 WWL 5 VNW pch L=4e-08 W=1.2e-07 
M20 VDD 6 17 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M22 7 5 VDD VNW pch L=4e-08 W=2.85e-07 
M23 VDD 5 7 VNW pch L=4e-08 W=2.85e-07 
M24 RBL1 9 7 VNW pch L=4e-08 W=2.2e-07 
M25 7 9 RBL1 VNW pch L=4e-08 W=2.2e-07 
M26 9 RWL1 VDD VNW pch L=4e-08 W=2.7e-07 
M27 10 5 VDD VNW pch L=4e-08 W=2.85e-07 
M28 VDD 5 10 VNW pch L=4e-08 W=2.85e-07 
M29 RBL2 12 10 VNW pch L=4e-08 W=2.2e-07 
M30 10 12 RBL2 VNW pch L=4e-08 W=2.2e-07 
M31 12 RWL2 VDD VNW pch L=4e-08 W=2.7e-07 
.ENDS


.SUBCKT RF2R1WS_X2M_A9TR RBL1 RBL2 VDD VNW VPW VSS RWL1 RWL2 WBL WWL
M0 VSS WWL 1 VPW nch L=4e-08 W=2.2e-07 
M1 4 WBL VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 WWL 4 VPW nch L=4e-08 W=2.9e-07 
M3 18 1 5 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 6 18 VPW nch L=4e-08 W=1.2e-07 
M5 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M6 7 5 VSS VPW nch L=4e-08 W=3.1e-07 
M7 VSS 5 7 VPW nch L=4e-08 W=3.1e-07 
M8 RBL1 RWL1 7 VPW nch L=4e-08 W=3.1e-07 
M9 7 RWL1 RBL1 VPW nch L=4e-08 W=3.1e-07 
M10 9 RWL1 VSS VPW nch L=4e-08 W=2.65e-07 
M11 10 5 VSS VPW nch L=4e-08 W=3.1e-07 
M12 VSS 5 10 VPW nch L=4e-08 W=3.1e-07 
M13 RBL2 RWL2 10 VPW nch L=4e-08 W=3.1e-07 
M14 10 RWL2 RBL2 VPW nch L=4e-08 W=3.1e-07 
M15 12 RWL2 VSS VPW nch L=4e-08 W=2.65e-07 
M16 VDD WWL 1 VNW pch L=4e-08 W=2.8e-07 
M17 4 WBL VDD VNW pch L=4e-08 W=3.8e-07 
M18 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M19 17 WWL 5 VNW pch L=4e-08 W=1.2e-07 
M20 VDD 6 17 VNW pch L=4e-08 W=1.2e-07 
M21 VDD 5 6 VNW pch L=4e-08 W=1.2e-07 
M22 7 5 VDD VNW pch L=4e-08 W=4e-07 
M23 VDD 5 7 VNW pch L=4e-08 W=4e-07 
M24 RBL1 9 7 VNW pch L=4e-08 W=3.1e-07 
M25 7 9 RBL1 VNW pch L=4e-08 W=3.1e-07 
M26 9 RWL1 VDD VNW pch L=4e-08 W=3.4e-07 
M27 10 5 VDD VNW pch L=4e-08 W=4e-07 
M28 VDD 5 10 VNW pch L=4e-08 W=4e-07 
M29 RBL2 12 10 VNW pch L=4e-08 W=3.1e-07 
M30 10 12 RBL2 VNW pch L=4e-08 W=3.1e-07 
M31 12 RWL2 VDD VNW pch L=4e-08 W=3.4e-07 
.ENDS


.SUBCKT RF2R2WS_X1M_A9TR RBL1 RBL2 VDD VNW VPW VSS RWL1 RWL2 WBL1 WBL2 WWL1 WWL2
M0 VSS WWL1 1 VPW nch L=4e-08 W=2.2e-07 
M1 4 WBL1 VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 WWL1 4 VPW nch L=4e-08 W=2.9e-07 
M3 23 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 24 6 23 VPW nch L=4e-08 W=1.6e-07 
M5 VSS 8 24 VPW nch L=4e-08 W=1.6e-07 
M6 6 WWL2 VSS VPW nch L=4e-08 W=2.2e-07 
M7 7 WWL2 5 VPW nch L=4e-08 W=2.9e-07 
M8 VSS WBL2 7 VPW nch L=4e-08 W=2.9e-07 
M9 VSS 5 8 VPW nch L=4e-08 W=1.2e-07 
M10 9 5 VSS VPW nch L=4e-08 W=3.1e-07 
M11 RBL1 RWL1 9 VPW nch L=4e-08 W=3.1e-07 
M12 11 RWL1 VSS VPW nch L=4e-08 W=1.6e-07 
M13 12 5 VSS VPW nch L=4e-08 W=3.1e-07 
M14 RBL2 RWL2 12 VPW nch L=4e-08 W=3.1e-07 
M15 14 RWL2 VSS VPW nch L=4e-08 W=1.6e-07 
M16 VDD WWL1 1 VNW pch L=4e-08 W=2.8e-07 
M17 4 WBL1 VDD VNW pch L=4e-08 W=3.8e-07 
M18 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M19 21 WWL1 5 VNW pch L=4e-08 W=1.6e-07 
M20 22 WWL2 21 VNW pch L=4e-08 W=1.6e-07 
M21 VDD 8 22 VNW pch L=4e-08 W=1.6e-07 
M22 6 WWL2 VDD VNW pch L=4e-08 W=2.8e-07 
M23 7 6 5 VNW pch L=4e-08 W=2.9e-07 
M24 VDD WBL2 7 VNW pch L=4e-08 W=3.8e-07 
M25 VDD 5 8 VNW pch L=4e-08 W=1.2e-07 
M26 9 5 VDD VNW pch L=4e-08 W=4e-07 
M27 RBL1 11 9 VNW pch L=4e-08 W=3.1e-07 
M28 11 RWL1 VDD VNW pch L=4e-08 W=2.1e-07 
M29 12 5 VDD VNW pch L=4e-08 W=4e-07 
M30 RBL2 14 12 VNW pch L=4e-08 W=3.1e-07 
M31 14 RWL2 VDD VNW pch L=4e-08 W=2.1e-07 
.ENDS


.SUBCKT RF2R2WS_X1P4M_A9TR RBL1 RBL2 VDD VNW VPW VSS RWL1 RWL2 WBL1 WBL2 WWL1 WWL2
M0 VSS WWL1 1 VPW nch L=4e-08 W=2.2e-07 
M1 4 WBL1 VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 WWL1 4 VPW nch L=4e-08 W=2.9e-07 
M3 23 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 24 6 23 VPW nch L=4e-08 W=1.6e-07 
M5 VSS 8 24 VPW nch L=4e-08 W=1.6e-07 
M6 6 WWL2 VSS VPW nch L=4e-08 W=2.2e-07 
M7 7 WWL2 5 VPW nch L=4e-08 W=2.9e-07 
M8 VSS WBL2 7 VPW nch L=4e-08 W=2.9e-07 
M9 VSS 5 8 VPW nch L=4e-08 W=1.2e-07 
M10 9 5 VSS VPW nch L=4e-08 W=2.2e-07 
M11 VSS 5 9 VPW nch L=4e-08 W=2.2e-07 
M12 RBL1 RWL1 9 VPW nch L=4e-08 W=2.2e-07 
M13 9 RWL1 RBL1 VPW nch L=4e-08 W=2.2e-07 
M14 11 RWL1 VSS VPW nch L=4e-08 W=2.1e-07 
M15 12 5 VSS VPW nch L=4e-08 W=2.2e-07 
M16 VSS 5 12 VPW nch L=4e-08 W=2.2e-07 
M17 RBL2 RWL2 12 VPW nch L=4e-08 W=2.2e-07 
M18 12 RWL2 RBL2 VPW nch L=4e-08 W=2.2e-07 
M19 14 RWL2 VSS VPW nch L=4e-08 W=2.1e-07 
M20 VDD WWL1 1 VNW pch L=4e-08 W=2.8e-07 
M21 4 WBL1 VDD VNW pch L=4e-08 W=3.8e-07 
M22 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M23 21 WWL1 5 VNW pch L=4e-08 W=1.6e-07 
M24 22 WWL2 21 VNW pch L=4e-08 W=1.6e-07 
M25 VDD 8 22 VNW pch L=4e-08 W=1.6e-07 
M26 6 WWL2 VDD VNW pch L=4e-08 W=2.8e-07 
M27 7 6 5 VNW pch L=4e-08 W=2.9e-07 
M28 VDD WBL2 7 VNW pch L=4e-08 W=3.8e-07 
M29 VDD 5 8 VNW pch L=4e-08 W=1.2e-07 
M30 9 5 VDD VNW pch L=4e-08 W=2.85e-07 
M31 VDD 5 9 VNW pch L=4e-08 W=2.85e-07 
M32 RBL1 11 9 VNW pch L=4e-08 W=2.2e-07 
M33 9 11 RBL1 VNW pch L=4e-08 W=2.2e-07 
M34 11 RWL1 VDD VNW pch L=4e-08 W=2.7e-07 
M35 12 5 VDD VNW pch L=4e-08 W=2.85e-07 
M36 VDD 5 12 VNW pch L=4e-08 W=2.85e-07 
M37 RBL2 14 12 VNW pch L=4e-08 W=2.2e-07 
M38 12 14 RBL2 VNW pch L=4e-08 W=2.2e-07 
M39 14 RWL2 VDD VNW pch L=4e-08 W=2.7e-07 
.ENDS


.SUBCKT RF2R2WS_X2M_A9TR RBL1 RBL2 VDD VNW VPW VSS RWL1 RWL2 WBL1 WBL2 WWL1 WWL2
M0 VSS WWL1 1 VPW nch L=4e-08 W=2.2e-07 
M1 4 WBL1 VSS VPW nch L=4e-08 W=2.9e-07 
M2 5 WWL1 4 VPW nch L=4e-08 W=2.9e-07 
M3 23 1 5 VPW nch L=4e-08 W=1.6e-07 
M4 24 6 23 VPW nch L=4e-08 W=1.6e-07 
M5 VSS 8 24 VPW nch L=4e-08 W=1.6e-07 
M6 6 WWL2 VSS VPW nch L=4e-08 W=2.2e-07 
M7 7 WWL2 5 VPW nch L=4e-08 W=2.9e-07 
M8 VSS WBL2 7 VPW nch L=4e-08 W=2.9e-07 
M9 VSS 5 8 VPW nch L=4e-08 W=1.2e-07 
M10 9 5 VSS VPW nch L=4e-08 W=3.1e-07 
M11 VSS 5 9 VPW nch L=4e-08 W=3.1e-07 
M12 RBL1 RWL1 9 VPW nch L=4e-08 W=3.1e-07 
M13 9 RWL1 RBL1 VPW nch L=4e-08 W=3.1e-07 
M14 11 RWL1 VSS VPW nch L=4e-08 W=2.65e-07 
M15 12 5 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 5 12 VPW nch L=4e-08 W=3.1e-07 
M17 RBL2 RWL2 12 VPW nch L=4e-08 W=3.1e-07 
M18 12 RWL2 RBL2 VPW nch L=4e-08 W=3.1e-07 
M19 14 RWL2 VSS VPW nch L=4e-08 W=2.65e-07 
M20 VDD WWL1 1 VNW pch L=4e-08 W=2.8e-07 
M21 4 WBL1 VDD VNW pch L=4e-08 W=3.8e-07 
M22 5 1 4 VNW pch L=4e-08 W=2.9e-07 
M23 21 WWL1 5 VNW pch L=4e-08 W=1.6e-07 
M24 22 WWL2 21 VNW pch L=4e-08 W=1.6e-07 
M25 VDD 8 22 VNW pch L=4e-08 W=1.6e-07 
M26 6 WWL2 VDD VNW pch L=4e-08 W=2.8e-07 
M27 7 6 5 VNW pch L=4e-08 W=2.9e-07 
M28 VDD WBL2 7 VNW pch L=4e-08 W=3.8e-07 
M29 VDD 5 8 VNW pch L=4e-08 W=1.2e-07 
M30 9 5 VDD VNW pch L=4e-08 W=4e-07 
M31 VDD 5 9 VNW pch L=4e-08 W=4e-07 
M32 RBL1 11 9 VNW pch L=4e-08 W=3.1e-07 
M33 9 11 RBL1 VNW pch L=4e-08 W=3.1e-07 
M34 11 RWL1 VDD VNW pch L=4e-08 W=3.4e-07 
M35 12 5 VDD VNW pch L=4e-08 W=4e-07 
M36 VDD 5 12 VNW pch L=4e-08 W=4e-07 
M37 RBL2 14 12 VNW pch L=4e-08 W=3.1e-07 
M38 12 14 RBL2 VNW pch L=4e-08 W=3.1e-07 
M39 14 RWL2 VDD VNW pch L=4e-08 W=3.4e-07 
.ENDS


.SUBCKT SDFFNQ_X1M_A9TR Q VDD VNW VPW VSS CKN D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=1.2e-07 
M4 4 D 21 VPW nch L=4e-08 W=1.2e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.2e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M9 7 10 6 VPW nch L=4e-08 W=1.2e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 7 8 VPW nch L=4e-08 W=2e-07 
M13 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M14 VSS CKN 10 VPW nch L=4e-08 W=1.2e-07 
M15 11 10 VSS VPW nch L=4e-08 W=1.2e-07 
M16 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M17 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M18 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M19 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M20 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M21 5 10 4 VNW pch L=4e-08 W=2e-07 
M22 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M24 6 5 VDD VNW pch L=4e-08 W=2e-07 
M25 7 11 6 VNW pch L=4e-08 W=2e-07 
M26 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 7 8 VNW pch L=4e-08 W=2e-07 
M29 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD CKN 10 VNW pch L=4e-08 W=2.5e-07 
M31 11 10 VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFNQ_X2M_A9TR Q VDD VNW VPW VSS CKN D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=1.2e-07 
M4 4 D 21 VPW nch L=4e-08 W=1.2e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.55e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=1.55e-07 
M9 7 10 6 VPW nch L=4e-08 W=1.55e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 8 7 VSS VPW nch L=4e-08 W=3.1e-07 
M13 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M14 VSS 8 Q VPW nch L=4e-08 W=2e-07 
M15 VSS CKN 10 VPW nch L=4e-08 W=1.3e-07 
M16 11 10 VSS VPW nch L=4e-08 W=1.3e-07 
M17 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M18 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M19 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M20 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M21 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M22 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M23 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M25 6 5 VDD VNW pch L=4e-08 W=3.1e-07 
M26 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M27 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M29 8 7 VDD VNW pch L=4e-08 W=3.1e-07 
M30 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M32 VDD CKN 10 VNW pch L=4e-08 W=2.7e-07 
M33 11 10 VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFNQ_X3M_A9TR Q VDD VNW VPW VSS CKN D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=1.2e-07 
M4 4 D 21 VPW nch L=4e-08 W=1.2e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.55e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=1.8e-07 
M9 7 10 6 VPW nch L=4e-08 W=1.55e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 8 7 VSS VPW nch L=4e-08 W=1.9e-07 
M13 VSS 7 8 VPW nch L=4e-08 W=1.9e-07 
M14 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M15 VSS 8 Q VPW nch L=4e-08 W=2e-07 
M16 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M17 VSS CKN 10 VPW nch L=4e-08 W=1.3e-07 
M18 11 10 VSS VPW nch L=4e-08 W=1.3e-07 
M19 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M20 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M21 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M22 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M23 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M24 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M25 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M27 6 5 VDD VNW pch L=4e-08 W=3.8e-07 
M28 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M29 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M31 8 7 VDD VNW pch L=4e-08 W=1.9e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=1.9e-07 
M33 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M35 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD CKN 10 VNW pch L=4e-08 W=2.7e-07 
M37 11 10 VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFNRPQ_X1M_A9TR Q VDD VNW VPW VSS CKN D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=1.2e-07 
M4 4 D 24 VPW nch L=4e-08 W=1.2e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.2e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=1.2e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.2e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=2e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M16 VSS CKN 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 10 VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=3.6e-07 
M22 4 D 18 VNW pch L=4e-08 W=3.6e-07 
M23 5 10 4 VNW pch L=4e-08 W=2e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M26 20 R VDD VNW pch L=4e-08 W=3.6e-07 
M27 6 5 20 VNW pch L=4e-08 W=3.6e-07 
M28 7 11 6 VNW pch L=4e-08 W=2e-07 
M29 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M30 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M31 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=2e-07 
M33 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD CKN 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 10 VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFNRPQ_X2M_A9TR Q VDD VNW VPW VSS CKN D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=1.3e-07 
M4 4 D 24 VPW nch L=4e-08 W=1.3e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.55e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=1.2e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.55e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=3.1e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M16 VSS 8 Q VPW nch L=4e-08 W=2e-07 
M17 VSS CKN 10 VPW nch L=4e-08 W=1.3e-07 
M18 11 10 VSS VPW nch L=4e-08 W=1.3e-07 
M19 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M20 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M21 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M22 18 SE VDD VNW pch L=4e-08 W=3.8e-07 
M23 4 D 18 VNW pch L=4e-08 W=3.8e-07 
M24 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M25 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M27 20 R VDD VNW pch L=4e-08 W=3.8e-07 
M28 6 5 20 VNW pch L=4e-08 W=3.8e-07 
M29 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M30 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M31 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M32 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M33 VDD 7 8 VNW pch L=4e-08 W=3.1e-07 
M34 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M36 VDD CKN 10 VNW pch L=4e-08 W=2.7e-07 
M37 11 10 VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFNRPQ_X3M_A9TR Q VDD VNW VPW VSS CKN D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=1.35e-07 
M4 4 D 24 VPW nch L=4e-08 W=1.35e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.55e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=1.2e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.55e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=3.8e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M16 VSS 8 Q VPW nch L=4e-08 W=2e-07 
M17 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M18 VSS CKN 10 VPW nch L=4e-08 W=1.3e-07 
M19 11 10 VSS VPW nch L=4e-08 W=1.3e-07 
M20 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M21 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M22 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M23 18 SE VDD VNW pch L=4e-08 W=3.8e-07 
M24 4 D 18 VNW pch L=4e-08 W=3.8e-07 
M25 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M26 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M28 20 R VDD VNW pch L=4e-08 W=3.8e-07 
M29 6 5 20 VNW pch L=4e-08 W=3.8e-07 
M30 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M31 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M32 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M33 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M34 VDD 7 8 VNW pch L=4e-08 W=3.8e-07 
M35 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M37 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M38 VDD CKN 10 VNW pch L=4e-08 W=2.7e-07 
M39 11 10 VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFNSQ_X1M_A9TR Q VDD VNW VPW VSS CKN D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=1.2e-07 
M4 4 D 22 VPW nch L=4e-08 W=1.2e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.2e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.5e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.5e-07 
M8 24 SN VSS VPW nch L=4e-08 W=1.8e-07 
M9 6 5 24 VPW nch L=4e-08 W=1.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.2e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=2e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M16 VSS CKN 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 10 VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=3.6e-07 
M22 4 D 18 VNW pch L=4e-08 W=3.6e-07 
M23 5 10 4 VNW pch L=4e-08 W=2e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.5e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.5e-07 
M26 6 SN VDD VNW pch L=4e-08 W=2e-07 
M27 VDD 5 6 VNW pch L=4e-08 W=2e-07 
M28 7 11 6 VNW pch L=4e-08 W=2e-07 
M29 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M31 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=2e-07 
M33 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD CKN 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 10 VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFNSQ_X2M_A9TR Q VDD VNW VPW VSS CKN D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=1.3e-07 
M4 4 D 22 VPW nch L=4e-08 W=1.3e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.55e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.5e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.5e-07 
M8 24 SN VSS VPW nch L=4e-08 W=2.8e-07 
M9 6 5 24 VPW nch L=4e-08 W=2.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.55e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=3.1e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M16 VSS 8 Q VPW nch L=4e-08 W=2e-07 
M17 VSS CKN 10 VPW nch L=4e-08 W=1.3e-07 
M18 11 10 VSS VPW nch L=4e-08 W=1.3e-07 
M19 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M20 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M21 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M22 18 SE VDD VNW pch L=4e-08 W=3.8e-07 
M23 4 D 18 VNW pch L=4e-08 W=3.8e-07 
M24 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M25 19 11 5 VNW pch L=4e-08 W=1.5e-07 
M26 VDD 6 19 VNW pch L=4e-08 W=1.5e-07 
M27 6 SN VDD VNW pch L=4e-08 W=3.1e-07 
M28 VDD 5 6 VNW pch L=4e-08 W=3.1e-07 
M29 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M30 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M32 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M33 VDD 7 8 VNW pch L=4e-08 W=3.1e-07 
M34 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M36 VDD CKN 10 VNW pch L=4e-08 W=2.7e-07 
M37 11 10 VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFNSQ_X3M_A9TR Q VDD VNW VPW VSS CKN D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=1.3e-07 
M4 4 D 22 VPW nch L=4e-08 W=1.3e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.55e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.5e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.5e-07 
M8 24 SN VSS VPW nch L=4e-08 W=2.8e-07 
M9 6 5 24 VPW nch L=4e-08 W=2.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.55e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=3.8e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M16 VSS 8 Q VPW nch L=4e-08 W=2e-07 
M17 Q 8 VSS VPW nch L=4e-08 W=2e-07 
M18 VSS CKN 10 VPW nch L=4e-08 W=1.3e-07 
M19 11 10 VSS VPW nch L=4e-08 W=1.3e-07 
M20 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M21 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M22 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M23 18 SE VDD VNW pch L=4e-08 W=3.8e-07 
M24 4 D 18 VNW pch L=4e-08 W=3.8e-07 
M25 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M26 19 11 5 VNW pch L=4e-08 W=1.5e-07 
M27 VDD 6 19 VNW pch L=4e-08 W=1.5e-07 
M28 6 SN VDD VNW pch L=4e-08 W=3.1e-07 
M29 VDD 5 6 VNW pch L=4e-08 W=3.1e-07 
M30 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M31 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M32 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M33 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M34 VDD 7 8 VNW pch L=4e-08 W=3.8e-07 
M35 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M37 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M38 VDD CKN 10 VNW pch L=4e-08 W=2.7e-07 
M39 11 10 VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFNSRPQ_X1M_A9TR Q VDD VNW VPW VSS CKN D R SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 26 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M3 27 3 VSS VPW nch L=4e-08 W=1.2e-07 
M4 4 D 27 VPW nch L=4e-08 W=1.2e-07 
M5 5 12 4 VPW nch L=4e-08 W=1.2e-07 
M6 28 11 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 7 28 VPW nch L=4e-08 W=1.2e-07 
M8 6 SN VSS VPW nch L=4e-08 W=1.8e-07 
M9 7 5 6 VPW nch L=4e-08 W=1.8e-07 
M10 6 R 7 VPW nch L=4e-08 W=1.8e-07 
M11 8 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 29 12 8 VPW nch L=4e-08 W=1.6e-07 
M13 30 9 29 VPW nch L=4e-08 W=1.6e-07 
M14 VSS SN 30 VPW nch L=4e-08 W=1.6e-07 
M15 31 R VSS VPW nch L=4e-08 W=1.6e-07 
M16 8 SN 31 VPW nch L=4e-08 W=1.6e-07 
M17 VSS 8 9 VPW nch L=4e-08 W=2e-07 
M18 Q 9 VSS VPW nch L=4e-08 W=2e-07 
M19 VSS CKN 11 VPW nch L=4e-08 W=1.2e-07 
M20 12 11 VSS VPW nch L=4e-08 W=1.2e-07 
M21 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M22 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M23 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M24 20 SE VDD VNW pch L=4e-08 W=3.6e-07 
M25 4 D 20 VNW pch L=4e-08 W=3.6e-07 
M26 5 11 4 VNW pch L=4e-08 W=2e-07 
M27 21 12 5 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 7 21 VNW pch L=4e-08 W=1.2e-07 
M29 7 SN VDD VNW pch L=4e-08 W=3.6e-07 
M30 22 5 7 VNW pch L=4e-08 W=3.6e-07 
M31 VDD R 22 VNW pch L=4e-08 W=3.6e-07 
M32 8 12 7 VNW pch L=4e-08 W=2e-07 
M33 23 11 8 VNW pch L=4e-08 W=1.6e-07 
M34 24 9 23 VNW pch L=4e-08 W=1.6e-07 
M35 VDD R 24 VNW pch L=4e-08 W=1.6e-07 
M36 8 SN VDD VNW pch L=4e-08 W=1.6e-07 
M37 VDD 8 9 VNW pch L=4e-08 W=2e-07 
M38 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M39 VDD CKN 11 VNW pch L=4e-08 W=2.5e-07 
M40 12 11 VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFNSRPQ_X2M_A9TR Q VDD VNW VPW VSS CKN D R SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 26 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M3 27 3 VSS VPW nch L=4e-08 W=1.4e-07 
M4 4 D 27 VPW nch L=4e-08 W=1.4e-07 
M5 5 12 4 VPW nch L=4e-08 W=1.55e-07 
M6 28 11 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 7 28 VPW nch L=4e-08 W=1.2e-07 
M8 6 SN VSS VPW nch L=4e-08 W=1.8e-07 
M9 7 5 6 VPW nch L=4e-08 W=1.8e-07 
M10 6 R 7 VPW nch L=4e-08 W=1.8e-07 
M11 8 11 7 VPW nch L=4e-08 W=1.55e-07 
M12 29 12 8 VPW nch L=4e-08 W=1.6e-07 
M13 30 9 29 VPW nch L=4e-08 W=1.6e-07 
M14 VSS SN 30 VPW nch L=4e-08 W=1.6e-07 
M15 31 R VSS VPW nch L=4e-08 W=1.6e-07 
M16 8 SN 31 VPW nch L=4e-08 W=1.6e-07 
M17 VSS 8 9 VPW nch L=4e-08 W=3.1e-07 
M18 Q 9 VSS VPW nch L=4e-08 W=2e-07 
M19 VSS 9 Q VPW nch L=4e-08 W=2e-07 
M20 VSS CKN 11 VPW nch L=4e-08 W=1.3e-07 
M21 12 11 VSS VPW nch L=4e-08 W=1.3e-07 
M22 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M23 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M24 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M25 20 SE VDD VNW pch L=4e-08 W=3.8e-07 
M26 4 D 20 VNW pch L=4e-08 W=3.8e-07 
M27 5 11 4 VNW pch L=4e-08 W=3.1e-07 
M28 21 12 5 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 7 21 VNW pch L=4e-08 W=1.2e-07 
M30 7 SN VDD VNW pch L=4e-08 W=3.6e-07 
M31 22 5 7 VNW pch L=4e-08 W=3.6e-07 
M32 VDD R 22 VNW pch L=4e-08 W=3.6e-07 
M33 8 12 7 VNW pch L=4e-08 W=3.1e-07 
M34 23 11 8 VNW pch L=4e-08 W=1.6e-07 
M35 24 9 23 VNW pch L=4e-08 W=1.6e-07 
M36 VDD R 24 VNW pch L=4e-08 W=1.6e-07 
M37 8 SN VDD VNW pch L=4e-08 W=1.6e-07 
M38 VDD 8 9 VNW pch L=4e-08 W=3.1e-07 
M39 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M41 VDD CKN 11 VNW pch L=4e-08 W=2.7e-07 
M42 12 11 VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFNSRPQ_X3M_A9TR Q VDD VNW VPW VSS CKN D R SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 26 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M3 27 3 VSS VPW nch L=4e-08 W=1.4e-07 
M4 4 D 27 VPW nch L=4e-08 W=1.4e-07 
M5 5 12 4 VPW nch L=4e-08 W=1.55e-07 
M6 28 11 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 7 28 VPW nch L=4e-08 W=1.2e-07 
M8 6 SN VSS VPW nch L=4e-08 W=1.8e-07 
M9 7 5 6 VPW nch L=4e-08 W=1.8e-07 
M10 6 R 7 VPW nch L=4e-08 W=1.8e-07 
M11 8 11 7 VPW nch L=4e-08 W=1.55e-07 
M12 29 12 8 VPW nch L=4e-08 W=1.6e-07 
M13 30 9 29 VPW nch L=4e-08 W=1.6e-07 
M14 VSS SN 30 VPW nch L=4e-08 W=1.6e-07 
M15 31 R VSS VPW nch L=4e-08 W=1.6e-07 
M16 8 SN 31 VPW nch L=4e-08 W=1.6e-07 
M17 VSS 8 9 VPW nch L=4e-08 W=3.8e-07 
M18 Q 9 VSS VPW nch L=4e-08 W=2e-07 
M19 VSS 9 Q VPW nch L=4e-08 W=2e-07 
M20 Q 9 VSS VPW nch L=4e-08 W=2e-07 
M21 VSS CKN 11 VPW nch L=4e-08 W=1.3e-07 
M22 12 11 VSS VPW nch L=4e-08 W=1.3e-07 
M23 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M24 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M25 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M26 20 SE VDD VNW pch L=4e-08 W=3.8e-07 
M27 4 D 20 VNW pch L=4e-08 W=3.8e-07 
M28 5 11 4 VNW pch L=4e-08 W=3.1e-07 
M29 21 12 5 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 7 21 VNW pch L=4e-08 W=1.2e-07 
M31 7 SN VDD VNW pch L=4e-08 W=3.6e-07 
M32 22 5 7 VNW pch L=4e-08 W=3.6e-07 
M33 VDD R 22 VNW pch L=4e-08 W=3.6e-07 
M34 8 12 7 VNW pch L=4e-08 W=3.1e-07 
M35 23 11 8 VNW pch L=4e-08 W=1.6e-07 
M36 24 9 23 VNW pch L=4e-08 W=1.6e-07 
M37 VDD R 24 VNW pch L=4e-08 W=1.6e-07 
M38 8 SN VDD VNW pch L=4e-08 W=1.6e-07 
M39 VDD 8 9 VNW pch L=4e-08 W=3.8e-07 
M40 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M41 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M42 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M43 VDD CKN 11 VNW pch L=4e-08 W=2.7e-07 
M44 12 11 VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFQN_X0P5M_A9TR QN VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=1.8e-07 
M4 4 D 21 VPW nch L=4e-08 W=1.8e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.2e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M9 7 10 6 VPW nch L=4e-08 W=1.2e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M13 QN 7 VSS VPW nch L=4e-08 W=1.55e-07 
M14 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M15 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M16 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M17 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M18 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M19 17 SE VDD VNW pch L=4e-08 W=2.6e-07 
M20 4 D 17 VNW pch L=4e-08 W=2.6e-07 
M21 5 10 4 VNW pch L=4e-08 W=1.2e-07 
M22 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M24 6 5 VDD VNW pch L=4e-08 W=1.8e-07 
M25 7 11 6 VNW pch L=4e-08 W=1.2e-07 
M26 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M29 QN 7 VDD VNW pch L=4e-08 W=2e-07 
M30 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M31 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFQN_X1M_A9TR QN VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 4 D 21 VPW nch L=4e-08 W=2.4e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.6e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=1.6e-07 
M9 7 10 6 VPW nch L=4e-08 W=1.6e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M13 QN 7 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M15 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M16 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M17 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M18 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M19 17 SE VDD VNW pch L=4e-08 W=3.3e-07 
M20 4 D 17 VNW pch L=4e-08 W=3.3e-07 
M21 5 10 4 VNW pch L=4e-08 W=1.6e-07 
M22 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M24 6 5 VDD VNW pch L=4e-08 W=2.3e-07 
M25 7 11 6 VNW pch L=4e-08 W=1.6e-07 
M26 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M29 QN 7 VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M31 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFQN_X2M_A9TR QN VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 21 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=2.5e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=2.5e-07 
M9 7 10 6 VPW nch L=4e-08 W=2.5e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M13 QN 7 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 7 QN VPW nch L=4e-08 W=3.1e-07 
M15 VSS 11 10 VPW nch L=4e-08 W=1.3e-07 
M16 11 CK VSS VPW nch L=4e-08 W=1.3e-07 
M17 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M18 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M19 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M20 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M21 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M22 5 10 4 VNW pch L=4e-08 W=2.5e-07 
M23 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M25 6 5 VDD VNW pch L=4e-08 W=3.35e-07 
M26 7 11 6 VNW pch L=4e-08 W=2.5e-07 
M27 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M30 QN 7 VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD 7 QN VNW pch L=4e-08 W=3.8e-07 
M32 VDD 11 10 VNW pch L=4e-08 W=2.7e-07 
M33 11 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFQN_X3M_A9TR QN VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 21 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M13 QN 7 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 7 QN VPW nch L=4e-08 W=3.1e-07 
M15 QN 7 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.4e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.4e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M21 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M22 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M23 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M24 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M26 6 5 VDD VNW pch L=4e-08 W=3.8e-07 
M27 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M28 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M31 QN 7 VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD 7 QN VNW pch L=4e-08 W=3.8e-07 
M33 QN 7 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.9e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=1.8e-07 
M4 4 D 21 VPW nch L=4e-08 W=1.8e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.2e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=1.2e-07 
M9 7 10 6 VPW nch L=4e-08 W=1.2e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M13 Q 8 VSS VPW nch L=4e-08 W=1.55e-07 
M14 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M15 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M16 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M17 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M18 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M19 17 SE VDD VNW pch L=4e-08 W=2.5e-07 
M20 4 D 17 VNW pch L=4e-08 W=2.5e-07 
M21 5 10 4 VNW pch L=4e-08 W=1.2e-07 
M22 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M24 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M25 7 11 6 VNW pch L=4e-08 W=1.2e-07 
M26 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 7 8 VNW pch L=4e-08 W=1.55e-07 
M29 Q 8 VDD VNW pch L=4e-08 W=2e-07 
M30 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M31 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFQ_X1M_A9TR Q VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 4 D 21 VPW nch L=4e-08 W=2.4e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.6e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=1.6e-07 
M9 7 10 6 VPW nch L=4e-08 W=1.6e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 7 8 VPW nch L=4e-08 W=1.75e-07 
M13 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M15 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M16 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M17 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M18 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M19 17 SE VDD VNW pch L=4e-08 W=3.1e-07 
M20 4 D 17 VNW pch L=4e-08 W=3.1e-07 
M21 5 10 4 VNW pch L=4e-08 W=1.6e-07 
M22 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M23 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M24 6 5 VDD VNW pch L=4e-08 W=2.05e-07 
M25 7 11 6 VNW pch L=4e-08 W=1.6e-07 
M26 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 7 8 VNW pch L=4e-08 W=2.45e-07 
M29 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M31 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFQ_X2M_A9TR Q VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 21 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=2.5e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=2.5e-07 
M9 7 10 6 VPW nch L=4e-08 W=2.5e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 8 7 VSS VPW nch L=4e-08 W=2.5e-07 
M13 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M15 VSS 11 10 VPW nch L=4e-08 W=1.3e-07 
M16 11 CK VSS VPW nch L=4e-08 W=1.3e-07 
M17 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M18 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M19 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M20 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M21 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M22 5 10 4 VNW pch L=4e-08 W=2.5e-07 
M23 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M25 6 5 VDD VNW pch L=4e-08 W=3.25e-07 
M26 7 11 6 VNW pch L=4e-08 W=2.5e-07 
M27 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M29 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M30 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M32 VDD 11 10 VNW pch L=4e-08 W=2.7e-07 
M33 11 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFQ_X3M_A9TR Q VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 21 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 8 7 VSS VPW nch L=4e-08 W=2.5e-07 
M13 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.4e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.4e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M21 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M22 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M23 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M24 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M26 6 5 VDD VNW pch L=4e-08 W=3.8e-07 
M27 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M28 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M30 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M31 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M33 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.9e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFQ_X4M_A9TR Q VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 21 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 8 7 VSS VPW nch L=4e-08 W=2.5e-07 
M13 VSS 7 8 VPW nch L=4e-08 W=2.5e-07 
M14 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M16 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M18 VSS 11 10 VPW nch L=4e-08 W=1.4e-07 
M19 11 CK VSS VPW nch L=4e-08 W=1.4e-07 
M20 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M21 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M22 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M23 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M24 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M25 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M26 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M28 6 5 VDD VNW pch L=4e-08 W=3.8e-07 
M29 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M30 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M32 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD 7 8 VNW pch L=4e-08 W=3.8e-07 
M34 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M36 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M37 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M38 VDD 11 10 VNW pch L=4e-08 W=2.9e-07 
M39 11 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFRPQN_X0P5M_A9TR QN VDD VNW VPW VSS CK D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=1.8e-07 
M4 4 D 24 VPW nch L=4e-08 W=1.8e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.2e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=1.2e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.2e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 QN 7 VSS VPW nch L=4e-08 W=1.65e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=2.7e-07 
M22 4 D 18 VNW pch L=4e-08 W=2.7e-07 
M23 5 10 4 VNW pch L=4e-08 W=1.2e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M26 20 R VDD VNW pch L=4e-08 W=2.7e-07 
M27 6 5 20 VNW pch L=4e-08 W=2.7e-07 
M28 7 11 6 VNW pch L=4e-08 W=1.2e-07 
M29 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M30 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M31 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M33 QN 7 VDD VNW pch L=4e-08 W=1.8e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFRPQN_X1M_A9TR QN VDD VNW VPW VSS CK D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 4 D 24 VPW nch L=4e-08 W=2.4e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.5e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=1.5e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=1.5e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.5e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 QN 7 VSS VPW nch L=4e-08 W=3.3e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=3.3e-07 
M22 4 D 18 VNW pch L=4e-08 W=3.3e-07 
M23 5 10 4 VNW pch L=4e-08 W=1.7e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M26 20 R VDD VNW pch L=4e-08 W=3.3e-07 
M27 6 5 20 VNW pch L=4e-08 W=3.3e-07 
M28 7 11 6 VNW pch L=4e-08 W=1.7e-07 
M29 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M30 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M31 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M33 QN 7 VDD VNW pch L=4e-08 W=3.6e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFRPQN_X2M_A9TR QN VDD VNW VPW VSS CK D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=3.3e-07 
M4 4 D 24 VPW nch L=4e-08 W=3.3e-07 
M5 5 11 4 VPW nch L=4e-08 W=2e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=2e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=2e-07 
M10 7 10 6 VPW nch L=4e-08 W=2e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 QN 7 VSS VPW nch L=4e-08 W=3.3e-07 
M16 VSS 7 QN VPW nch L=4e-08 W=3.3e-07 
M17 VSS 11 10 VPW nch L=4e-08 W=1.3e-07 
M18 11 CK VSS VPW nch L=4e-08 W=1.3e-07 
M19 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M20 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M21 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M22 18 SE VDD VNW pch L=4e-08 W=3.6e-07 
M23 4 D 18 VNW pch L=4e-08 W=3.6e-07 
M24 5 10 4 VNW pch L=4e-08 W=3e-07 
M25 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M27 20 R VDD VNW pch L=4e-08 W=3.8e-07 
M28 6 5 20 VNW pch L=4e-08 W=3.8e-07 
M29 7 11 6 VNW pch L=4e-08 W=3e-07 
M30 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M31 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M32 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M33 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M34 QN 7 VDD VNW pch L=4e-08 W=3.6e-07 
M35 VDD 7 QN VNW pch L=4e-08 W=3.6e-07 
M36 VDD 11 10 VNW pch L=4e-08 W=2.7e-07 
M37 11 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFRPQN_X3M_A9TR QN VDD VNW VPW VSS CK D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=3.3e-07 
M4 4 D 24 VPW nch L=4e-08 W=3.3e-07 
M5 5 11 4 VPW nch L=4e-08 W=2e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=2e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=2e-07 
M10 7 10 6 VPW nch L=4e-08 W=2e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 QN 7 VSS VPW nch L=4e-08 W=3.4e-07 
M16 VSS 7 QN VPW nch L=4e-08 W=3.4e-07 
M17 QN 7 VSS VPW nch L=4e-08 W=3.4e-07 
M18 VSS 11 10 VPW nch L=4e-08 W=1.3e-07 
M19 11 CK VSS VPW nch L=4e-08 W=1.3e-07 
M20 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M21 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M22 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M23 18 SE VDD VNW pch L=4e-08 W=3.6e-07 
M24 4 D 18 VNW pch L=4e-08 W=3.6e-07 
M25 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M26 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M28 20 R VDD VNW pch L=4e-08 W=3.8e-07 
M29 6 5 20 VNW pch L=4e-08 W=3.8e-07 
M30 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M31 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M32 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M33 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M34 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M35 QN 7 VDD VNW pch L=4e-08 W=3.5e-07 
M36 VDD 7 QN VNW pch L=4e-08 W=3.5e-07 
M37 QN 7 VDD VNW pch L=4e-08 W=3.5e-07 
M38 VDD 11 10 VNW pch L=4e-08 W=2.7e-07 
M39 11 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFRPQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=1.8e-07 
M4 4 D 24 VPW nch L=4e-08 W=1.8e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.2e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=1.2e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=1.2e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.2e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=1.55e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=2.5e-07 
M22 4 D 18 VNW pch L=4e-08 W=2.5e-07 
M23 5 10 4 VNW pch L=4e-08 W=1.2e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M26 20 R VDD VNW pch L=4e-08 W=2.5e-07 
M27 6 5 20 VNW pch L=4e-08 W=2.5e-07 
M28 7 11 6 VNW pch L=4e-08 W=1.2e-07 
M29 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M30 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M31 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=1.35e-07 
M33 Q 8 VDD VNW pch L=4e-08 W=2e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFRPQ_X1M_A9TR Q VDD VNW VPW VSS CK D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 4 D 24 VPW nch L=4e-08 W=2.4e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.6e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=1.6e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=1.6e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.55e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.95e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=3.1e-07 
M22 4 D 18 VNW pch L=4e-08 W=3.1e-07 
M23 5 10 4 VNW pch L=4e-08 W=1.6e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M26 20 R VDD VNW pch L=4e-08 W=3.2e-07 
M27 6 5 20 VNW pch L=4e-08 W=3.2e-07 
M28 7 11 6 VNW pch L=4e-08 W=1.55e-07 
M29 21 10 7 VNW pch L=4e-08 W=1.55e-07 
M30 22 8 21 VNW pch L=4e-08 W=1.55e-07 
M31 VDD R 22 VNW pch L=4e-08 W=1.55e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=2.25e-07 
M33 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFRPQ_X2M_A9TR Q VDD VNW VPW VSS CK D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=3.3e-07 
M4 4 D 24 VPW nch L=4e-08 W=3.3e-07 
M5 5 11 4 VPW nch L=4e-08 W=2.5e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=2.5e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=2.5e-07 
M10 7 10 6 VPW nch L=4e-08 W=2.5e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=3e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M17 VSS 11 10 VPW nch L=4e-08 W=1.3e-07 
M18 11 CK VSS VPW nch L=4e-08 W=1.3e-07 
M19 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M20 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M21 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M22 18 SE VDD VNW pch L=4e-08 W=3.6e-07 
M23 4 D 18 VNW pch L=4e-08 W=3.6e-07 
M24 5 10 4 VNW pch L=4e-08 W=2.5e-07 
M25 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M27 20 R VDD VNW pch L=4e-08 W=3.8e-07 
M28 6 5 20 VNW pch L=4e-08 W=3.8e-07 
M29 7 11 6 VNW pch L=4e-08 W=2.5e-07 
M30 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M31 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M32 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M33 VDD 7 8 VNW pch L=4e-08 W=3.4e-07 
M34 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M36 VDD 11 10 VNW pch L=4e-08 W=2.7e-07 
M37 11 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFRPQ_X3M_A9TR Q VDD VNW VPW VSS CK D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=3.3e-07 
M4 4 D 24 VPW nch L=4e-08 W=3.3e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=2.5e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=2.5e-07 
M10 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=3.4e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M17 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M18 VSS 11 10 VPW nch L=4e-08 W=1.4e-07 
M19 11 CK VSS VPW nch L=4e-08 W=1.4e-07 
M20 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M21 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M22 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M23 18 SE VDD VNW pch L=4e-08 W=3.6e-07 
M24 4 D 18 VNW pch L=4e-08 W=3.6e-07 
M25 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M26 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M28 20 R VDD VNW pch L=4e-08 W=3.8e-07 
M29 6 5 20 VNW pch L=4e-08 W=3.8e-07 
M30 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M31 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M32 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M33 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M34 VDD 7 8 VNW pch L=4e-08 W=3.8e-07 
M35 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M37 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M38 VDD 11 10 VNW pch L=4e-08 W=2.9e-07 
M39 11 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFRPQ_X4M_A9TR Q VDD VNW VPW VSS CK D R SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 23 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 23 VPW nch L=4e-08 W=1.2e-07 
M3 24 3 VSS VPW nch L=4e-08 W=3.3e-07 
M4 4 D 24 VPW nch L=4e-08 W=3.3e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 25 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 25 VPW nch L=4e-08 W=1.2e-07 
M8 6 R VSS VPW nch L=4e-08 W=2.5e-07 
M9 VSS 5 6 VPW nch L=4e-08 W=2.5e-07 
M10 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M11 26 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 VSS 8 26 VPW nch L=4e-08 W=1.2e-07 
M13 7 R VSS VPW nch L=4e-08 W=1.2e-07 
M14 8 7 VSS VPW nch L=4e-08 W=3e-07 
M15 VSS 7 8 VPW nch L=4e-08 W=3e-07 
M16 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M18 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M20 VSS 11 10 VPW nch L=4e-08 W=1.4e-07 
M21 11 CK VSS VPW nch L=4e-08 W=1.4e-07 
M22 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M23 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M24 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M25 18 SE VDD VNW pch L=4e-08 W=3.6e-07 
M26 4 D 18 VNW pch L=4e-08 W=3.6e-07 
M27 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M28 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M30 20 R VDD VNW pch L=4e-08 W=3.8e-07 
M31 6 5 20 VNW pch L=4e-08 W=3.8e-07 
M32 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M33 21 10 7 VNW pch L=4e-08 W=1.6e-07 
M34 22 8 21 VNW pch L=4e-08 W=1.6e-07 
M35 VDD R 22 VNW pch L=4e-08 W=1.6e-07 
M36 8 7 VDD VNW pch L=4e-08 W=3.2e-07 
M37 VDD 7 8 VNW pch L=4e-08 W=3.2e-07 
M38 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M39 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M40 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M41 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M42 VDD 11 10 VNW pch L=4e-08 W=2.9e-07 
M43 11 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFSQN_X0P5M_A9TR QN VDD VNW VPW VSS CK D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=1.8e-07 
M4 4 D 22 VPW nch L=4e-08 W=1.8e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.2e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.2e-07 
M8 24 5 VSS VPW nch L=4e-08 W=1.8e-07 
M9 6 SN 24 VPW nch L=4e-08 W=1.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.2e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 QN 7 VSS VPW nch L=4e-08 W=1.55e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=2.6e-07 
M22 4 D 18 VNW pch L=4e-08 W=2.6e-07 
M23 5 10 4 VNW pch L=4e-08 W=1.2e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M26 6 5 VDD VNW pch L=4e-08 W=1.55e-07 
M27 VDD SN 6 VNW pch L=4e-08 W=1.55e-07 
M28 7 11 6 VNW pch L=4e-08 W=1.2e-07 
M29 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M31 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M33 QN 7 VDD VNW pch L=4e-08 W=2e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFSQN_X1M_A9TR QN VDD VNW VPW VSS CK D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 4 D 22 VPW nch L=4e-08 W=2.4e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.6e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.2e-07 
M8 24 5 VSS VPW nch L=4e-08 W=2.45e-07 
M9 6 SN 24 VPW nch L=4e-08 W=2.45e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.6e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 QN 7 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=3.2e-07 
M22 4 D 18 VNW pch L=4e-08 W=3.2e-07 
M23 5 10 4 VNW pch L=4e-08 W=1.6e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M26 6 5 VDD VNW pch L=4e-08 W=2.05e-07 
M27 VDD SN 6 VNW pch L=4e-08 W=2.05e-07 
M28 7 11 6 VNW pch L=4e-08 W=1.6e-07 
M29 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M31 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M33 QN 7 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFSQN_X2M_A9TR QN VDD VNW VPW VSS CK D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 22 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=2.5e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.2e-07 
M8 24 5 VSS VPW nch L=4e-08 W=3.8e-07 
M9 6 SN 24 VPW nch L=4e-08 W=3.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=2.5e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 QN 7 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 7 QN VPW nch L=4e-08 W=3.1e-07 
M17 VSS 11 10 VPW nch L=4e-08 W=1.3e-07 
M18 11 CK VSS VPW nch L=4e-08 W=1.3e-07 
M19 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M20 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M21 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M22 18 SE VDD VNW pch L=4e-08 W=3.8e-07 
M23 4 D 18 VNW pch L=4e-08 W=3.8e-07 
M24 5 10 4 VNW pch L=4e-08 W=2.5e-07 
M25 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M27 6 5 VDD VNW pch L=4e-08 W=3.2e-07 
M28 VDD SN 6 VNW pch L=4e-08 W=3.2e-07 
M29 7 11 6 VNW pch L=4e-08 W=2.5e-07 
M30 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M32 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M33 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M34 QN 7 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 7 QN VNW pch L=4e-08 W=3.8e-07 
M36 VDD 11 10 VNW pch L=4e-08 W=2.7e-07 
M37 11 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFSQN_X3M_A9TR QN VDD VNW VPW VSS CK D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 22 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.2e-07 
M8 24 5 VSS VPW nch L=4e-08 W=3.8e-07 
M9 6 SN 24 VPW nch L=4e-08 W=3.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 QN 7 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 7 QN VPW nch L=4e-08 W=3.1e-07 
M17 QN 7 VSS VPW nch L=4e-08 W=3.1e-07 
M18 VSS 11 10 VPW nch L=4e-08 W=1.4e-07 
M19 11 CK VSS VPW nch L=4e-08 W=1.4e-07 
M20 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M21 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M22 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M23 18 SE VDD VNW pch L=4e-08 W=3.8e-07 
M24 4 D 18 VNW pch L=4e-08 W=3.8e-07 
M25 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M26 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M28 6 5 VDD VNW pch L=4e-08 W=3.2e-07 
M29 VDD SN 6 VNW pch L=4e-08 W=3.2e-07 
M30 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M31 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M32 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M33 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M34 VDD 7 8 VNW pch L=4e-08 W=1.2e-07 
M35 QN 7 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 7 QN VNW pch L=4e-08 W=3.8e-07 
M37 QN 7 VDD VNW pch L=4e-08 W=3.8e-07 
M38 VDD 11 10 VNW pch L=4e-08 W=2.9e-07 
M39 11 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFSQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=1.8e-07 
M4 4 D 22 VPW nch L=4e-08 W=1.8e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.2e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.2e-07 
M8 24 SN VSS VPW nch L=4e-08 W=1.8e-07 
M9 6 5 24 VPW nch L=4e-08 W=1.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.2e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.2e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=1.55e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=2.6e-07 
M22 4 D 18 VNW pch L=4e-08 W=2.6e-07 
M23 5 10 4 VNW pch L=4e-08 W=1.2e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M26 6 SN VDD VNW pch L=4e-08 W=1.55e-07 
M27 VDD 5 6 VNW pch L=4e-08 W=1.55e-07 
M28 7 11 6 VNW pch L=4e-08 W=1.2e-07 
M29 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M31 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=1.6e-07 
M33 Q 8 VDD VNW pch L=4e-08 W=2e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFSQ_X1M_A9TR Q VDD VNW VPW VSS CK D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 4 D 22 VPW nch L=4e-08 W=2.4e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.6e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.2e-07 
M8 24 SN VSS VPW nch L=4e-08 W=2.4e-07 
M9 6 5 24 VPW nch L=4e-08 W=2.4e-07 
M10 7 10 6 VPW nch L=4e-08 W=1.6e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=1.65e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=1.2e-07 
M17 11 CK VSS VPW nch L=4e-08 W=1.2e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M21 18 SE VDD VNW pch L=4e-08 W=3.2e-07 
M22 4 D 18 VNW pch L=4e-08 W=3.2e-07 
M23 5 10 4 VNW pch L=4e-08 W=1.6e-07 
M24 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M26 6 SN VDD VNW pch L=4e-08 W=2.05e-07 
M27 VDD 5 6 VNW pch L=4e-08 W=2.05e-07 
M28 7 11 6 VNW pch L=4e-08 W=1.6e-07 
M29 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M31 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M32 VDD 7 8 VNW pch L=4e-08 W=2.55e-07 
M33 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=2.5e-07 
M35 11 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFSQ_X2M_A9TR Q VDD VNW VPW VSS CK D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 22 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=2.5e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.2e-07 
M8 24 SN VSS VPW nch L=4e-08 W=3.8e-07 
M9 6 5 24 VPW nch L=4e-08 W=3.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=2.5e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=2.5e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M17 VSS 11 10 VPW nch L=4e-08 W=1.3e-07 
M18 11 CK VSS VPW nch L=4e-08 W=1.3e-07 
M19 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M20 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M21 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M22 18 SE VDD VNW pch L=4e-08 W=3.8e-07 
M23 4 D 18 VNW pch L=4e-08 W=3.8e-07 
M24 5 10 4 VNW pch L=4e-08 W=2.5e-07 
M25 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M26 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M27 6 SN VDD VNW pch L=4e-08 W=3.25e-07 
M28 VDD 5 6 VNW pch L=4e-08 W=3.25e-07 
M29 7 11 6 VNW pch L=4e-08 W=2.5e-07 
M30 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M32 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M33 VDD 7 8 VNW pch L=4e-08 W=3.8e-07 
M34 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M36 VDD 11 10 VNW pch L=4e-08 W=2.7e-07 
M37 11 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFSQ_X3M_A9TR Q VDD VNW VPW VSS CK D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 22 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.2e-07 
M8 24 SN VSS VPW nch L=4e-08 W=3.8e-07 
M9 6 5 24 VPW nch L=4e-08 W=3.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 VSS 7 8 VPW nch L=4e-08 W=2.5e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M17 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M18 VSS 11 10 VPW nch L=4e-08 W=1.4e-07 
M19 11 CK VSS VPW nch L=4e-08 W=1.4e-07 
M20 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M21 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M22 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M23 18 SE VDD VNW pch L=4e-08 W=3.8e-07 
M24 4 D 18 VNW pch L=4e-08 W=3.8e-07 
M25 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M26 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M28 6 SN VDD VNW pch L=4e-08 W=3.25e-07 
M29 VDD 5 6 VNW pch L=4e-08 W=3.25e-07 
M30 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M31 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M32 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M33 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M34 VDD 7 8 VNW pch L=4e-08 W=3.8e-07 
M35 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M37 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M38 VDD 11 10 VNW pch L=4e-08 W=2.9e-07 
M39 11 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFSQ_X4M_A9TR Q VDD VNW VPW VSS CK D SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 21 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 21 VPW nch L=4e-08 W=1.2e-07 
M3 22 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 22 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 23 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 23 VPW nch L=4e-08 W=1.2e-07 
M8 24 SN VSS VPW nch L=4e-08 W=3.8e-07 
M9 6 5 24 VPW nch L=4e-08 W=3.8e-07 
M10 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M11 25 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 26 8 25 VPW nch L=4e-08 W=1.6e-07 
M13 VSS SN 26 VPW nch L=4e-08 W=1.6e-07 
M14 8 7 VSS VPW nch L=4e-08 W=1.9e-07 
M15 VSS 7 8 VPW nch L=4e-08 W=1.9e-07 
M16 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M18 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M20 VSS 11 10 VPW nch L=4e-08 W=1.4e-07 
M21 11 CK VSS VPW nch L=4e-08 W=1.4e-07 
M22 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M23 17 3 4 VNW pch L=4e-08 W=1.55e-07 
M24 VDD SI 17 VNW pch L=4e-08 W=1.55e-07 
M25 18 SE VDD VNW pch L=4e-08 W=3.8e-07 
M26 4 D 18 VNW pch L=4e-08 W=3.8e-07 
M27 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M28 19 11 5 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 6 19 VNW pch L=4e-08 W=1.2e-07 
M30 6 SN VDD VNW pch L=4e-08 W=3.25e-07 
M31 VDD 5 6 VNW pch L=4e-08 W=3.25e-07 
M32 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M33 20 10 7 VNW pch L=4e-08 W=1.2e-07 
M34 VDD 8 20 VNW pch L=4e-08 W=1.2e-07 
M35 7 SN VDD VNW pch L=4e-08 W=1.2e-07 
M36 8 7 VDD VNW pch L=4e-08 W=3.4e-07 
M37 VDD 7 8 VNW pch L=4e-08 W=3.4e-07 
M38 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M39 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M40 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M41 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M42 VDD 11 10 VNW pch L=4e-08 W=2.9e-07 
M43 11 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFSRPQ_X0P5M_A9TR Q VDD VNW VPW VSS CK D R SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 26 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M3 27 3 VSS VPW nch L=4e-08 W=1.8e-07 
M4 4 D 27 VPW nch L=4e-08 W=1.8e-07 
M5 5 12 4 VPW nch L=4e-08 W=1.2e-07 
M6 28 11 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 7 28 VPW nch L=4e-08 W=1.2e-07 
M8 6 SN VSS VPW nch L=4e-08 W=1.8e-07 
M9 7 5 6 VPW nch L=4e-08 W=1.8e-07 
M10 6 R 7 VPW nch L=4e-08 W=1.8e-07 
M11 8 11 7 VPW nch L=4e-08 W=1.2e-07 
M12 29 12 8 VPW nch L=4e-08 W=1.6e-07 
M13 30 9 29 VPW nch L=4e-08 W=1.6e-07 
M14 VSS SN 30 VPW nch L=4e-08 W=1.6e-07 
M15 31 R VSS VPW nch L=4e-08 W=1.6e-07 
M16 8 SN 31 VPW nch L=4e-08 W=1.6e-07 
M17 VSS 8 9 VPW nch L=4e-08 W=1.2e-07 
M18 Q 9 VSS VPW nch L=4e-08 W=1.55e-07 
M19 VSS 12 11 VPW nch L=4e-08 W=1.2e-07 
M20 12 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M22 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M23 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M24 20 SE VDD VNW pch L=4e-08 W=2.6e-07 
M25 4 D 20 VNW pch L=4e-08 W=2.6e-07 
M26 5 11 4 VNW pch L=4e-08 W=1.2e-07 
M27 21 12 5 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 7 21 VNW pch L=4e-08 W=1.2e-07 
M29 7 SN VDD VNW pch L=4e-08 W=2.6e-07 
M30 22 5 7 VNW pch L=4e-08 W=2.6e-07 
M31 VDD R 22 VNW pch L=4e-08 W=2.6e-07 
M32 8 12 7 VNW pch L=4e-08 W=1.2e-07 
M33 23 11 8 VNW pch L=4e-08 W=1.6e-07 
M34 24 9 23 VNW pch L=4e-08 W=1.6e-07 
M35 VDD R 24 VNW pch L=4e-08 W=1.6e-07 
M36 8 SN VDD VNW pch L=4e-08 W=1.6e-07 
M37 VDD 8 9 VNW pch L=4e-08 W=1.3e-07 
M38 Q 9 VDD VNW pch L=4e-08 W=2e-07 
M39 VDD 12 11 VNW pch L=4e-08 W=2.5e-07 
M40 12 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFSRPQ_X1M_A9TR Q VDD VNW VPW VSS CK D R SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 26 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M3 27 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 4 D 27 VPW nch L=4e-08 W=2.4e-07 
M5 5 12 4 VPW nch L=4e-08 W=1.6e-07 
M6 28 11 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 7 28 VPW nch L=4e-08 W=1.2e-07 
M8 6 SN VSS VPW nch L=4e-08 W=2.4e-07 
M9 7 5 6 VPW nch L=4e-08 W=2.4e-07 
M10 6 R 7 VPW nch L=4e-08 W=2.4e-07 
M11 8 11 7 VPW nch L=4e-08 W=1.6e-07 
M12 29 12 8 VPW nch L=4e-08 W=1.6e-07 
M13 30 9 29 VPW nch L=4e-08 W=1.6e-07 
M14 VSS SN 30 VPW nch L=4e-08 W=1.6e-07 
M15 31 R VSS VPW nch L=4e-08 W=1.6e-07 
M16 8 SN 31 VPW nch L=4e-08 W=1.6e-07 
M17 VSS 8 9 VPW nch L=4e-08 W=2e-07 
M18 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 12 11 VPW nch L=4e-08 W=1.2e-07 
M20 12 CK VSS VPW nch L=4e-08 W=1.2e-07 
M21 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M22 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M23 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M24 20 SE VDD VNW pch L=4e-08 W=3.1e-07 
M25 4 D 20 VNW pch L=4e-08 W=3.1e-07 
M26 5 11 4 VNW pch L=4e-08 W=1.6e-07 
M27 21 12 5 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 7 21 VNW pch L=4e-08 W=1.2e-07 
M29 7 SN VDD VNW pch L=4e-08 W=3.2e-07 
M30 22 5 7 VNW pch L=4e-08 W=3.2e-07 
M31 VDD R 22 VNW pch L=4e-08 W=3.2e-07 
M32 8 12 7 VNW pch L=4e-08 W=1.6e-07 
M33 23 11 8 VNW pch L=4e-08 W=1.6e-07 
M34 24 9 23 VNW pch L=4e-08 W=1.6e-07 
M35 VDD R 24 VNW pch L=4e-08 W=1.6e-07 
M36 8 SN VDD VNW pch L=4e-08 W=1.6e-07 
M37 VDD 8 9 VNW pch L=4e-08 W=2.2e-07 
M38 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M39 VDD 12 11 VNW pch L=4e-08 W=2.5e-07 
M40 12 CK VDD VNW pch L=4e-08 W=1.3e-07 
.ENDS


.SUBCKT SDFFSRPQ_X2M_A9TR Q VDD VNW VPW VSS CK D R SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 26 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M3 27 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 27 VPW nch L=4e-08 W=3.1e-07 
M5 5 12 4 VPW nch L=4e-08 W=2.5e-07 
M6 28 11 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 7 28 VPW nch L=4e-08 W=1.2e-07 
M8 6 SN VSS VPW nch L=4e-08 W=2.95e-07 
M9 7 5 6 VPW nch L=4e-08 W=2.95e-07 
M10 6 R 7 VPW nch L=4e-08 W=2.95e-07 
M11 8 11 7 VPW nch L=4e-08 W=2.5e-07 
M12 29 12 8 VPW nch L=4e-08 W=1.6e-07 
M13 30 9 29 VPW nch L=4e-08 W=1.6e-07 
M14 VSS SN 30 VPW nch L=4e-08 W=1.6e-07 
M15 31 R VSS VPW nch L=4e-08 W=1.6e-07 
M16 8 SN 31 VPW nch L=4e-08 W=1.6e-07 
M17 VSS 8 9 VPW nch L=4e-08 W=3e-07 
M18 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M20 VSS 12 11 VPW nch L=4e-08 W=1.3e-07 
M21 12 CK VSS VPW nch L=4e-08 W=1.3e-07 
M22 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M23 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M24 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M25 20 SE VDD VNW pch L=4e-08 W=3.8e-07 
M26 4 D 20 VNW pch L=4e-08 W=3.8e-07 
M27 5 11 4 VNW pch L=4e-08 W=2.5e-07 
M28 21 12 5 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 7 21 VNW pch L=4e-08 W=1.2e-07 
M30 7 SN VDD VNW pch L=4e-08 W=3.8e-07 
M31 22 5 7 VNW pch L=4e-08 W=3.8e-07 
M32 VDD R 22 VNW pch L=4e-08 W=3.8e-07 
M33 8 12 7 VNW pch L=4e-08 W=2.5e-07 
M34 23 11 8 VNW pch L=4e-08 W=1.6e-07 
M35 24 9 23 VNW pch L=4e-08 W=1.6e-07 
M36 VDD R 24 VNW pch L=4e-08 W=1.6e-07 
M37 8 SN VDD VNW pch L=4e-08 W=1.6e-07 
M38 VDD 8 9 VNW pch L=4e-08 W=3.35e-07 
M39 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M41 VDD 12 11 VNW pch L=4e-08 W=2.7e-07 
M42 12 CK VDD VNW pch L=4e-08 W=1.4e-07 
.ENDS


.SUBCKT SDFFSRPQ_X3M_A9TR Q VDD VNW VPW VSS CK D R SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 26 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M3 27 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 27 VPW nch L=4e-08 W=3.1e-07 
M5 5 12 4 VPW nch L=4e-08 W=3.1e-07 
M6 28 11 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 7 28 VPW nch L=4e-08 W=1.2e-07 
M8 6 SN VSS VPW nch L=4e-08 W=2.95e-07 
M9 7 5 6 VPW nch L=4e-08 W=2.95e-07 
M10 6 R 7 VPW nch L=4e-08 W=2.95e-07 
M11 8 11 7 VPW nch L=4e-08 W=3.1e-07 
M12 29 12 8 VPW nch L=4e-08 W=1.6e-07 
M13 30 9 29 VPW nch L=4e-08 W=1.6e-07 
M14 VSS SN 30 VPW nch L=4e-08 W=1.6e-07 
M15 31 R VSS VPW nch L=4e-08 W=1.6e-07 
M16 8 SN 31 VPW nch L=4e-08 W=1.6e-07 
M17 VSS 8 9 VPW nch L=4e-08 W=3.1e-07 
M18 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M20 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M21 VSS 12 11 VPW nch L=4e-08 W=1.4e-07 
M22 12 CK VSS VPW nch L=4e-08 W=1.4e-07 
M23 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M24 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M25 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M26 20 SE VDD VNW pch L=4e-08 W=3.8e-07 
M27 4 D 20 VNW pch L=4e-08 W=3.8e-07 
M28 5 11 4 VNW pch L=4e-08 W=3.1e-07 
M29 21 12 5 VNW pch L=4e-08 W=1.2e-07 
M30 VDD 7 21 VNW pch L=4e-08 W=1.2e-07 
M31 7 SN VDD VNW pch L=4e-08 W=3.8e-07 
M32 22 5 7 VNW pch L=4e-08 W=3.8e-07 
M33 VDD R 22 VNW pch L=4e-08 W=3.8e-07 
M34 8 12 7 VNW pch L=4e-08 W=3.1e-07 
M35 23 11 8 VNW pch L=4e-08 W=1.6e-07 
M36 24 9 23 VNW pch L=4e-08 W=1.6e-07 
M37 VDD R 24 VNW pch L=4e-08 W=1.6e-07 
M38 8 SN VDD VNW pch L=4e-08 W=1.6e-07 
M39 VDD 8 9 VNW pch L=4e-08 W=3.8e-07 
M40 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M41 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M42 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M43 VDD 12 11 VNW pch L=4e-08 W=2.9e-07 
M44 12 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFSRPQ_X4M_A9TR Q VDD VNW VPW VSS CK D R SE SI SN
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 26 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 26 VPW nch L=4e-08 W=1.2e-07 
M3 27 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 27 VPW nch L=4e-08 W=3.1e-07 
M5 5 12 4 VPW nch L=4e-08 W=3.1e-07 
M6 28 11 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 7 28 VPW nch L=4e-08 W=1.2e-07 
M8 6 SN VSS VPW nch L=4e-08 W=2.95e-07 
M9 7 5 6 VPW nch L=4e-08 W=2.95e-07 
M10 6 R 7 VPW nch L=4e-08 W=2.95e-07 
M11 8 11 7 VPW nch L=4e-08 W=3.1e-07 
M12 29 12 8 VPW nch L=4e-08 W=1.6e-07 
M13 30 9 29 VPW nch L=4e-08 W=1.6e-07 
M14 VSS SN 30 VPW nch L=4e-08 W=1.6e-07 
M15 31 R VSS VPW nch L=4e-08 W=1.6e-07 
M16 8 SN 31 VPW nch L=4e-08 W=1.6e-07 
M17 9 8 VSS VPW nch L=4e-08 W=3e-07 
M18 VSS 8 9 VPW nch L=4e-08 W=3e-07 
M19 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M20 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M21 Q 9 VSS VPW nch L=4e-08 W=3.1e-07 
M22 VSS 9 Q VPW nch L=4e-08 W=3.1e-07 
M23 VSS 12 11 VPW nch L=4e-08 W=1.4e-07 
M24 12 CK VSS VPW nch L=4e-08 W=1.4e-07 
M25 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M26 19 3 4 VNW pch L=4e-08 W=1.55e-07 
M27 VDD SI 19 VNW pch L=4e-08 W=1.55e-07 
M28 20 SE VDD VNW pch L=4e-08 W=3.8e-07 
M29 4 D 20 VNW pch L=4e-08 W=3.8e-07 
M30 5 11 4 VNW pch L=4e-08 W=3.1e-07 
M31 21 12 5 VNW pch L=4e-08 W=1.2e-07 
M32 VDD 7 21 VNW pch L=4e-08 W=1.2e-07 
M33 7 SN VDD VNW pch L=4e-08 W=3.8e-07 
M34 22 5 7 VNW pch L=4e-08 W=3.8e-07 
M35 VDD R 22 VNW pch L=4e-08 W=3.8e-07 
M36 8 12 7 VNW pch L=4e-08 W=3.1e-07 
M37 23 11 8 VNW pch L=4e-08 W=1.6e-07 
M38 24 9 23 VNW pch L=4e-08 W=1.6e-07 
M39 VDD R 24 VNW pch L=4e-08 W=1.6e-07 
M40 8 SN VDD VNW pch L=4e-08 W=1.6e-07 
M41 9 8 VDD VNW pch L=4e-08 W=3.2e-07 
M42 VDD 8 9 VNW pch L=4e-08 W=3.2e-07 
M43 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M44 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M45 Q 9 VDD VNW pch L=4e-08 W=3.8e-07 
M46 VDD 9 Q VNW pch L=4e-08 W=3.8e-07 
M47 VDD 12 11 VNW pch L=4e-08 W=2.9e-07 
M48 12 CK VDD VNW pch L=4e-08 W=1.5e-07 
.ENDS


.SUBCKT SDFFYQ_X1M_A9TR Q VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=2.4e-07 
M4 4 D 21 VPW nch L=4e-08 W=2.4e-07 
M5 5 11 4 VPW nch L=4e-08 W=1.6e-07 
M6 22 10 5 VPW nch L=4e-08 W=2.4e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=2.4e-07 
M8 6 5 VSS VPW nch L=4e-08 W=1.6e-07 
M9 7 10 6 VPW nch L=4e-08 W=1.6e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.6e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.6e-07 
M12 VSS 7 8 VPW nch L=4e-08 W=1.9e-07 
M13 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 11 10 VPW nch L=4e-08 W=2.2e-07 
M15 11 CK VSS VPW nch L=4e-08 W=2.2e-07 
M16 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M17 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M18 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M19 17 SE VDD VNW pch L=4e-08 W=3.3e-07 
M20 4 D 17 VNW pch L=4e-08 W=3.3e-07 
M21 5 10 4 VNW pch L=4e-08 W=1.6e-07 
M22 18 11 5 VNW pch L=4e-08 W=2.4e-07 
M23 VDD 6 18 VNW pch L=4e-08 W=2.4e-07 
M24 6 5 VDD VNW pch L=4e-08 W=2.05e-07 
M25 7 11 6 VNW pch L=4e-08 W=1.6e-07 
M26 19 10 7 VNW pch L=4e-08 W=2.4e-07 
M27 VDD 8 19 VNW pch L=4e-08 W=2.4e-07 
M28 VDD 7 8 VNW pch L=4e-08 W=2.3e-07 
M29 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD 11 10 VNW pch L=4e-08 W=3.3e-07 
M31 11 CK VDD VNW pch L=4e-08 W=2.4e-07 
.ENDS


.SUBCKT SDFFYQ_X2M_A9TR Q VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 21 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=2.5e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=2.5e-07 
M9 7 10 6 VPW nch L=4e-08 W=2.5e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 8 7 VSS VPW nch L=4e-08 W=2.5e-07 
M13 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M15 VSS 11 10 VPW nch L=4e-08 W=2.3e-07 
M16 11 CK VSS VPW nch L=4e-08 W=2.3e-07 
M17 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M18 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M19 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M20 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M21 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M22 5 10 4 VNW pch L=4e-08 W=2.5e-07 
M23 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M24 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M25 6 5 VDD VNW pch L=4e-08 W=3.15e-07 
M26 7 11 6 VNW pch L=4e-08 W=2.5e-07 
M27 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M28 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M29 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M30 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M32 VDD 11 10 VNW pch L=4e-08 W=3.45e-07 
M33 11 CK VDD VNW pch L=4e-08 W=2.5e-07 
.ENDS


.SUBCKT SDFFYQ_X3M_A9TR Q VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 21 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 8 7 VSS VPW nch L=4e-08 W=2.5e-07 
M13 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M14 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M15 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M16 VSS 11 10 VPW nch L=4e-08 W=2.4e-07 
M17 11 CK VSS VPW nch L=4e-08 W=2.4e-07 
M18 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M19 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M20 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M21 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M22 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M23 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M24 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M25 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M26 6 5 VDD VNW pch L=4e-08 W=3.8e-07 
M27 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M28 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M29 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M30 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M31 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M33 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD 11 10 VNW pch L=4e-08 W=3.6e-07 
M35 11 CK VDD VNW pch L=4e-08 W=2.6e-07 
.ENDS


.SUBCKT SDFFYQ_X4M_A9TR Q VDD VNW VPW VSS CK D SE SI
M0 3 SE VSS VPW nch L=4e-08 W=1.2e-07 
M1 20 SE 4 VPW nch L=4e-08 W=1.2e-07 
M2 VSS SI 20 VPW nch L=4e-08 W=1.2e-07 
M3 21 3 VSS VPW nch L=4e-08 W=3.1e-07 
M4 4 D 21 VPW nch L=4e-08 W=3.1e-07 
M5 5 11 4 VPW nch L=4e-08 W=3.1e-07 
M6 22 10 5 VPW nch L=4e-08 W=1.2e-07 
M7 VSS 6 22 VPW nch L=4e-08 W=1.2e-07 
M8 6 5 VSS VPW nch L=4e-08 W=3.1e-07 
M9 7 10 6 VPW nch L=4e-08 W=3.1e-07 
M10 23 11 7 VPW nch L=4e-08 W=1.2e-07 
M11 VSS 8 23 VPW nch L=4e-08 W=1.2e-07 
M12 8 7 VSS VPW nch L=4e-08 W=2.5e-07 
M13 VSS 7 8 VPW nch L=4e-08 W=2.5e-07 
M14 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M15 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M16 Q 8 VSS VPW nch L=4e-08 W=3.1e-07 
M17 VSS 8 Q VPW nch L=4e-08 W=3.1e-07 
M18 VSS 11 10 VPW nch L=4e-08 W=2.4e-07 
M19 11 CK VSS VPW nch L=4e-08 W=2.4e-07 
M20 3 SE VDD VNW pch L=4e-08 W=1.7e-07 
M21 16 3 4 VNW pch L=4e-08 W=1.55e-07 
M22 VDD SI 16 VNW pch L=4e-08 W=1.55e-07 
M23 17 SE VDD VNW pch L=4e-08 W=3.8e-07 
M24 4 D 17 VNW pch L=4e-08 W=3.8e-07 
M25 5 10 4 VNW pch L=4e-08 W=3.1e-07 
M26 18 11 5 VNW pch L=4e-08 W=1.2e-07 
M27 VDD 6 18 VNW pch L=4e-08 W=1.2e-07 
M28 6 5 VDD VNW pch L=4e-08 W=3.8e-07 
M29 7 11 6 VNW pch L=4e-08 W=3.1e-07 
M30 19 10 7 VNW pch L=4e-08 W=1.2e-07 
M31 VDD 8 19 VNW pch L=4e-08 W=1.2e-07 
M32 8 7 VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD 7 8 VNW pch L=4e-08 W=3.8e-07 
M34 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M35 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M36 Q 8 VDD VNW pch L=4e-08 W=3.8e-07 
M37 VDD 8 Q VNW pch L=4e-08 W=3.8e-07 
M38 VDD 11 10 VNW pch L=4e-08 W=3.6e-07 
M39 11 CK VDD VNW pch L=4e-08 W=2.6e-07 
.ENDS


.SUBCKT TIEHI_X1M_A9TR Y VDD VNW VPW VSS
M0 3 2 VSS VPW nch L=4e-08 W=1.2e-07 
M1 VSS 3 3 VPW nch L=4e-08 W=1.2e-07 
M2 VDD 3 2 VNW pch L=4e-08 W=1.2e-07 
M3 Y 3 VDD VNW pch L=4e-08 W=4e-07 
.ENDS


.SUBCKT TIELO_X1M_A9TR Y VDD VNW VPW VSS
M0 VSS 4 1 VPW nch L=4e-08 W=1.2e-07 
M1 Y 4 VSS VPW nch L=4e-08 W=4e-07 
M2 4 1 VDD VNW pch L=4e-08 W=1.2e-07 
M3 VDD 4 4 VNW pch L=4e-08 W=1.2e-07 
.ENDS


.SUBCKT XNOR2_X0P5M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y A 4 VPW nch L=4e-08 W=1.2e-07 
M2 6 3 Y VPW nch L=4e-08 W=1.2e-07 
M3 VSS B 6 VPW nch L=4e-08 W=1.2e-07 
M4 4 6 VSS VPW nch L=4e-08 W=1.2e-07 
M5 3 A VDD VNW pch L=4e-08 W=1.9e-07 
M6 Y 3 4 VNW pch L=4e-08 W=1.9e-07 
M7 6 A Y VNW pch L=4e-08 W=1.9e-07 
M8 VDD B 6 VNW pch L=4e-08 W=1.9e-07 
M9 4 6 VDD VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT XNOR2_X0P7M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=1.7e-07 
M1 Y A 4 VPW nch L=4e-08 W=1.7e-07 
M2 6 3 Y VPW nch L=4e-08 W=1.7e-07 
M3 VSS B 6 VPW nch L=4e-08 W=1.7e-07 
M4 4 6 VSS VPW nch L=4e-08 W=1.7e-07 
M5 3 A VDD VNW pch L=4e-08 W=2.35e-07 
M6 Y 3 4 VNW pch L=4e-08 W=2.35e-07 
M7 6 A Y VNW pch L=4e-08 W=2.35e-07 
M8 VDD B 6 VNW pch L=4e-08 W=2.35e-07 
M9 4 6 VDD VNW pch L=4e-08 W=2.35e-07 
.ENDS


.SUBCKT XNOR2_X1M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=2.45e-07 
M1 Y A 4 VPW nch L=4e-08 W=2.45e-07 
M2 5 3 Y VPW nch L=4e-08 W=2.45e-07 
M3 VSS B 5 VPW nch L=4e-08 W=2.45e-07 
M4 4 5 VSS VPW nch L=4e-08 W=2.45e-07 
M5 3 A VDD VNW pch L=4e-08 W=3.8e-07 
M6 Y A 5 VNW pch L=4e-08 W=3.8e-07 
M7 4 3 Y VNW pch L=4e-08 W=3.8e-07 
M8 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M9 4 5 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XNOR2_X1P4M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=1.9e-07 
M1 VSS A 3 VPW nch L=4e-08 W=1.9e-07 
M2 Y A 4 VPW nch L=4e-08 W=3.8e-07 
M3 5 3 Y VPW nch L=4e-08 W=3.8e-07 
M4 VSS B 5 VPW nch L=4e-08 W=3.8e-07 
M5 4 5 VSS VPW nch L=4e-08 W=1.9e-07 
M6 VSS 5 4 VPW nch L=4e-08 W=1.9e-07 
M7 3 A VDD VNW pch L=4e-08 W=3.3e-07 
M8 VDD A 3 VNW pch L=4e-08 W=3.3e-07 
M9 Y A 5 VNW pch L=4e-08 W=4e-07 
M10 4 3 Y VNW pch L=4e-08 W=4e-07 
M11 5 B VDD VNW pch L=4e-08 W=3.3e-07 
M12 VDD B 5 VNW pch L=4e-08 W=3.3e-07 
M13 4 5 VDD VNW pch L=4e-08 W=3.3e-07 
M14 VDD 5 4 VNW pch L=4e-08 W=3.3e-07 
.ENDS


.SUBCKT XNOR2_X2M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS A 3 VPW nch L=4e-08 W=2.45e-07 
M2 5 A Y VPW nch L=4e-08 W=2.45e-07 
M3 Y A 5 VPW nch L=4e-08 W=2.45e-07 
M4 6 3 Y VPW nch L=4e-08 W=2.45e-07 
M5 Y 3 6 VPW nch L=4e-08 W=2.45e-07 
M6 VSS B 6 VPW nch L=4e-08 W=3.7e-07 
M7 5 6 VSS VPW nch L=4e-08 W=2.45e-07 
M8 VSS 6 5 VPW nch L=4e-08 W=2.45e-07 
M9 3 A VDD VNW pch L=4e-08 W=3.8e-07 
M10 VDD A 3 VNW pch L=4e-08 W=3.8e-07 
M11 6 A Y VNW pch L=4e-08 W=3.8e-07 
M12 Y A 6 VNW pch L=4e-08 W=3.8e-07 
M13 5 3 Y VNW pch L=4e-08 W=3.8e-07 
M14 Y 3 5 VNW pch L=4e-08 W=3.8e-07 
M15 6 B VDD VNW pch L=4e-08 W=3.8e-07 
M16 VDD B 6 VNW pch L=4e-08 W=3.8e-07 
M17 5 6 VDD VNW pch L=4e-08 W=3.8e-07 
M18 VDD 6 5 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XNOR2_X3M_A9TR Y VDD VNW VPW VSS A B
M0 VSS A 1 VPW nch L=4e-08 W=2.45e-07 
M1 1 A VSS VPW nch L=4e-08 W=2.45e-07 
M2 VSS A 1 VPW nch L=4e-08 W=2.45e-07 
M3 Y A 4 VPW nch L=4e-08 W=2.45e-07 
M4 4 A Y VPW nch L=4e-08 W=2.45e-07 
M5 Y A 4 VPW nch L=4e-08 W=2.45e-07 
M6 5 1 Y VPW nch L=4e-08 W=2.45e-07 
M7 Y 1 5 VPW nch L=4e-08 W=2.45e-07 
M8 5 1 Y VPW nch L=4e-08 W=2.45e-07 
M9 VSS B 5 VPW nch L=4e-08 W=2.45e-07 
M10 5 B VSS VPW nch L=4e-08 W=2.45e-07 
M11 VSS B 5 VPW nch L=4e-08 W=2.45e-07 
M12 4 5 VSS VPW nch L=4e-08 W=2.45e-07 
M13 VSS 5 4 VPW nch L=4e-08 W=2.45e-07 
M14 4 5 VSS VPW nch L=4e-08 W=2.45e-07 
M15 VDD A 1 VNW pch L=4e-08 W=3.8e-07 
M16 1 A VDD VNW pch L=4e-08 W=3.8e-07 
M17 VDD A 1 VNW pch L=4e-08 W=3.8e-07 
M18 Y A 5 VNW pch L=4e-08 W=3.8e-07 
M19 5 A Y VNW pch L=4e-08 W=3.8e-07 
M20 Y A 5 VNW pch L=4e-08 W=3.8e-07 
M21 4 1 Y VNW pch L=4e-08 W=3.8e-07 
M22 Y 1 4 VNW pch L=4e-08 W=3.8e-07 
M23 4 1 Y VNW pch L=4e-08 W=3.8e-07 
M24 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M25 5 B VDD VNW pch L=4e-08 W=3.8e-07 
M26 VDD B 5 VNW pch L=4e-08 W=3.8e-07 
M27 4 5 VDD VNW pch L=4e-08 W=3.8e-07 
M28 VDD 5 4 VNW pch L=4e-08 W=3.8e-07 
M29 4 5 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XNOR2_X4M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS A 3 VPW nch L=4e-08 W=2.45e-07 
M2 3 A VSS VPW nch L=4e-08 W=2.45e-07 
M3 VSS A 3 VPW nch L=4e-08 W=2.45e-07 
M4 5 A Y VPW nch L=4e-08 W=2.45e-07 
M5 Y A 5 VPW nch L=4e-08 W=2.45e-07 
M6 5 A Y VPW nch L=4e-08 W=2.45e-07 
M7 Y A 5 VPW nch L=4e-08 W=2.45e-07 
M8 6 3 Y VPW nch L=4e-08 W=2.45e-07 
M9 Y 3 6 VPW nch L=4e-08 W=2.45e-07 
M10 6 3 Y VPW nch L=4e-08 W=2.45e-07 
M11 Y 3 6 VPW nch L=4e-08 W=2.45e-07 
M12 VSS B 6 VPW nch L=4e-08 W=3.3e-07 
M13 6 B VSS VPW nch L=4e-08 W=3.3e-07 
M14 VSS B 6 VPW nch L=4e-08 W=3.3e-07 
M15 5 6 VSS VPW nch L=4e-08 W=2.45e-07 
M16 VSS 6 5 VPW nch L=4e-08 W=2.45e-07 
M17 5 6 VSS VPW nch L=4e-08 W=2.45e-07 
M18 VSS 6 5 VPW nch L=4e-08 W=2.45e-07 
M19 3 A VDD VNW pch L=4e-08 W=3.8e-07 
M20 VDD A 3 VNW pch L=4e-08 W=3.8e-07 
M21 3 A VDD VNW pch L=4e-08 W=3.8e-07 
M22 VDD A 3 VNW pch L=4e-08 W=3.8e-07 
M23 6 A Y VNW pch L=4e-08 W=3.8e-07 
M24 Y A 6 VNW pch L=4e-08 W=3.8e-07 
M25 6 A Y VNW pch L=4e-08 W=3.8e-07 
M26 Y A 6 VNW pch L=4e-08 W=3.8e-07 
M27 5 3 Y VNW pch L=4e-08 W=3.8e-07 
M28 Y 3 5 VNW pch L=4e-08 W=3.8e-07 
M29 5 3 Y VNW pch L=4e-08 W=3.8e-07 
M30 Y 3 5 VNW pch L=4e-08 W=3.8e-07 
M31 6 B VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD B 6 VNW pch L=4e-08 W=3.8e-07 
M33 6 B VDD VNW pch L=4e-08 W=3.8e-07 
M34 VDD B 6 VNW pch L=4e-08 W=3.8e-07 
M35 5 6 VDD VNW pch L=4e-08 W=3.8e-07 
M36 VDD 6 5 VNW pch L=4e-08 W=3.8e-07 
M37 5 6 VDD VNW pch L=4e-08 W=3.8e-07 
M38 VDD 6 5 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XNOR3_X0P5M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 B VSS VPW nch L=4e-08 W=1.2e-07 
M2 6 B 1 VPW nch L=4e-08 W=1.2e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 1 5 VPW nch L=4e-08 W=1.2e-07 
M5 7 6 VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 9 6 VPW nch L=4e-08 W=1.2e-07 
M7 7 A 8 VPW nch L=4e-08 W=1.2e-07 
M8 VSS A 9 VPW nch L=4e-08 W=1.2e-07 
M9 Y 8 VSS VPW nch L=4e-08 W=1.55e-07 
M10 VDD C 1 VNW pch L=4e-08 W=1.9e-07 
M11 4 B VDD VNW pch L=4e-08 W=1.9e-07 
M12 6 B 5 VNW pch L=4e-08 W=1.9e-07 
M13 1 4 6 VNW pch L=4e-08 W=1.9e-07 
M14 VDD 1 5 VNW pch L=4e-08 W=1.9e-07 
M15 7 6 VDD VNW pch L=4e-08 W=1.9e-07 
M16 8 9 7 VNW pch L=4e-08 W=1.9e-07 
M17 6 A 8 VNW pch L=4e-08 W=1.9e-07 
M18 VDD A 9 VNW pch L=4e-08 W=1.9e-07 
M19 Y 8 VDD VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT XNOR3_X0P7M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=1.7e-07 
M1 4 B VSS VPW nch L=4e-08 W=1.7e-07 
M2 6 B 1 VPW nch L=4e-08 W=1.7e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.7e-07 
M4 VSS 1 5 VPW nch L=4e-08 W=1.7e-07 
M5 7 6 VSS VPW nch L=4e-08 W=1.7e-07 
M6 8 9 6 VPW nch L=4e-08 W=1.7e-07 
M7 7 A 8 VPW nch L=4e-08 W=1.7e-07 
M8 VSS A 9 VPW nch L=4e-08 W=1.7e-07 
M9 Y 8 VSS VPW nch L=4e-08 W=2.15e-07 
M10 VDD C 1 VNW pch L=4e-08 W=2.65e-07 
M11 4 B VDD VNW pch L=4e-08 W=2.65e-07 
M12 6 B 5 VNW pch L=4e-08 W=2.65e-07 
M13 1 4 6 VNW pch L=4e-08 W=2.65e-07 
M14 VDD 1 5 VNW pch L=4e-08 W=2.65e-07 
M15 7 6 VDD VNW pch L=4e-08 W=2.65e-07 
M16 8 9 7 VNW pch L=4e-08 W=2.65e-07 
M17 6 A 8 VNW pch L=4e-08 W=2.65e-07 
M18 VDD A 9 VNW pch L=4e-08 W=2.65e-07 
M19 Y 8 VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT XNOR3_X1M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=2.45e-07 
M1 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M2 6 B 1 VPW nch L=4e-08 W=2.45e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M4 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M5 7 6 VSS VPW nch L=4e-08 W=2.45e-07 
M6 8 9 6 VPW nch L=4e-08 W=2.45e-07 
M7 7 A 8 VPW nch L=4e-08 W=2.45e-07 
M8 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M9 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M11 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M12 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M13 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M14 VDD 1 5 VNW pch L=4e-08 W=3.8e-07 
M15 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M16 8 9 7 VNW pch L=4e-08 W=3.8e-07 
M17 6 A 8 VNW pch L=4e-08 W=3.8e-07 
M18 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M19 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XNOR3_X1P4M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=2.45e-07 
M1 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M2 6 B 1 VPW nch L=4e-08 W=2.45e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M4 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M5 7 6 VSS VPW nch L=4e-08 W=2.45e-07 
M6 8 9 6 VPW nch L=4e-08 W=2.45e-07 
M7 7 A 8 VPW nch L=4e-08 W=2.45e-07 
M8 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M9 Y 8 VSS VPW nch L=4e-08 W=2.3e-07 
M10 VSS 8 Y VPW nch L=4e-08 W=2.3e-07 
M11 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M12 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M13 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M14 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M15 VDD 1 5 VNW pch L=4e-08 W=3.8e-07 
M16 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M17 8 9 7 VNW pch L=4e-08 W=3.8e-07 
M18 6 A 8 VNW pch L=4e-08 W=3.8e-07 
M19 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M20 Y 8 VDD VNW pch L=4e-08 W=2.8e-07 
M21 VDD 8 Y VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT XNOR3_X2M_A9TR Y VDD VNW VPW VSS A B C
M0 3 C VSS VPW nch L=4e-08 W=1.75e-07 
M1 VSS C 3 VPW nch L=4e-08 W=1.75e-07 
M2 4 B VSS VPW nch L=4e-08 W=3.5e-07 
M3 6 B 3 VPW nch L=4e-08 W=3.5e-07 
M4 5 4 6 VPW nch L=4e-08 W=3.5e-07 
M5 VSS 3 5 VPW nch L=4e-08 W=1.75e-07 
M6 5 3 VSS VPW nch L=4e-08 W=1.75e-07 
M7 7 6 VSS VPW nch L=4e-08 W=1.75e-07 
M8 VSS 6 7 VPW nch L=4e-08 W=1.75e-07 
M9 8 9 6 VPW nch L=4e-08 W=3.5e-07 
M10 7 A 8 VPW nch L=4e-08 W=3.5e-07 
M11 VSS A 9 VPW nch L=4e-08 W=3.5e-07 
M12 Y 8 VSS VPW nch L=4e-08 W=3.5e-07 
M13 VSS 8 Y VPW nch L=4e-08 W=3.5e-07 
M14 3 C VDD VNW pch L=4e-08 W=3e-07 
M15 VDD C 3 VNW pch L=4e-08 W=3e-07 
M16 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M17 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M18 3 4 6 VNW pch L=4e-08 W=3.8e-07 
M19 VDD 3 5 VNW pch L=4e-08 W=3e-07 
M20 5 3 VDD VNW pch L=4e-08 W=3e-07 
M21 7 6 VDD VNW pch L=4e-08 W=3e-07 
M22 VDD 6 7 VNW pch L=4e-08 W=3e-07 
M23 8 9 7 VNW pch L=4e-08 W=3.8e-07 
M24 6 A 8 VNW pch L=4e-08 W=3.8e-07 
M25 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M26 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XNOR3_X3M_A9TR Y VDD VNW VPW VSS A B C
M0 3 C VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS C 3 VPW nch L=4e-08 W=2.45e-07 
M2 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M3 VSS B 4 VPW nch L=4e-08 W=2.45e-07 
M4 3 B 5 VPW nch L=4e-08 W=2.45e-07 
M5 5 B 3 VPW nch L=4e-08 W=2.45e-07 
M6 6 4 5 VPW nch L=4e-08 W=2.45e-07 
M7 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M8 VSS 3 6 VPW nch L=4e-08 W=2.45e-07 
M9 6 3 VSS VPW nch L=4e-08 W=2.45e-07 
M10 7 5 VSS VPW nch L=4e-08 W=2.45e-07 
M11 VSS 5 7 VPW nch L=4e-08 W=2.45e-07 
M12 5 9 8 VPW nch L=4e-08 W=2.45e-07 
M13 8 9 5 VPW nch L=4e-08 W=2.45e-07 
M14 7 A 8 VPW nch L=4e-08 W=2.45e-07 
M15 8 A 7 VPW nch L=4e-08 W=2.45e-07 
M16 9 A VSS VPW nch L=4e-08 W=2.45e-07 
M17 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M18 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 8 Y VPW nch L=4e-08 W=3.1e-07 
M20 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M21 3 C VDD VNW pch L=4e-08 W=3.8e-07 
M22 VDD C 3 VNW pch L=4e-08 W=3.8e-07 
M23 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M24 VDD B 4 VNW pch L=4e-08 W=3.8e-07 
M25 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M26 5 B 6 VNW pch L=4e-08 W=3.8e-07 
M27 3 4 5 VNW pch L=4e-08 W=3.8e-07 
M28 5 4 3 VNW pch L=4e-08 W=3.8e-07 
M29 6 3 VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD 3 6 VNW pch L=4e-08 W=3.8e-07 
M31 7 5 VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD 5 7 VNW pch L=4e-08 W=3.8e-07 
M33 7 9 8 VNW pch L=4e-08 W=3.8e-07 
M34 8 9 7 VNW pch L=4e-08 W=3.8e-07 
M35 5 A 8 VNW pch L=4e-08 W=3.8e-07 
M36 8 A 5 VNW pch L=4e-08 W=3.8e-07 
M37 9 A VDD VNW pch L=4e-08 W=3.8e-07 
M38 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M39 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
M41 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XNOR3_X4M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=2.45e-07 
M1 1 C VSS VPW nch L=4e-08 W=2.45e-07 
M2 VSS C 1 VPW nch L=4e-08 W=2.45e-07 
M3 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M4 VSS B 4 VPW nch L=4e-08 W=2.45e-07 
M5 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M6 6 B 1 VPW nch L=4e-08 W=2.45e-07 
M7 1 B 6 VPW nch L=4e-08 W=2.45e-07 
M8 6 B 1 VPW nch L=4e-08 W=2.45e-07 
M9 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M10 6 4 5 VPW nch L=4e-08 W=2.45e-07 
M11 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M12 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M13 5 1 VSS VPW nch L=4e-08 W=2.45e-07 
M14 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M15 7 6 VSS VPW nch L=4e-08 W=2.45e-07 
M16 VSS 6 7 VPW nch L=4e-08 W=2.45e-07 
M17 7 6 VSS VPW nch L=4e-08 W=2.45e-07 
M18 6 9 8 VPW nch L=4e-08 W=3.65e-07 
M19 8 9 6 VPW nch L=4e-08 W=3.65e-07 
M20 7 A 8 VPW nch L=4e-08 W=3.65e-07 
M21 8 A 7 VPW nch L=4e-08 W=3.65e-07 
M22 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M23 9 A VSS VPW nch L=4e-08 W=2.45e-07 
M24 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M25 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M26 VSS 8 Y VPW nch L=4e-08 W=3.1e-07 
M27 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M28 VSS 8 Y VPW nch L=4e-08 W=3.1e-07 
M29 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M30 1 C VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M32 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M33 VDD B 4 VNW pch L=4e-08 W=3.8e-07 
M34 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M35 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M36 5 B 6 VNW pch L=4e-08 W=3.8e-07 
M37 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M38 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M39 6 4 1 VNW pch L=4e-08 W=3.8e-07 
M40 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M41 5 1 VDD VNW pch L=4e-08 W=3.8e-07 
M42 VDD 1 5 VNW pch L=4e-08 W=3.8e-07 
M43 5 1 VDD VNW pch L=4e-08 W=3.8e-07 
M44 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M45 VDD 6 7 VNW pch L=4e-08 W=3.8e-07 
M46 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M47 8 9 7 VNW pch L=4e-08 W=3.8e-07 
M48 7 9 8 VNW pch L=4e-08 W=3.8e-07 
M49 8 9 7 VNW pch L=4e-08 W=3.8e-07 
M50 6 A 8 VNW pch L=4e-08 W=3.8e-07 
M51 8 A 6 VNW pch L=4e-08 W=3.8e-07 
M52 6 A 8 VNW pch L=4e-08 W=3.8e-07 
M53 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M54 9 A VDD VNW pch L=4e-08 W=3.8e-07 
M55 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M56 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M57 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
M58 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M59 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XOR2_X0P5M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=1.2e-07 
M1 Y 3 4 VPW nch L=4e-08 W=1.2e-07 
M2 6 A Y VPW nch L=4e-08 W=1.2e-07 
M3 VSS B 6 VPW nch L=4e-08 W=1.2e-07 
M4 4 6 VSS VPW nch L=4e-08 W=1.2e-07 
M5 3 A VDD VNW pch L=4e-08 W=1.9e-07 
M6 Y A 4 VNW pch L=4e-08 W=1.9e-07 
M7 6 3 Y VNW pch L=4e-08 W=1.9e-07 
M8 VDD B 6 VNW pch L=4e-08 W=1.9e-07 
M9 4 6 VDD VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT XOR2_X0P7M_A9TR Y VDD VNW VPW VSS A B
M0 3 A VSS VPW nch L=4e-08 W=1.7e-07 
M1 Y 3 4 VPW nch L=4e-08 W=1.7e-07 
M2 6 A Y VPW nch L=4e-08 W=1.7e-07 
M3 VSS B 6 VPW nch L=4e-08 W=1.7e-07 
M4 4 6 VSS VPW nch L=4e-08 W=1.7e-07 
M5 3 A VDD VNW pch L=4e-08 W=2.35e-07 
M6 Y A 4 VNW pch L=4e-08 W=2.35e-07 
M7 6 3 Y VNW pch L=4e-08 W=2.35e-07 
M8 VDD B 6 VNW pch L=4e-08 W=2.35e-07 
M9 4 6 VDD VNW pch L=4e-08 W=2.35e-07 
.ENDS


.SUBCKT XOR2_X1M_A9TR Y VDD VNW VPW VSS A B
M0 VSS B 1 VPW nch L=4e-08 W=2.45e-07 
M1 4 A VSS VPW nch L=4e-08 W=2.45e-07 
M2 Y A 1 VPW nch L=4e-08 W=2.45e-07 
M3 5 4 Y VPW nch L=4e-08 W=2.45e-07 
M4 5 1 VSS VPW nch L=4e-08 W=2.45e-07 
M5 VDD B 1 VNW pch L=4e-08 W=3.8e-07 
M6 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M7 Y A 5 VNW pch L=4e-08 W=3.8e-07 
M8 1 4 Y VNW pch L=4e-08 W=3.8e-07 
M9 5 1 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XOR2_X1P4M_A9TR Y VDD VNW VPW VSS A B
M0 3 B VSS VPW nch L=4e-08 W=1.9e-07 
M1 VSS B 3 VPW nch L=4e-08 W=1.9e-07 
M2 4 A VSS VPW nch L=4e-08 W=1.9e-07 
M3 VSS A 4 VPW nch L=4e-08 W=1.9e-07 
M4 Y A 3 VPW nch L=4e-08 W=3.8e-07 
M5 5 4 Y VPW nch L=4e-08 W=3.8e-07 
M6 5 3 VSS VPW nch L=4e-08 W=1.9e-07 
M7 VSS 3 5 VPW nch L=4e-08 W=1.9e-07 
M8 3 B VDD VNW pch L=4e-08 W=3.3e-07 
M9 VDD B 3 VNW pch L=4e-08 W=3.3e-07 
M10 4 A VDD VNW pch L=4e-08 W=3.3e-07 
M11 VDD A 4 VNW pch L=4e-08 W=3.3e-07 
M12 Y A 5 VNW pch L=4e-08 W=4e-07 
M13 3 4 Y VNW pch L=4e-08 W=4e-07 
M14 5 3 VDD VNW pch L=4e-08 W=3.3e-07 
M15 VDD 3 5 VNW pch L=4e-08 W=3.3e-07 
.ENDS


.SUBCKT XOR2_X2M_A9TR Y VDD VNW VPW VSS A B
M0 3 B VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.45e-07 
M2 4 A VSS VPW nch L=4e-08 W=2.45e-07 
M3 VSS A 4 VPW nch L=4e-08 W=2.45e-07 
M4 3 A Y VPW nch L=4e-08 W=2.45e-07 
M5 Y A 3 VPW nch L=4e-08 W=2.45e-07 
M6 6 4 Y VPW nch L=4e-08 W=2.45e-07 
M7 Y 4 6 VPW nch L=4e-08 W=2.45e-07 
M8 6 3 VSS VPW nch L=4e-08 W=2.45e-07 
M9 VSS 3 6 VPW nch L=4e-08 W=2.45e-07 
M10 3 B VDD VNW pch L=4e-08 W=3.8e-07 
M11 VDD B 3 VNW pch L=4e-08 W=3.8e-07 
M12 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M13 VDD A 4 VNW pch L=4e-08 W=3.8e-07 
M14 6 A Y VNW pch L=4e-08 W=3.8e-07 
M15 Y A 6 VNW pch L=4e-08 W=3.8e-07 
M16 3 4 Y VNW pch L=4e-08 W=3.8e-07 
M17 Y 4 3 VNW pch L=4e-08 W=3.8e-07 
M18 6 3 VDD VNW pch L=4e-08 W=3.8e-07 
M19 VDD 3 6 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XOR2_X3M_A9TR Y VDD VNW VPW VSS A B
M0 VSS B 1 VPW nch L=4e-08 W=2.45e-07 
M1 1 B VSS VPW nch L=4e-08 W=2.45e-07 
M2 VSS B 1 VPW nch L=4e-08 W=2.45e-07 
M3 4 A VSS VPW nch L=4e-08 W=2.45e-07 
M4 VSS A 4 VPW nch L=4e-08 W=2.45e-07 
M5 4 A VSS VPW nch L=4e-08 W=2.45e-07 
M6 Y A 1 VPW nch L=4e-08 W=2.45e-07 
M7 1 A Y VPW nch L=4e-08 W=2.45e-07 
M8 Y A 1 VPW nch L=4e-08 W=2.45e-07 
M9 5 4 Y VPW nch L=4e-08 W=2.45e-07 
M10 Y 4 5 VPW nch L=4e-08 W=2.45e-07 
M11 5 4 Y VPW nch L=4e-08 W=2.45e-07 
M12 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M13 5 1 VSS VPW nch L=4e-08 W=2.45e-07 
M14 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M15 VDD B 1 VNW pch L=4e-08 W=3.8e-07 
M16 1 B VDD VNW pch L=4e-08 W=3.8e-07 
M17 VDD B 1 VNW pch L=4e-08 W=3.8e-07 
M18 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M19 VDD A 4 VNW pch L=4e-08 W=3.8e-07 
M20 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M21 Y A 5 VNW pch L=4e-08 W=3.8e-07 
M22 5 A Y VNW pch L=4e-08 W=3.8e-07 
M23 Y A 5 VNW pch L=4e-08 W=3.8e-07 
M24 1 4 Y VNW pch L=4e-08 W=3.8e-07 
M25 Y 4 1 VNW pch L=4e-08 W=3.8e-07 
M26 1 4 Y VNW pch L=4e-08 W=3.8e-07 
M27 5 1 VDD VNW pch L=4e-08 W=3.8e-07 
M28 VDD 1 5 VNW pch L=4e-08 W=3.8e-07 
M29 5 1 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XOR2_X4M_A9TR Y VDD VNW VPW VSS A B
M0 3 B VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS B 3 VPW nch L=4e-08 W=2.45e-07 
M2 3 B VSS VPW nch L=4e-08 W=2.45e-07 
M3 VSS B 3 VPW nch L=4e-08 W=2.45e-07 
M4 4 A VSS VPW nch L=4e-08 W=2.45e-07 
M5 VSS A 4 VPW nch L=4e-08 W=2.45e-07 
M6 4 A VSS VPW nch L=4e-08 W=2.45e-07 
M7 VSS A 4 VPW nch L=4e-08 W=2.45e-07 
M8 3 A Y VPW nch L=4e-08 W=2.45e-07 
M9 Y A 3 VPW nch L=4e-08 W=2.45e-07 
M10 3 A Y VPW nch L=4e-08 W=2.45e-07 
M11 Y A 3 VPW nch L=4e-08 W=2.45e-07 
M12 6 4 Y VPW nch L=4e-08 W=2.45e-07 
M13 Y 4 6 VPW nch L=4e-08 W=2.45e-07 
M14 6 4 Y VPW nch L=4e-08 W=2.45e-07 
M15 Y 4 6 VPW nch L=4e-08 W=2.45e-07 
M16 6 3 VSS VPW nch L=4e-08 W=2.45e-07 
M17 VSS 3 6 VPW nch L=4e-08 W=2.45e-07 
M18 6 3 VSS VPW nch L=4e-08 W=2.45e-07 
M19 VSS 3 6 VPW nch L=4e-08 W=2.45e-07 
M20 3 B VDD VNW pch L=4e-08 W=3.8e-07 
M21 VDD B 3 VNW pch L=4e-08 W=3.8e-07 
M22 3 B VDD VNW pch L=4e-08 W=3.8e-07 
M23 VDD B 3 VNW pch L=4e-08 W=3.8e-07 
M24 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M25 VDD A 4 VNW pch L=4e-08 W=3.8e-07 
M26 4 A VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD A 4 VNW pch L=4e-08 W=3.8e-07 
M28 6 A Y VNW pch L=4e-08 W=3.8e-07 
M29 Y A 6 VNW pch L=4e-08 W=3.8e-07 
M30 6 A Y VNW pch L=4e-08 W=3.8e-07 
M31 Y A 6 VNW pch L=4e-08 W=3.8e-07 
M32 3 4 Y VNW pch L=4e-08 W=3.8e-07 
M33 Y 4 3 VNW pch L=4e-08 W=3.8e-07 
M34 3 4 Y VNW pch L=4e-08 W=3.8e-07 
M35 Y 4 3 VNW pch L=4e-08 W=3.8e-07 
M36 6 3 VDD VNW pch L=4e-08 W=3.8e-07 
M37 VDD 3 6 VNW pch L=4e-08 W=3.8e-07 
M38 6 3 VDD VNW pch L=4e-08 W=3.8e-07 
M39 VDD 3 6 VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XOR3_X0P5M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=1.2e-07 
M1 4 B VSS VPW nch L=4e-08 W=1.2e-07 
M2 6 B 1 VPW nch L=4e-08 W=1.2e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.2e-07 
M4 VSS 1 5 VPW nch L=4e-08 W=1.2e-07 
M5 7 6 VSS VPW nch L=4e-08 W=1.2e-07 
M6 8 9 7 VPW nch L=4e-08 W=1.2e-07 
M7 8 A 6 VPW nch L=4e-08 W=1.2e-07 
M8 VSS A 9 VPW nch L=4e-08 W=1.2e-07 
M9 Y 8 VSS VPW nch L=4e-08 W=1.55e-07 
M10 VDD C 1 VNW pch L=4e-08 W=1.9e-07 
M11 4 B VDD VNW pch L=4e-08 W=1.9e-07 
M12 6 B 5 VNW pch L=4e-08 W=1.9e-07 
M13 1 4 6 VNW pch L=4e-08 W=1.9e-07 
M14 VDD 1 5 VNW pch L=4e-08 W=1.9e-07 
M15 7 6 VDD VNW pch L=4e-08 W=1.9e-07 
M16 8 9 6 VNW pch L=4e-08 W=1.9e-07 
M17 7 A 8 VNW pch L=4e-08 W=1.9e-07 
M18 VDD A 9 VNW pch L=4e-08 W=1.9e-07 
M19 Y 8 VDD VNW pch L=4e-08 W=1.9e-07 
.ENDS


.SUBCKT XOR3_X0P7M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=1.7e-07 
M1 4 B VSS VPW nch L=4e-08 W=1.7e-07 
M2 6 B 1 VPW nch L=4e-08 W=1.7e-07 
M3 5 4 6 VPW nch L=4e-08 W=1.7e-07 
M4 VSS 1 5 VPW nch L=4e-08 W=1.7e-07 
M5 7 6 VSS VPW nch L=4e-08 W=1.7e-07 
M6 8 9 7 VPW nch L=4e-08 W=1.7e-07 
M7 6 A 8 VPW nch L=4e-08 W=1.7e-07 
M8 VSS A 9 VPW nch L=4e-08 W=1.7e-07 
M9 Y 8 VSS VPW nch L=4e-08 W=2.15e-07 
M10 VDD C 1 VNW pch L=4e-08 W=2.65e-07 
M11 4 B VDD VNW pch L=4e-08 W=2.65e-07 
M12 6 B 5 VNW pch L=4e-08 W=2.65e-07 
M13 1 4 6 VNW pch L=4e-08 W=2.65e-07 
M14 VDD 1 5 VNW pch L=4e-08 W=2.65e-07 
M15 7 6 VDD VNW pch L=4e-08 W=2.65e-07 
M16 8 9 6 VNW pch L=4e-08 W=2.65e-07 
M17 7 A 8 VNW pch L=4e-08 W=2.65e-07 
M18 VDD A 9 VNW pch L=4e-08 W=2.65e-07 
M19 Y 8 VDD VNW pch L=4e-08 W=2.65e-07 
.ENDS


.SUBCKT XOR3_X1M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=2.45e-07 
M1 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M2 6 B 1 VPW nch L=4e-08 W=2.45e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M4 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M5 7 6 VSS VPW nch L=4e-08 W=2.45e-07 
M6 8 9 7 VPW nch L=4e-08 W=2.45e-07 
M7 6 A 8 VPW nch L=4e-08 W=2.45e-07 
M8 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M9 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M10 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M11 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M12 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M13 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M14 VDD 1 5 VNW pch L=4e-08 W=3.8e-07 
M15 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M16 8 9 6 VNW pch L=4e-08 W=3.8e-07 
M17 7 A 8 VNW pch L=4e-08 W=3.8e-07 
M18 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M19 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XOR3_X1P4M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=2.45e-07 
M1 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M2 6 B 1 VPW nch L=4e-08 W=2.45e-07 
M3 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M4 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M5 7 6 VSS VPW nch L=4e-08 W=2.45e-07 
M6 8 9 7 VPW nch L=4e-08 W=2.45e-07 
M7 6 A 8 VPW nch L=4e-08 W=2.45e-07 
M8 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M9 Y 8 VSS VPW nch L=4e-08 W=2.3e-07 
M10 VSS 8 Y VPW nch L=4e-08 W=2.3e-07 
M11 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M12 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M13 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M14 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M15 VDD 1 5 VNW pch L=4e-08 W=3.8e-07 
M16 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M17 8 9 6 VNW pch L=4e-08 W=3.8e-07 
M18 7 A 8 VNW pch L=4e-08 W=3.8e-07 
M19 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M20 Y 8 VDD VNW pch L=4e-08 W=2.8e-07 
M21 VDD 8 Y VNW pch L=4e-08 W=2.8e-07 
.ENDS


.SUBCKT XOR3_X2M_A9TR Y VDD VNW VPW VSS A B C
M0 3 C VSS VPW nch L=4e-08 W=1.75e-07 
M1 VSS C 3 VPW nch L=4e-08 W=1.75e-07 
M2 4 B VSS VPW nch L=4e-08 W=3.5e-07 
M3 6 B 3 VPW nch L=4e-08 W=3.5e-07 
M4 5 4 6 VPW nch L=4e-08 W=3.5e-07 
M5 VSS 3 5 VPW nch L=4e-08 W=1.75e-07 
M6 5 3 VSS VPW nch L=4e-08 W=1.75e-07 
M7 7 6 VSS VPW nch L=4e-08 W=1.75e-07 
M8 VSS 6 7 VPW nch L=4e-08 W=1.75e-07 
M9 8 9 7 VPW nch L=4e-08 W=3.5e-07 
M10 6 A 8 VPW nch L=4e-08 W=3.5e-07 
M11 VSS A 9 VPW nch L=4e-08 W=3.5e-07 
M12 Y 8 VSS VPW nch L=4e-08 W=3.5e-07 
M13 VSS 8 Y VPW nch L=4e-08 W=3.5e-07 
M14 3 C VDD VNW pch L=4e-08 W=3e-07 
M15 VDD C 3 VNW pch L=4e-08 W=3e-07 
M16 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M17 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M18 3 4 6 VNW pch L=4e-08 W=3.8e-07 
M19 VDD 3 5 VNW pch L=4e-08 W=3e-07 
M20 5 3 VDD VNW pch L=4e-08 W=3e-07 
M21 7 6 VDD VNW pch L=4e-08 W=3e-07 
M22 VDD 6 7 VNW pch L=4e-08 W=3e-07 
M23 8 9 6 VNW pch L=4e-08 W=3.8e-07 
M24 7 A 8 VNW pch L=4e-08 W=3.8e-07 
M25 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M26 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M27 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XOR3_X3M_A9TR Y VDD VNW VPW VSS A B C
M0 3 C VSS VPW nch L=4e-08 W=2.45e-07 
M1 VSS C 3 VPW nch L=4e-08 W=2.45e-07 
M2 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M3 VSS B 4 VPW nch L=4e-08 W=2.45e-07 
M4 3 B 5 VPW nch L=4e-08 W=2.45e-07 
M5 5 B 3 VPW nch L=4e-08 W=2.45e-07 
M6 6 4 5 VPW nch L=4e-08 W=2.45e-07 
M7 5 4 6 VPW nch L=4e-08 W=2.45e-07 
M8 VSS 3 6 VPW nch L=4e-08 W=2.45e-07 
M9 6 3 VSS VPW nch L=4e-08 W=2.45e-07 
M10 7 5 VSS VPW nch L=4e-08 W=2.45e-07 
M11 VSS 5 7 VPW nch L=4e-08 W=2.45e-07 
M12 5 A 8 VPW nch L=4e-08 W=2.45e-07 
M13 8 A 5 VPW nch L=4e-08 W=2.45e-07 
M14 7 9 8 VPW nch L=4e-08 W=2.45e-07 
M15 8 9 7 VPW nch L=4e-08 W=2.45e-07 
M16 9 A VSS VPW nch L=4e-08 W=2.45e-07 
M17 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M18 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M19 VSS 8 Y VPW nch L=4e-08 W=3.1e-07 
M20 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M21 3 C VDD VNW pch L=4e-08 W=3.8e-07 
M22 VDD C 3 VNW pch L=4e-08 W=3.8e-07 
M23 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M24 VDD B 4 VNW pch L=4e-08 W=3.8e-07 
M25 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M26 5 B 6 VNW pch L=4e-08 W=3.8e-07 
M27 3 4 5 VNW pch L=4e-08 W=3.8e-07 
M28 5 4 3 VNW pch L=4e-08 W=3.8e-07 
M29 6 3 VDD VNW pch L=4e-08 W=3.8e-07 
M30 VDD 3 6 VNW pch L=4e-08 W=3.8e-07 
M31 7 5 VDD VNW pch L=4e-08 W=3.8e-07 
M32 VDD 5 7 VNW pch L=4e-08 W=3.8e-07 
M33 7 A 8 VNW pch L=4e-08 W=3.8e-07 
M34 8 A 7 VNW pch L=4e-08 W=3.8e-07 
M35 5 9 8 VNW pch L=4e-08 W=3.8e-07 
M36 8 9 5 VNW pch L=4e-08 W=3.8e-07 
M37 9 A VDD VNW pch L=4e-08 W=3.8e-07 
M38 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M39 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
M41 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
.ENDS


.SUBCKT XOR3_X4M_A9TR Y VDD VNW VPW VSS A B C
M0 VSS C 1 VPW nch L=4e-08 W=2.45e-07 
M1 1 C VSS VPW nch L=4e-08 W=2.45e-07 
M2 VSS C 1 VPW nch L=4e-08 W=2.45e-07 
M3 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M4 VSS B 4 VPW nch L=4e-08 W=2.45e-07 
M5 4 B VSS VPW nch L=4e-08 W=2.45e-07 
M6 1 B 6 VPW nch L=4e-08 W=3.7e-07 
M7 6 B 1 VPW nch L=4e-08 W=3.7e-07 
M8 5 4 6 VPW nch L=4e-08 W=3.7e-07 
M9 6 4 5 VPW nch L=4e-08 W=3.7e-07 
M10 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M11 5 1 VSS VPW nch L=4e-08 W=2.45e-07 
M12 VSS 1 5 VPW nch L=4e-08 W=2.45e-07 
M13 7 6 VSS VPW nch L=4e-08 W=2.45e-07 
M14 VSS 6 7 VPW nch L=4e-08 W=2.45e-07 
M15 7 6 VSS VPW nch L=4e-08 W=2.45e-07 
M16 6 A 8 VPW nch L=4e-08 W=3.7e-07 
M17 8 A 6 VPW nch L=4e-08 W=3.7e-07 
M18 7 9 8 VPW nch L=4e-08 W=3.7e-07 
M19 8 9 7 VPW nch L=4e-08 W=3.7e-07 
M20 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M21 9 A VSS VPW nch L=4e-08 W=2.45e-07 
M22 VSS A 9 VPW nch L=4e-08 W=2.45e-07 
M23 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M24 VSS 8 Y VPW nch L=4e-08 W=3.1e-07 
M25 Y 8 VSS VPW nch L=4e-08 W=3.1e-07 
M26 VSS 8 Y VPW nch L=4e-08 W=3.1e-07 
M27 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M28 1 C VDD VNW pch L=4e-08 W=3.8e-07 
M29 VDD C 1 VNW pch L=4e-08 W=3.8e-07 
M30 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M31 VDD B 4 VNW pch L=4e-08 W=3.8e-07 
M32 4 B VDD VNW pch L=4e-08 W=3.8e-07 
M33 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M34 5 B 6 VNW pch L=4e-08 W=3.8e-07 
M35 6 B 5 VNW pch L=4e-08 W=3.8e-07 
M36 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M37 6 4 1 VNW pch L=4e-08 W=3.8e-07 
M38 1 4 6 VNW pch L=4e-08 W=3.8e-07 
M39 5 1 VDD VNW pch L=4e-08 W=3.8e-07 
M40 VDD 1 5 VNW pch L=4e-08 W=3.8e-07 
M41 5 1 VDD VNW pch L=4e-08 W=3.8e-07 
M42 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M43 VDD 6 7 VNW pch L=4e-08 W=3.8e-07 
M44 7 6 VDD VNW pch L=4e-08 W=3.8e-07 
M45 8 A 7 VNW pch L=4e-08 W=3.8e-07 
M46 7 A 8 VNW pch L=4e-08 W=3.8e-07 
M47 8 A 7 VNW pch L=4e-08 W=3.8e-07 
M48 6 9 8 VNW pch L=4e-08 W=3.8e-07 
M49 8 9 6 VNW pch L=4e-08 W=3.8e-07 
M50 6 9 8 VNW pch L=4e-08 W=3.8e-07 
M51 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M52 9 A VDD VNW pch L=4e-08 W=3.8e-07 
M53 VDD A 9 VNW pch L=4e-08 W=3.8e-07 
M54 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M55 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
M56 Y 8 VDD VNW pch L=4e-08 W=3.8e-07 
M57 VDD 8 Y VNW pch L=4e-08 W=3.8e-07 
.ENDS

