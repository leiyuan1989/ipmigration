* Created:  04/09/2012

.SUBCKT PLVT11LL_CKT DRN GATE SRC BULK 
+ 
.ENDS

.SUBCKT NLVT11LL_CKT DRN GATE SRC BULK 
+ 
.ENDS
****Sub-Circuit for LVT_AD1HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AD1HSV1 A B CI CO S VDD VSS
XX14 m CI net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX18 S net098 VSS VPW NLVT11LL_CKT W=190.00n L=40.00n
XX20 bn B VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX27 net0175 CI net0171 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX28 net0171 m VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 m net43 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX22 cn CI VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX29 net0167 B VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX30 net0175 A net0167 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX32 CO net0175 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX3 net0217 bn net43 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 net0147 B net43 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net0217 A VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX16 net43 cn net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 net0147 net0217 VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX13 m cn net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX17 S net098 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX11 m net43 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX25 net0175 A net0106 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX21 cn CI VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX19 bn B VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX8 net0147 bn net43 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX26 net0175 B net0106 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX24 net0106 m VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX23 net0106 CI VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net0217 B net43 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX31 CO net0175 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX4 net0147 net0217 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX5 net0217 A VDD VNW PLVT11LL_CKT W=400.00n L=40.00n
XX15 net43 CI net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_AD1HSV1
****Sub-Circuit for LVT_ADH1HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_ADH1HSV1 A B CO S VDD VSS
XX18 S net098 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX20 bn B VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX33 net0106 B net0171 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX28 net0171 A VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX32 CO net0106 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX3 net0217 bn net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 net0147 B net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net0217 A VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 net0147 net0217 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX17 S net098 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX19 bn B VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX8 net0147 bn net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX24 net0106 B VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX23 net0106 A VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net0217 B net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX31 CO net0106 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX4 net0147 net0217 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net0217 A VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
.ENDS LVT_ADH1HSV1
****Sub-Circuit for LVT_AND2HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND2HSV1 A1 A2 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_AND2HSV1
****Sub-Circuit for LVT_AND2HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND2HSV2 A1 A2 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_AND2HSV2
****Sub-Circuit for LVT_AND2HSV4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND2HSV4 A1 A2 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=620.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_AND2HSV4
****Sub-Circuit for LVT_AND2HSV8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND2HSV8 A1 A2 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AND2HSV8
****Sub-Circuit for LVT_AND3HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND3HSV1 A1 A2 A3 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=260.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 net_043 A3 VSS VPW NLVT11LL_CKT W=260.00n L=40.00n
XXN1 net18 A2 net_043 VPW NLVT11LL_CKT W=260.00n L=40.00n
XX5 net11 A3 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_AND3HSV1
****Sub-Circuit for LVT_AND3HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND3HSV2 A1 A2 A3 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=260.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 net_043 A3 VSS VPW NLVT11LL_CKT W=260.00n L=40.00n
XXN1 net18 A2 net_043 VPW NLVT11LL_CKT W=260.00n L=40.00n
XX5 net11 A3 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_AND3HSV2
****Sub-Circuit for LVT_AND3HSV4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND3HSV4 A1 A2 A3 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=260.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=620.00n L=40.00n
XX4 net_043 A3 VSS VPW NLVT11LL_CKT W=260.00n L=40.00n
XXN1 net18 A2 net_043 VPW NLVT11LL_CKT W=260.00n L=40.00n
XX5 net11 A3 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_AND3HSV4
****Sub-Circuit for LVT_AND3HSV8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND3HSV8 A1 A2 A3 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX4 net_043 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net_043 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX5 net11 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AND3HSV8
****Sub-Circuit for LVT_AND4HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND4HSV1 A1 A2 A3 A4 Z VDD VSS
XX6 net_042 A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 net_054 A3 net_042 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net_054 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net11 A4 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX5 net11 A3 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_AND4HSV1
****Sub-Circuit for LVT_AND4HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND4HSV2 A1 A2 A3 A4 Z VDD VSS
XX6 net_042 A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 net_054 A3 net_042 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net_054 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net11 A4 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX5 net11 A3 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_AND4HSV2
****Sub-Circuit for LVT_AND4HSV4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND4HSV4 A1 A2 A3 A4 Z VDD VSS
XX6 net_042 A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=620.00n L=40.00n
XX4 net_054 A3 net_042 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net_054 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net11 A4 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX5 net11 A3 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_AND4HSV4
****Sub-Circuit for LVT_AND4HSV8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AND4HSV8 A1 A2 A3 A4 Z VDD VSS
XX6 net_042 A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX4 net_054 A3 net_042 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net_054 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net11 A4 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net11 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AND4HSV8
****Sub-Circuit for LVT_AOI211HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI211HSV1 A1 A2 B C ZN VDD VSS
XX6 ZN B VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 net4 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN C VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net4 A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net3 A1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net3 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net2 B net3 VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN C net2 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_AOI211HSV1
****Sub-Circuit for LVT_AOI211HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI211HSV2 A1 A2 B C ZN VDD VSS
XX6 ZN B VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net4 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN C VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net4 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net3 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net3 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net2 B net3 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN C net2 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AOI211HSV2
****Sub-Circuit for LVT_AOI21HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI21HSV1 A1 A2 B ZN VDD VSS
XX6 ZN B VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 net4 VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net4 A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net3 A1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net3 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN B net3 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_AOI21HSV1
****Sub-Circuit for LVT_AOI21HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI21HSV2 A1 A2 B ZN VDD VSS
XX6 ZN B VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net4 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net4 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net3 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net3 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 ZN B net3 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AOI21HSV2
****Sub-Circuit for LVT_AOI221HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI221HSV1 A1 A2 B1 B2 C ZN VDD VSS
XX6 ZN C VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 N3 B2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 N14 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN B1 N3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 N14 A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 N9 B1 N11 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX7 N11 A1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 N11 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 N9 B2 N11 VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN C N9 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_AOI221HSV1
****Sub-Circuit for LVT_AOI221HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI221HSV2 A1 A2 B1 B2 C ZN VDD VSS
XX6 ZN C VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 N3 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 N14 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B1 N3 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 N14 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 N9 B1 N11 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX7 N11 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 N11 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 N9 B2 N11 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN C N9 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AOI221HSV2
****Sub-Circuit for LVT_AOI222HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI222HSV1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX6 ZN C1 net4 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX10 net4 C2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 net5 B2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 net6 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN B1 net5 VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net6 A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 net2 B2 net1 VNW PLVT11LL_CKT W=310.0n L=40.00n
XX11 ZN A2 net2 VNW PLVT11LL_CKT W=310.0n L=40.00n
XX7 net1 C1 VDD VNW PLVT11LL_CKT W=310.0n L=40.00n
XX5 net1 C2 VDD VNW PLVT11LL_CKT W=310.0n L=40.00n
XX0 net2 B1 net1 VNW PLVT11LL_CKT W=310.0n L=40.00n
XXP1 ZN A1 net2 VNW PLVT11LL_CKT W=310.0n L=40.00n
.ENDS LVT_AOI222HSV1
****Sub-Circuit for LVT_AOI222HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI222HSV2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX6 ZN C1 net4 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX10 net4 C2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 net5 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net6 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B1 net5 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net6 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 net2 B2 net1 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX11 ZN A2 net2 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX7 net1 C1 VDD VNW PLVT11LL_CKT W=455.0n L=40.00n
XX5 net1 C2 VDD VNW PLVT11LL_CKT W=455.0n L=40.00n
XX0 net2 B1 net1 VNW PLVT11LL_CKT W=455.0n L=40.00n
XXP1 ZN A1 net2 VNW PLVT11LL_CKT W=455.0n L=40.00n
.ENDS LVT_AOI222HSV2
****Sub-Circuit for LVT_AOI22HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI22HSV1 A1 A2 B1 B2 ZN VDD VSS
XX9 N64 B2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 N49 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN B1 N64 VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 N49 A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 ZN B2 N69 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX7 N69 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 N69 A1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN B1 N69 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_AOI22HSV1
****Sub-Circuit for LVT_AOI22HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI22HSV2 A1 A2 B1 B2 ZN VDD VSS
XX9 N64 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 N49 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B1 N64 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 N49 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 ZN B2 N69 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX7 N69 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 N69 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 ZN B1 N69 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AOI22HSV2
****Sub-Circuit for LVT_AOI31HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI31HSV1 A1 A2 A3 B ZN VDD VSS
XX6 ZN B VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 net3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 net4 A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net3 A2 net4 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 net1 A3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX7 net1 A1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net1 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN B net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_AOI31HSV1
****Sub-Circuit for LVT_AOI31HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI31HSV2 A1 A2 A3 B ZN VDD VSS
XX6 ZN B VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net3 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 net4 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net3 A2 net4 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 net1 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX7 net1 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net1 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 ZN B net1 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AOI31HSV2
****Sub-Circuit for LVT_AOI32HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI32HSV1 A1 A2 A3 B1 B2 ZN VDD VSS
XX6 ZN B1 net5 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 net3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 net4 A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX11 net5 B2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net3 A2 net4 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 net1 A3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX10 ZN B2 net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX7 net1 A1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net1 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN B1 net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_AOI32HSV1
****Sub-Circuit for LVT_AOI32HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI32HSV2 A1 A2 A3 B1 B2 ZN VDD VSS
XX6 ZN B1 net5 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net3 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 net4 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX11 net5 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net3 A2 net4 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 net1 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX10 ZN B2 net1 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX7 net1 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net1 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 ZN B1 net1 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AOI32HSV2
****Sub-Circuit for LVT_AOI33HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI33HSV1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX12 net_69 B3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 ZN B1 net5 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 net3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 net4 A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX11 net5 B2 net_69 VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net3 A2 net4 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 net1 A3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX10 ZN B2 net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX7 net1 A1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net1 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX13 ZN B3 net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN B1 net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_AOI33HSV1
****Sub-Circuit for LVT_AOI33HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_AOI33HSV2 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX12 net_69 B3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 ZN B1 net5 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net3 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 net4 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX11 net5 B2 net_69 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net3 A2 net4 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 net1 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX10 ZN B2 net1 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX7 net1 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net1 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX13 ZN B3 net1 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 ZN B1 net1 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_AOI33HSV2
****Sub-Circuit for LVT_BUFHSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV1 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_BUFHSV1
****Sub-Circuit for LVT_BUFHSV12, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV12 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=1.86u L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=720.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=2.73u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=1.08u L=40.00n
.ENDS LVT_BUFHSV12
****Sub-Circuit for LVT_BUFHSV16, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV16 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=2.48u L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=930.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=3.64u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=1.365u L=40.00n
.ENDS LVT_BUFHSV16
****Sub-Circuit for LVT_BUFHSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV2 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_BUFHSV2
****Sub-Circuit for LVT_BUFHSV20, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV20 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=3.1u L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=4.55u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
.ENDS LVT_BUFHSV20
****Sub-Circuit for LVT_BUFHSV24, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV24 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=3.72u L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=1.55u L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=5.46u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=2.275u L=40.00n
.ENDS LVT_BUFHSV24
****Sub-Circuit for LVT_BUFHSV3, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV3 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=190.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=700.00n L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_BUFHSV3
****Sub-Circuit for LVT_BUFHSV4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV4 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=620.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=240.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
.ENDS LVT_BUFHSV4
****Sub-Circuit for LVT_BUFHSV6, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV6 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=930.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=1.365u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_BUFHSV6
****Sub-Circuit for LVT_BUFHSV8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_BUFHSV8 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=480.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=740.00n L=40.00n
.ENDS LVT_BUFHSV8
****Sub-Circuit for LVT_CKMUX2HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CKMUX2HSV1 I0 I1 S Z VDD VSS
XX47 net41 S net64 VPW NLVT11LL_CKT W=270.00n L=40.00n
XX51 Z net64 VSS VPW NLVT11LL_CKT W=180.00n L=40.00n
XX49 net39 I0 VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX31 net41 I1 VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX53 net43 S VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX36 net39 net43 net64 VPW NLVT11LL_CKT W=270.00n L=40.00n
XX50 net39 I0 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX52 Z net64 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX48 net41 net43 net64 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX32 net41 I1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 net43 S VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX39 net39 S net64 VNW PLVT11LL_CKT W=300.00n L=40.00n
.ENDS LVT_CKMUX2HSV1
****Sub-Circuit for LVT_CKMUX2HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CKMUX2HSV2 I0 I1 S Z VDD VSS
XX47 net41 S net64 VPW NLVT11LL_CKT W=270n L=40.00n
XX51 Z net64 VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XX49 net39 I0 VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX31 net41 I1 VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX53 net43 S VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX36 net39 net43 net64 VPW NLVT11LL_CKT W=270.00n L=40.00n
XX50 net39 I0 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX52 Z net64 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX48 net41 net43 net64 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX32 net41 I1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 net43 S VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX39 net39 S net64 VNW PLVT11LL_CKT W=300.00n L=40.00n
.ENDS LVT_CKMUX2HSV2
****Sub-Circuit for LVT_CLKAND2HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKAND2HSV1 A1 A2 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=180.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_CLKAND2HSV1
****Sub-Circuit for LVT_CLKAND2HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKAND2HSV2 A1 A2 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_CLKAND2HSV2
****Sub-Circuit for LVT_CLKAND2HSV4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKAND2HSV4 A1 A2 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=620.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=1.365u L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_CLKAND2HSV4
****Sub-Circuit for LVT_CLKAND2HSV8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKAND2HSV8 A1 A2 Z VDD VSS
XX1 net11 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net11 VSS VPW NLVT11LL_CKT W=1.215u L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 Z net11 VDD VNW PLVT11LL_CKT W=2.73u L=40.00n
XX0 net11 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net11 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_CLKAND2HSV8
****Sub-Circuit for LVT_CLKBUFHSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV1 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=180.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_CLKBUFHSV1
****Sub-Circuit for LVT_CLKBUFHSV12, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV12 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=1.35u L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=450.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=2.73u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
.ENDS LVT_CLKBUFHSV12
****Sub-Circuit for LVT_CLKBUFHSV16, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV16 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=1.8u L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=590.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=3.64u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=1.2u L=40.00n
.ENDS LVT_CLKBUFHSV16
****Sub-Circuit for LVT_CLKBUFHSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV2 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_CLKBUFHSV2
****Sub-Circuit for LVT_CLKBUFHSV20, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV20 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=2.295u L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=765.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=4.55u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=1.6u L=40.00n
.ENDS LVT_CLKBUFHSV20
****Sub-Circuit for LVT_CLKBUFHSV24, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV24 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=2.7u L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=900.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=5.46u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
.ENDS LVT_CLKBUFHSV24
****Sub-Circuit for LVT_CLKBUFHSV3, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV3 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=380.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=190.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=700.00n L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=350.00n L=40.00n
.ENDS LVT_CLKBUFHSV3
****Sub-Circuit for LVT_CLKBUFHSV4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV4 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=500.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=260.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=445.00n L=40.00n
.ENDS LVT_CLKBUFHSV4
****Sub-Circuit for LVT_CLKBUFHSV6, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV6 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=720.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=240.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=1.365u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_CLKBUFHSV6
****Sub-Circuit for LVT_CLKBUFHSV8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKBUFHSV8 I Z VDD VSS
XX2 Z net7 VSS VPW NLVT11LL_CKT W=930.00n L=40.00n
XX0 net7 I VSS VPW NLVT11LL_CKT W=300.00n L=40.00n
XX3 Z net7 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX1 net7 I VDD VNW PLVT11LL_CKT W=610.00n L=40.00n
.ENDS LVT_CLKBUFHSV8
****Sub-Circuit for LVT_CLKLANQHSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV1 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=200.00n L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=155.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=320.00n L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=155.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV1
****Sub-Circuit for LVT_CLKLANQHSV12, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV12 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=1.86u L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=2.73u L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV12
****Sub-Circuit for LVT_CLKLANQHSV16, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV16 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=2.48u L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=3.64u L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV16
****Sub-Circuit for LVT_CLKLANQHSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV2 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV2
****Sub-Circuit for LVT_CLKLANQHSV20, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV20 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=3.1u L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=4.55u L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV20
****Sub-Circuit for LVT_CLKLANQHSV24, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV24 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=155.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=3.72u L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=155.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=5.46u L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV24
****Sub-Circuit for LVT_CLKLANQHSV3, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV3 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=440.00n L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=670.00n L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV3
****Sub-Circuit for LVT_CLKLANQHSV4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV4 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=560.00n L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV4
****Sub-Circuit for LVT_CLKLANQHSV6, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV6 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=795.00n L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=1.365u L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV6
****Sub-Circuit for LVT_CLKLANQHSV8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKLANQHSV8 CK E Q TE VDD VSS
XX6 net0112 TE VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX9 net0112 E VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX52 nt12 net076 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX1 c cn VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX2 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Q net0106 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX36 net0128 c nt12 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net0106 c net068 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net068 net076 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net076 net0128 VSS VPW NLVT11LL_CKT W=225.00n L=40.00n
XX15 net0128 cn net0112 VPW NLVT11LL_CKT W=225.00n L=40.00n
XX17 net0128 c net170 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX0 net076 net0128 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX53 nt11 net076 VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 c cn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 cn CK VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 Q net0106 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX39 net0128 cn nt11 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX18 net0106 c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net0106 net076 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0171 TE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX10 net170 E net0171 VNW PLVT11LL_CKT W=280.00n L=40.00n
.ENDS LVT_CLKLANQHSV8
****Sub-Circuit for LVT_CLKNAND2HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNAND2HSV1 A1 A2 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=280.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
.ENDS LVT_CLKNAND2HSV1
****Sub-Circuit for LVT_CLKNAND2HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNAND2HSV2 A1 A2 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=330.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=330.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_CLKNAND2HSV2
****Sub-Circuit for LVT_CLKNAND2HSV3, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNAND2HSV3 A1 A2 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=440.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=440.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
.ENDS LVT_CLKNAND2HSV3
****Sub-Circuit for LVT_CLKNAND2HSV4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNAND2HSV4 A1 A2 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=600.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=600.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
.ENDS LVT_CLKNAND2HSV4
****Sub-Circuit for LVT_CLKNAND2HSV8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNAND2HSV8 A1 A2 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=1.2u L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=1.2u L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
.ENDS LVT_CLKNAND2HSV8
****Sub-Circuit for LVT_CLKNHSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV1 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=180.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=315.0n L=40.00n
.ENDS LVT_CLKNHSV1
****Sub-Circuit for LVT_CLKNHSV12, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV12 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=1.3u L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=2.73u L=40.00n
.ENDS LVT_CLKNHSV12
****Sub-Circuit for LVT_CLKNHSV16, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV16 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=1.86u L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=3.64u L=40.00n
.ENDS LVT_CLKNHSV16
****Sub-Circuit for LVT_CLKNHSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV2 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=455.0n L=40.00n
.ENDS LVT_CLKNHSV2
****Sub-Circuit for LVT_CLKNHSV20, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV20 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=2.32u L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=4.55u L=40.00n
.ENDS LVT_CLKNHSV20
****Sub-Circuit for LVT_CLKNHSV24, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV24 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=2.695u L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=5.46u L=40.00n
.ENDS LVT_CLKNHSV24
****Sub-Circuit for LVT_CLKNHSV3, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV3 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=400.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=700.0n L=40.00n
.ENDS LVT_CLKNHSV3
****Sub-Circuit for LVT_CLKNHSV4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV4 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=490.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
.ENDS LVT_CLKNHSV4
****Sub-Circuit for LVT_CLKNHSV6, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV6 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=720.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=1.365u L=40.00n
.ENDS LVT_CLKNHSV6
****Sub-Circuit for LVT_CLKNHSV8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKNHSV8 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=915.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
.ENDS LVT_CLKNHSV8
****Sub-Circuit for LVT_CLKXOR2HSV1, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKXOR2HSV1 A1 A2 Z VDD VSS
XX57 Z xna1a2 VSS VPW NLVT11LL_CKT W=180.00n L=40.00n
XX47 a2n a1n xna1a2 VPW NLVT11LL_CKT W=280.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX55 a2nn a2n VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX36 a2nn A1 xna1a2 VPW NLVT11LL_CKT W=280.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX58 Z xna1a2 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX48 a2n A1 xna1a2 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX56 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX39 a2nn a1n xna1a2 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_CLKXOR2HSV1
****Sub-Circuit for LVT_CLKXOR2HSV2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_CLKXOR2HSV2 A1 A2 Z VDD VSS
XX57 Z xna1a2 VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XX47 a2n a1n xna1a2 VPW NLVT11LL_CKT W=280.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX55 a2nn a2n VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX36 a2nn A1 xna1a2 VPW NLVT11LL_CKT W=280.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX58 Z xna1a2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX48 a2n A1 xna1a2 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX56 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX39 a2nn a1n xna1a2 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_CLKXOR2HSV2
****Sub-Circuit for LVT_DELHS2, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_DELHS2 I Z VDD VSS
XX9 net040 net026 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX4 net026 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX5 net050 net026 net040 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 net13 net050 net048 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX11 net048 net050 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net13 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 net071 net026 VDD VNW PLVT11LL_CKT W=210.0n L=40.00n
XX6 net026 I VDD VNW PLVT11LL_CKT W=210.0n L=40.00n
XX7 net050 net026 net071 VNW PLVT11LL_CKT W=210.0n L=40.00n
XX1 net13 net050 net091 VNW PLVT11LL_CKT W=210.0n L=40.00n
XX10 net091 net050 VDD VNW PLVT11LL_CKT W=210.0n L=40.00n
XX3 Z net13 VDD VNW PLVT11LL_CKT W=455.0n L=40.00n
.ENDS LVT_DELHS2
****Sub-Circuit for LVT_DHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DHSV1 CK D Q QN VDD VSS
XX8 net122 D VDD VNW PLVT11LL_CKT W=235.00n L=40.00n
XX1 net163 net171 VDD VNW PLVT11LL_CKT W=400.00n L=40.00n
XX43 Q s VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX2 net163 cn net210 VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net139 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net139 c net210 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 QN net210 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX18 s net210 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net127 cn net171 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net163 net127 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX10 net171 c net122 VNW PLVT11LL_CKT W=235.00n L=40.00n
XX42 Q s VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net167 D VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX0 net163 net171 VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX3 net163 c net210 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net194 cn net210 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net194 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 QN net210 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX17 s net210 VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net178 c net171 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS net163 net178 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX9 net171 cn net167 VPW NLVT11LL_CKT W=220.00n L=40.00n
.ENDS LVT_DHSV1
****Sub-Circuit for LVT_DHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DHSV2 CK D Q QN VDD VSS
XX42 Q s VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net0217 c net43 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn net43 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 QN net43 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 s net43 VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net52 c net0204 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS net0217 net52 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX9 net0204 cn net69 VPW NLVT11LL_CKT W=220.00n L=40.00n
XX7 net69 D VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX0 net0217 net0204 VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX43 Q s VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net0217 cn net43 VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c net43 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 QN net43 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 s net43 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn net0204 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net0217 net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX10 net0204 c net128 VNW PLVT11LL_CKT W=235.00n L=40.00n
XX8 net128 D VDD VNW PLVT11LL_CKT W=235.00n L=40.00n
XX1 net0217 net0204 VDD VNW PLVT11LL_CKT W=400.00n L=40.00n
.ENDS LVT_DHSV2
****Sub-Circuit for LVT_DQHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DQHSV1 CK D Q VDD VSS
XX8 net111 D VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX1 net148 net156 VDD VNW PLVT11LL_CKT W=400.00n L=40.00n
XX43 Q s VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX2 net148 cn net191 VNW PLVT11LL_CKT W=260.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=400.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net124 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net124 c net191 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX18 s net191 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net116 cn net156 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net148 net116 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX5 net156 c net111 VNW PLVT11LL_CKT W=250.00n L=40.00n
XX42 Q s VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net152 D VSS VPW NLVT11LL_CKT W=240.00n L=40.00n
XX0 net148 net156 VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XX3 net148 c net191 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net175 cn net191 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net175 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX17 s net191 VSS VPW NLVT11LL_CKT W=200.00n L=40.00n
XX12 net163 c net156 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS net148 net163 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX9 net156 cn net152 VPW NLVT11LL_CKT W=240.00n L=40.00n
.ENDS LVT_DQHSV1
****Sub-Circuit for LVT_DQHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DQHSV2 CK D Q VDD VSS
XX42 Q s VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net0217 c net43 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn net43 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX17 s net43 VSS VPW NLVT11LL_CKT W=200.00n L=40.00n
XX12 net52 c net0181 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS net0217 net52 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX9 net0181 cn net69 VPW NLVT11LL_CKT W=240.00n L=40.00n
XX7 net69 D VSS VPW NLVT11LL_CKT W=240.00n L=40.00n
XX0 net0217 net0181 VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XX43 Q s VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net0217 cn net43 VNW PLVT11LL_CKT W=260.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=400.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c net43 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX18 s net43 VDD VNW PLVT11LL_CKT W=390.00n L=40.00n
XX14 net117 cn net0181 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net0217 net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX5 net0181 c net128 VNW PLVT11LL_CKT W=260.00n L=40.00n
XX8 net128 D VDD VNW PLVT11LL_CKT W=260.00n L=40.00n
XX1 net0217 net0181 VDD VNW PLVT11LL_CKT W=400.00n L=40.00n
.ENDS LVT_DQHSV2
****Sub-Circuit for LVT_DRNHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DRNHSV1 CK D Q QN RDN VDD VSS
XX21 net128 c net135 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX8 net128 RDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX1 net184 net128 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX43 Q net144 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 net135 D VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX19 QN net231 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX2 net184 cn net231 VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD net144 net152 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net152 c net231 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX15 net144 RDN VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX18 net144 net231 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net140 cn net128 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net184 net140 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX42 Q net144 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net188 RDN VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XX0 net184 net128 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX20 QN net231 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX16 net144 RDN net208 VPW NLVT11LL_CKT W=220.00n L=40.00n
XX6 net128 cn net192 VPW NLVT11LL_CKT W=250.00n L=40.00n
XX3 net184 c net231 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net215 cn net231 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net144 net215 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX17 net208 net231 VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX10 VSS RDN net207 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX12 net199 c net128 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net207 net184 net199 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net192 D net188 VPW NLVT11LL_CKT W=250.00n L=40.00n
.ENDS LVT_DRNHSV1
****Sub-Circuit for LVT_DRNHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DRNHSV2 CK D Q QN RDN VDD VSS
XX42 Q net0117 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX20 QN net43 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net0117 RDN net0108 VPW NLVT11LL_CKT W=220.00n L=40.00n
XX6 net0177 cn net0181 VPW NLVT11LL_CKT W=250.00n L=40.00n
XX3 net0217 c net43 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn net43 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net0117 net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX17 net0108 net43 VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX10 VSS RDN net0161 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX12 net52 c net0177 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net0161 net0217 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net0181 D net69 VPW NLVT11LL_CKT W=250.00n L=40.00n
XX7 net69 RDN VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XX0 net0217 net0177 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX43 Q net0117 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net128 D VDD VNW PLVT11LL_CKT W=230.00n L=40.00n
XX19 QN net43 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net0217 cn net43 VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD net0117 net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c net43 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX15 net0117 RDN VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX18 net0117 net43 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn net0177 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net0217 net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX21 net0177 c net128 VNW PLVT11LL_CKT W=230.00n L=40.00n
XX8 net0177 RDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX1 net0217 net0177 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
.ENDS LVT_DRNHSV2
****Sub-Circuit for LVT_DRNQHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DRNQHSV1 CK D Q RDN VDD VSS
XX19 net117 c net124 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX8 net117 RDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX1 net169 net117 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX43 Q net133 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 net124 D VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX2 net169 cn net216 VNW PLVT11LL_CKT W=305.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD net133 net141 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net141 c net216 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX15 net133 RDN VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX18 net133 net216 VDD VNW PLVT11LL_CKT W=350.00n L=40.00n
XX14 net129 cn net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net169 net129 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX42 Q net133 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net173 RDN VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XX0 net169 net117 VSS VPW NLVT11LL_CKT W=265.00n L=40.00n
XX16 net133 RDN net193 VPW NLVT11LL_CKT W=270.00n L=40.00n
XX6 net117 cn net177 VPW NLVT11LL_CKT W=250.00n L=40.00n
XX3 net169 c net216 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net200 cn net216 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net133 net200 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX17 net193 net216 VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX10 VSS RDN net192 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX12 net184 c net117 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net192 net169 net184 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net177 D net173 VPW NLVT11LL_CKT W=250.00n L=40.00n
.ENDS LVT_DRNQHSV1
****Sub-Circuit for LVT_DRNQHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DRNQHSV2 CK D Q RDN VDD VSS
XX42 Q net0117 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net0117 RDN net0108 VPW NLVT11LL_CKT W=270.00n L=40.00n
XX6 net0177 cn net0181 VPW NLVT11LL_CKT W=250.00n L=40.00n
XX3 net0217 c net43 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn net43 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS net0117 net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX17 net0108 net43 VSS VPW NLVT11LL_CKT W=270.00n L=40.00n
XX10 VSS RDN net0161 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX12 net52 c net0177 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net0161 net0217 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net0181 D net69 VPW NLVT11LL_CKT W=250.00n L=40.00n
XX7 net69 RDN VSS VPW NLVT11LL_CKT W=250.00n L=40.00n
XX0 net0217 net0177 VSS VPW NLVT11LL_CKT W=265.00n L=40.00n
XX43 Q net0117 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net128 D VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX2 net0217 cn net43 VNW PLVT11LL_CKT W=305.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD net0117 net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c net43 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX15 net0117 RDN VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX18 net0117 net43 VDD VNW PLVT11LL_CKT W=350.00n L=40.00n
XX14 net117 cn net0177 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net0217 net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX19 net0177 c net128 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX8 net0177 RDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX1 net0217 net0177 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
.ENDS LVT_DRNQHSV2
****Sub-Circuit for LVT_DRSNHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DRSNHSV1 CK D Q QN RDN SDN VDD VSS
XX5 net147 c net154 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX8 net147 RDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX32 net143 net147 VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX39 VDD SDN net258 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX43 Q net263 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 net154 D VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX31 net143 SDN VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX19 QN net258 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX21 n RDN VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX40 net187 c net258 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX2 net143 cn net258 VNW PLVT11LL_CKT W=265.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD n net167 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX25 net167 net263 net187 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX41 net263 net258 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net159 cn net147 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net143 net159 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX44 net287 net263 net238 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net219 D net215 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX45 net258 cn net287 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX38 net238 SDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net215 RDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX42 Q net263 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX20 QN net258 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX22 n RDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX47 net263 net258 VSS VPW NLVT11LL_CKT W=315.00n L=40.00n
XX6 net147 cn net219 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX3 net143 c net258 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX33 net143 SDN net247 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX34 net247 net147 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=235.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 net258 n net238 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX10 VSS RDN net234 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX12 net226 c net147 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net234 net143 net226 VPW NLVT11LL_CKT W=150.00n L=40.00n
.ENDS LVT_DRSNHSV1
****Sub-Circuit for LVT_DRSNHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DRSNHSV2 CK D Q QN RDN SDN VDD VSS
XX44 net0224 net0226 net0381 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX45 net0320 cn net0224 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX38 net0381 SDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX42 Q net0226 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX20 QN net0320 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX22 n RDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX47 net0226 net0320 VSS VPW NLVT11LL_CKT W=315.00n L=40.00n
XX6 net0177 cn net0181 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX3 net0217 c net0320 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX33 net0217 SDN net0211 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX34 net0211 net0177 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=235.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 net0320 n net0381 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX10 VSS RDN net0161 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX12 net52 c net0177 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net0161 net0217 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net0181 D net69 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX7 net69 RDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX39 VDD SDN net0320 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX43 Q net0226 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net128 D VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX31 net0217 SDN VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX19 QN net0320 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX21 n RDN VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX40 net0305 c net0320 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX2 net0217 cn net0320 VNW PLVT11LL_CKT W=265.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD n net109 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX25 net109 net0226 net0305 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX41 net0226 net0320 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn net0177 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net0217 net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX5 net0177 c net128 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX8 net0177 RDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX32 net0217 net0177 VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
.ENDS LVT_DRSNHSV2
****Sub-Circuit for LVT_DSNHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DSNHSV1 CK D Q QN SDN VDD VSS
XX13 VDD net122 net134 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX5 net218 c net129 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX45 net178 c net209 VNW PLVT11LL_CKT W=130.00n L=40.00n
XX32 net122 net218 VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX43 Q net214 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 net129 D VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX31 net122 SDN VDD VNW PLVT11LL_CKT W=355.00n L=40.00n
XX19 QN net209 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX2 net122 cn net209 VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX44 VDD net214 net178 VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD SDN net209 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX41 net214 net209 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net134 cn net218 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS net122 net185 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX49 net238 net214 net230 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX50 net209 cn net238 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX38 net230 SDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX42 Q net214 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX20 QN net209 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX51 net218 cn net210 VPW NLVT11LL_CKT W=145.00n L=40.00n
XX47 net214 net209 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX48 net210 D VSS VPW NLVT11LL_CKT W=145.00n L=40.00n
XX3 net122 c net209 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX33 net122 SDN net198 VPW NLVT11LL_CKT W=285.00n L=40.00n
XX34 net198 net218 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX12 net185 c net218 VPW NLVT11LL_CKT W=120.00n L=40.00n
.ENDS LVT_DSNHSV1
****Sub-Circuit for LVT_DSNHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DSNHSV2 CK D Q QN SDN VDD VSS
XX49 net0188 net0226 net0381 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX50 net0320 cn net0188 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX38 net0381 SDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX42 Q net0226 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX20 QN net0320 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX51 net69 cn net0187 VPW NLVT11LL_CKT W=145.00n L=40.00n
XX47 net0226 net0320 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX48 net0187 D VSS VPW NLVT11LL_CKT W=145.00n L=40.00n
XX3 net0217 c net0320 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX33 net0217 SDN net0211 VPW NLVT11LL_CKT W=285.00n L=40.00n
XX34 net0211 net69 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX12 net52 c net69 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS net0217 net52 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX45 net0128 c net0320 VNW PLVT11LL_CKT W=130.00n L=40.00n
XX43 Q net0226 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net128 D VDD VNW PLVT11LL_CKT W=220.00n L=40.00n
XX31 net0217 SDN VDD VNW PLVT11LL_CKT W=355.00n L=40.00n
XX19 QN net0320 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net0217 cn net0320 VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX44 VDD net0226 net0128 VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD SDN net0320 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX41 net0226 net0320 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn net69 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net0217 net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX5 net69 c net128 VNW PLVT11LL_CKT W=220.00n L=40.00n
XX32 net0217 net69 VDD VNW PLVT11LL_CKT W=290.00n L=40.00n
.ENDS LVT_DSNHSV2
****Sub-Circuit for LVT_DXHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DXHSV1 CK DA DB Q QN SA VDD VSS
XX8 net191 SA VDD VNW PLVT11LL_CKT W=220.00n L=40.00n
XX1 net200 net256 VDD VNW PLVT11LL_CKT W=330.00n L=40.00n
XX43 Q s VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 sn SA VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 net188 sn net191 VNW PLVT11LL_CKT W=220.00n L=40.00n
XX16 net188 DB net191 VNW PLVT11LL_CKT W=220.00n L=40.00n
XX2 net200 cn net255 VNW PLVT11LL_CKT W=285.00n L=40.00n
XX22 net256 c net188 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net160 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net160 c net255 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 QN net255 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX18 s net255 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net148 cn net256 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net200 net148 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX10 net191 DA VDD VNW PLVT11LL_CKT W=220.00n L=40.00n
XX42 Q s VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net204 SA VSS VPW NLVT11LL_CKT W=170.00n L=40.00n
XX0 net200 net256 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX5 sn SA VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX31 net256 cn net216 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX3 net200 c net255 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net239 cn net255 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net239 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 QN net255 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX17 s net255 VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net223 c net256 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS net200 net223 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX9 net216 DA net204 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX15 net212 DB VSS VPW NLVT11LL_CKT W=170.00n L=40.00n
XX6 net216 sn net212 VPW NLVT11LL_CKT W=170.00n L=40.00n
.ENDS LVT_DXHSV1
****Sub-Circuit for LVT_DXHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_DXHSV2 CK DA DB Q QN SA VDD VSS
XX42 Q s VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX5 sn SA VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX31 net0207 cn net0216 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX3 net0260 c net43 VPW NLVT11LL_CKT W=230.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn net43 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 QN net43 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 s net43 VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net52 c net0207 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS net0260 net52 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX9 net0216 DA net69 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX15 net0296 DB VSS VPW NLVT11LL_CKT W=170.00n L=40.00n
XX6 net0216 sn net0296 VPW NLVT11LL_CKT W=170.00n L=40.00n
XX7 net69 SA VSS VPW NLVT11LL_CKT W=170.00n L=40.00n
XX0 net0260 net0207 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX43 Q s VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 sn SA VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 net0143 sn net128 VNW PLVT11LL_CKT W=230.00n L=40.00n
XX16 net0143 DB net128 VNW PLVT11LL_CKT W=230.00n L=40.00n
XX2 net0260 cn net43 VNW PLVT11LL_CKT W=285.00n L=40.00n
XX22 net0207 c net0143 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c net43 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 QN net43 VDD VNW PLVT11LL_CKT W=450.00n L=40.00n
XX18 s net43 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn net0207 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD net0260 net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX10 net128 DA VDD VNW PLVT11LL_CKT W=230.00n L=40.00n
XX8 net128 SA VDD VNW PLVT11LL_CKT W=230.00n L=40.00n
XX1 net0260 net0207 VDD VNW PLVT11LL_CKT W=330.00n L=40.00n
.ENDS LVT_DXHSV2
****Sub-Circuit for LVT_FDCAPHS16, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_FDCAPHS16 VDD VSS
XX1 VSS net3 net4 VPW NLVT11LL_CKT W=300.0n L=40.00n m=11
XX0 net3 net4 VDD VNW PLVT11LL_CKT W=340.00n L=40n m=11
.ENDS LVT_FDCAPHS16
****Sub-Circuit for LVT_FDCAPHS32, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_FDCAPHS32 VDD VSS
XX1 VSS net7 net8 VPW NLVT11LL_CKT W=300.0n L=40.00n m=23
XX0 net7 net8 VDD VNW PLVT11LL_CKT W=340.00n L=40.00n m=23
.ENDS LVT_FDCAPHS32
****Sub-Circuit for LVT_FDCAPHS4, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_FDCAPHS4 VDD VSS
XX1 VSS net7 net8 VPW NLVT11LL_CKT W=285.000n L=80.00n
XX0 net7 net8 VDD VNW PLVT11LL_CKT W=350.00n L=80.00n
.ENDS LVT_FDCAPHS4
****Sub-Circuit for LVT_FDCAPHS64, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_FDCAPHS64 VDD VSS
XX1 VSS net7 net8 VPW NLVT11LL_CKT W=300.0n L=40.00n m=48
XX0 net7 net8 VDD VNW PLVT11LL_CKT W=340.00n L=40.00n m=48
.ENDS LVT_FDCAPHS64
****Sub-Circuit for LVT_FDCAPHS8, Wed Sep  5 13:54:26 CST 2012****
.SUBCKT LVT_FDCAPHS8 VDD VSS
XX1 VSS net7 net8 VPW NLVT11LL_CKT W=300.0n L=40.00n m=5
XX0 net7 net8 VDD VNW PLVT11LL_CKT W=340.00n L=40.00n m=5
.ENDS LVT_FDCAPHS8
****Sub-Circuit for LVT_FILLTIEHS, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_FILLTIEHS VDD VSS
.ENDS LVT_FILLTIEHS
****Sub-Circuit for LVT_F_DIODEHS2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_F_DIODEHS2 A VDD VSS
DD1 A VNW PDIO11LLLVT PJ=1.36u AREA=0.0756p 
DD0 VPW A NDIO11LLLVT PJ=1.08u AREA=0.056p
.ENDS LVT_F_DIODEHS2
****Sub-Circuit for LVT_F_DIODEHS4, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_F_DIODEHS4 A VDD VSS
DD1 A VNW PDIO11LLLVT PJ=2.68u AREA=0.1824p 
DD0 VPW A NDIO11LLLVT PJ=2.12u AREA=0.1292p
.ENDS LVT_F_DIODEHS4
****Sub-Circuit for LVT_F_DIODEHS8, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_F_DIODEHS8 A VDD VSS
DD1 A VNW PDIO11LLLVT PJ=6.48u AREA=0.4032p 
DD0 VPW A NDIO11LLLVT PJ=5.08u AREA=0.2856p
.ENDS LVT_F_DIODEHS8
****Sub-Circuit for LVT_F_FILLHS1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_F_FILLHS1 VDD VSS
.ENDS LVT_F_FILLHS1
****Sub-Circuit for LVT_F_FILLHS16, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_F_FILLHS16 VDD VSS
.ENDS LVT_F_FILLHS16
****Sub-Circuit for LVT_F_FILLHS2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_F_FILLHS2 VDD VSS
.ENDS LVT_F_FILLHS2
****Sub-Circuit for LVT_F_FILLHS4, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_F_FILLHS4 VDD VSS
.ENDS LVT_F_FILLHS4
****Sub-Circuit for LVT_F_FILLHS8, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_F_FILLHS8 VDD VSS
.ENDS LVT_F_FILLHS8
****Sub-Circuit for LVT_I2NAND4HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_I2NAND4HSV1 A1 A2 B1 B2 ZN VDD VSS
XX9 a2n A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX6 a1n A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 net031 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN a1n net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net039 B1 net031 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 a2n net039 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 a2n A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX7 a1n A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN B2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 ZN B1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN a1n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_I2NAND4HSV1
****Sub-Circuit for LVT_I2NAND4HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_I2NAND4HSV2 A1 A2 B1 B2 ZN VDD VSS
XX9 a2n A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX6 a1n A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 net031 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN a1n net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net039 B1 net031 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 a2n net039 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 a2n A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX7 a1n A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN B2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX5 ZN B1 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX0 ZN a2n VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XXP1 ZN a1n VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
.ENDS LVT_I2NAND4HSV2
****Sub-Circuit for LVT_I2NOR4HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_I2NOR4HSV1 A1 A2 B1 B2 ZN VDD VSS
XX9 a2n A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX6 a1n A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 ZN B2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN a1n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 ZN B1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 ZN a2n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 a2n A2 VDD VNW PLVT11LL_CKT W=210.0n L=40.00n
XX7 a1n A1 VDD VNW PLVT11LL_CKT W=210.0n L=40.00n
XX4 net0139 B1 net0143 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX5 ZN B2 net0139 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX0 net0147 a1n VDD VNW PLVT11LL_CKT W=455.0n L=40.00n
XXP1 net0143 a2n net0147 VNW PLVT11LL_CKT W=455.0n L=40.00n
.ENDS LVT_I2NOR4HSV1
****Sub-Circuit for LVT_I2NOR4HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_I2NOR4HSV2 A1 A2 B1 B2 ZN VDD VSS
XX9 a2n A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX6 a1n A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 ZN B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN a1n VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 ZN B1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN a2n VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 a2n A2 VDD VNW PLVT11LL_CKT W=210.0n L=40.00n
XX7 a1n A1 VDD VNW PLVT11LL_CKT W=210.0n L=40.00n
XX4 net0139 B1 net0143 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX5 ZN B2 net0139 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX0 net0147 a1n VDD VNW PLVT11LL_CKT W=455.0n L=40.00n
XXP1 net0143 a2n net0147 VNW PLVT11LL_CKT W=455.0n L=40.00n
.ENDS LVT_I2NOR4HSV2
****Sub-Circuit for LVT_IAO21HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_IAO21HSV1 A1 A2 B ZN VDD VSS
XX3 net24 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 net24 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 ZN B VSS VPW NLVT11LL_CKT W=210.0n L=40.00n
XXN1 ZN net24 VSS VPW NLVT11LL_CKT W=210.0n L=40.00n
XX4 net24 A1 net056 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net056 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN net24 net064 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net064 B VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_IAO21HSV1
****Sub-Circuit for LVT_IAO21HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_IAO21HSV2 A1 A2 B ZN VDD VSS
XX3 net24 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 net24 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 ZN B VSS VPW NLVT11LL_CKT W=310.0n L=40.00n
XXN1 ZN net24 VSS VPW NLVT11LL_CKT W=310.0n L=40.00n
XX4 net24 A1 net056 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net056 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN net24 net064 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net064 B VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_IAO21HSV2
****Sub-Circuit for LVT_IAO22HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_IAO22HSV1 A1 A2 B1 B2 ZN VDD VSS
XX3 net24 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 net24 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 ZN B1 net050 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net050 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN net24 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 net061 B2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net24 A1 net074 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net074 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN net24 net061 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net061 B1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_IAO22HSV1
****Sub-Circuit for LVT_IAO22HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_IAO22HSV2 A1 A2 B1 B2 ZN VDD VSS
XX3 net24 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 net24 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 ZN B1 net050 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net050 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN net24 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 net061 B2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net24 A1 net074 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net074 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN net24 net061 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net061 B1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_IAO22HSV2
****Sub-Circuit for LVT_INAND2HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INAND2HSV1 A1 B1 ZN VDD VSS
XX3 net021 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 ZN net021 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 B1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 net021 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX0 ZN B1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN net021 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_INAND2HSV1
****Sub-Circuit for LVT_INAND2HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INAND2HSV2 A1 B1 ZN VDD VSS
XX3 net021 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 ZN net021 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 B1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 net021 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX0 ZN B1 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XXP1 ZN net021 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
.ENDS LVT_INAND2HSV2
****Sub-Circuit for LVT_INAND3HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INAND3HSV1 A1 B1 B2 ZN VDD VSS
XX5 net029 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net021 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 ZN net021 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 B1 net029 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 ZN B2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 net021 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX0 ZN B1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN net021 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_INAND3HSV1
****Sub-Circuit for LVT_INAND3HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INAND3HSV2 A1 B1 B2 ZN VDD VSS
XX5 net029 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net021 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 ZN net021 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 B1 net029 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 ZN B2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net021 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX0 ZN B1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN net021 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_INAND3HSV2
****Sub-Circuit for LVT_INAND4HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INAND4HSV1 A1 B1 B2 B3 ZN VDD VSS
XX8 net040 B3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX5 net029 B2 net040 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net021 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 ZN net021 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 B1 net029 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 ZN B3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX6 ZN B2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 net021 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX0 ZN B1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN net021 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_INAND4HSV1
****Sub-Circuit for LVT_INAND4HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INAND4HSV2 A1 B1 B2 B3 ZN VDD VSS
XX8 net040 B3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX5 net029 B2 net040 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net021 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 ZN net021 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 B1 net029 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 ZN B3 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX6 ZN B2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX4 net021 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX0 ZN B1 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XXP1 ZN net021 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
.ENDS LVT_INAND4HSV2
****Sub-Circuit for LVT_INHSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV1 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=310.0n L=40.00n
.ENDS LVT_INHSV1
****Sub-Circuit for LVT_INHSV12, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV12 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=1.4u L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=2.73u L=40.00n
.ENDS LVT_INHSV12
****Sub-Circuit for LVT_INHSV16, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV16 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=2.48u L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=3.64u L=40.00n
.ENDS LVT_INHSV16
****Sub-Circuit for LVT_INHSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV2 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=455.0n L=40.00n
.ENDS LVT_INHSV2
****Sub-Circuit for LVT_INHSV20, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV20 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=3.1u L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=4.55u L=40.00n
.ENDS LVT_INHSV20
****Sub-Circuit for LVT_INHSV24, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV24 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=3.72u L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=5.46u L=40.00n
.ENDS LVT_INHSV24
****Sub-Circuit for LVT_INHSV3, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV3 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=700.0n L=40.00n
.ENDS LVT_INHSV3
****Sub-Circuit for LVT_INHSV4, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV4 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=620.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=910.0n L=40.00n
.ENDS LVT_INHSV4
****Sub-Circuit for LVT_INHSV6, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV6 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=930.00n L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=1.365u L=40.00n
.ENDS LVT_INHSV6
****Sub-Circuit for LVT_INHSV8, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INHSV8 I ZN VDD VSS
XXN1 ZN I VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XXP1 ZN I VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
.ENDS LVT_INHSV8
****Sub-Circuit for LVT_INOR2HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INOR2HSV1 A1 B1 ZN VDD VSS
XX2 net27 A1 VSS VPW NLVT11LL_CKT W=140.0n L=40.00n
XX0 ZN B1 VSS VPW NLVT11LL_CKT W=285.0n L=40.00n
XXN1 ZN net27 VSS VPW NLVT11LL_CKT W=285.0n L=40.00n
XX1 ZN net27 net42 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX3 net27 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net42 B1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_INOR2HSV1
****Sub-Circuit for LVT_INOR2HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INOR2HSV2 A1 B1 ZN VDD VSS
XX2 net27 A1 VSS VPW NLVT11LL_CKT W=140.0n L=40.00n
XX0 ZN B1 VSS VPW NLVT11LL_CKT W=285.0n L=40.00n
XXN1 ZN net27 VSS VPW NLVT11LL_CKT W=285.0n L=40.00n
XX1 ZN net27 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX3 net27 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net42 B1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_INOR2HSV2
****Sub-Circuit for LVT_INOR3HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INOR3HSV1 A1 B1 B2 ZN VDD VSS
XX5 ZN net27 VSS VPW NLVT11LL_CKT W=210.0n L=40.00n
XX2 net27 A1 VSS VPW NLVT11LL_CKT W=140.0n L=40.00n
XX0 ZN B1 VSS VPW NLVT11LL_CKT W=210.0n L=40.00n
XXN1 ZN B2 VSS VPW NLVT11LL_CKT W=210.0n L=40.00n
XX4 net061 B2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 ZN net27 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX3 net27 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net42 B1 net061 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_INOR3HSV1
****Sub-Circuit for LVT_INOR3HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INOR3HSV2 A1 B1 B2 ZN VDD VSS
XX5 ZN net27 VSS VPW NLVT11LL_CKT W=310.0n L=40.00n
XX2 net27 A1 VSS VPW NLVT11LL_CKT W=140.0n L=40.00n
XX0 ZN B1 VSS VPW NLVT11LL_CKT W=310.0n L=40.00n
XXN1 ZN B2 VSS VPW NLVT11LL_CKT W=310.0n L=40.00n
XX4 net061 B2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 ZN net27 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX3 net27 A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 net42 B1 net061 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_INOR3HSV2
****Sub-Circuit for LVT_INOR4HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INOR4HSV1 A1 B1 B2 B3 ZN VDD VSS
XX7 ZN B3 VSS VPW NLVT11LL_CKT W=210.0n L=40.00n
XX5 ZN net27 VSS VPW NLVT11LL_CKT W=210.0n L=40.00n
XX2 net27 A1 VSS VPW NLVT11LL_CKT W=140.0n L=40.00n
XX0 ZN B1 VSS VPW NLVT11LL_CKT W=210.0n L=40.00n
XXN1 ZN B2 VSS VPW NLVT11LL_CKT W=210.0n L=40.00n
XX4 net061 B2 net070 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX6 net070 B3 VDD VNW PLVT11LL_CKT W=455.0n L=40.00n
XX1 ZN net27 net42 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX3 net27 A1 VDD VNW PLVT11LL_CKT W=210.0n L=40.00n
XXP1 net42 B1 net061 VNW PLVT11LL_CKT W=455.0n L=40.00n
.ENDS LVT_INOR4HSV1
****Sub-Circuit for LVT_INOR4HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_INOR4HSV2 A1 B1 B2 B3 ZN VDD VSS
XX7 ZN B3 VSS VPW NLVT11LL_CKT W=310.0n L=40.00n
XX5 ZN net27 VSS VPW NLVT11LL_CKT W=310.0n L=40.00n
XX2 net27 A1 VSS VPW NLVT11LL_CKT W=140.0n L=40.00n
XX0 ZN B1 VSS VPW NLVT11LL_CKT W=310.0n L=40.00n
XXN1 ZN B2 VSS VPW NLVT11LL_CKT W=310.0n L=40.00n
XX4 net061 B2 net070 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX6 net070 B3 VDD VNW PLVT11LL_CKT W=455.0n L=40.00n
XX1 ZN net27 net42 VNW PLVT11LL_CKT W=455.0n L=40.00n
XX3 net27 A1 VDD VNW PLVT11LL_CKT W=210.0n L=40.00n
XXP1 net42 B1 net061 VNW PLVT11LL_CKT W=455.0n L=40.00n
.ENDS LVT_INOR4HSV2
****Sub-Circuit for LVT_IOA21HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_IOA21HSV1 A1 A2 B ZN VDD VSS
XX2 ZN net038 net030 VPW NLVT11LL_CKT W=310n L=40.00n
XX3 net030 B VSS VPW NLVT11LL_CKT W=310n L=40.00n
XX1 net038 A1 net18 VPW NLVT11LL_CKT W=280n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=280n L=40.00n
XX4 ZN B VDD VNW PLVT11LL_CKT W=310n L=40.00n
XX5 ZN net038 VDD VNW PLVT11LL_CKT W=310n L=40.00n
XX0 net038 A2 VDD VNW PLVT11LL_CKT W=210n L=40.00n
XXP1 net038 A1 VDD VNW PLVT11LL_CKT W=210n L=40.00n
.ENDS LVT_IOA21HSV1
****Sub-Circuit for LVT_IOA21HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_IOA21HSV2 A1 A2 B ZN VDD VSS
XX2 ZN net038 net030 VPW NLVT11LL_CKT W=310n L=40.00n
XX3 net030 B VSS VPW NLVT11LL_CKT W=310n L=40.00n
XX1 net038 A1 net18 VPW NLVT11LL_CKT W=280n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=280n L=40.00n
XX4 ZN B VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 ZN net038 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net038 A2 VDD VNW PLVT11LL_CKT W=210n L=40.00n
XXP1 net038 A1 VDD VNW PLVT11LL_CKT W=210n L=40.00n
.ENDS LVT_IOA21HSV2
****Sub-Circuit for LVT_IOA22HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_IOA22HSV1 A1 A2 B1 B2 ZN VDD VSS
XX6 net030 B2 VSS VPW NLVT11LL_CKT W=310n L=40.00n
XX2 ZN net038 net030 VPW NLVT11LL_CKT W=310n L=40.00n
XX3 net030 B1 VSS VPW NLVT11LL_CKT W=310n L=40.00n
XX1 net038 A1 net18 VPW NLVT11LL_CKT W=280n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=280n L=40.00n
XX4 ZN B1 net063 VNW PLVT11LL_CKT W=430n L=40.00n
XX5 ZN net038 VDD VNW PLVT11LL_CKT W=310n L=40.00n
XX7 net063 B2 VDD VNW PLVT11LL_CKT W=430n L=40.00n
XX0 net038 A2 VDD VNW PLVT11LL_CKT W=210n L=40.00n
XXP1 net038 A1 VDD VNW PLVT11LL_CKT W=210n L=40.00n
.ENDS LVT_IOA22HSV1
****Sub-Circuit for LVT_IOA22HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_IOA22HSV2 A1 A2 B1 B2 ZN VDD VSS
XX6 net030 B2 VSS VPW NLVT11LL_CKT W=310n L=40.00n
XX2 ZN net038 net030 VPW NLVT11LL_CKT W=310n L=40.00n
XX3 net030 B1 VSS VPW NLVT11LL_CKT W=310n L=40.00n
XX1 net038 A1 net18 VPW NLVT11LL_CKT W=280n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=280n L=40.00n
XX4 ZN B1 net063 VNW PLVT11LL_CKT W=430n L=40.00n
XX5 ZN net038 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX7 net063 B2 VDD VNW PLVT11LL_CKT W=430n L=40.00n
XX0 net038 A2 VDD VNW PLVT11LL_CKT W=210n L=40.00n
XXP1 net038 A1 VDD VNW PLVT11LL_CKT W=210n L=40.00n
.ENDS LVT_IOA22HSV2
****Sub-Circuit for LVT_LALHSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_LALHSV1 D EN Q QN VDD VSS
XX46 Q net0104 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX30 cn c VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX27 c EN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX19 QN net_0154 VSS VPW NLVT11LL_CKT W=210n L=40.00n
XX12 net52 cn net0104 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 VSS net_0154 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net0104 c net69 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX7 net69 D VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX0 net_0154 net0104 VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX4 net128 D VDD VNW PLVT11LL_CKT W=400n L=40.00n
XX29 cn c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX28 c EN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX20 QN net_0154 VDD VNW PLVT11LL_CKT W=310n L=40.00n
XX47 Q net0104 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX14 net117 c net0104 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 VDD net_0154 net117 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX10 net0104 cn net128 VNW PLVT11LL_CKT W=400n L=40.00n
XX1 net_0154 net0104 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
.ENDS LVT_LALHSV1
****Sub-Circuit for LVT_LALHSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_LALHSV2 D EN Q QN VDD VSS
XX46 Q net0104 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX30 cn c VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX27 c EN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX19 QN net_0154 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 net52 cn net0104 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 VSS net_0154 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net0104 c net69 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX7 net69 D VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX0 net_0154 net0104 VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX4 net128 D VDD VNW PLVT11LL_CKT W=400n L=40.00n
XX29 cn c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX28 c EN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX20 QN net_0154 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX47 Q net0104 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX14 net117 c net0104 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 VDD net_0154 net117 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX10 net0104 cn net128 VNW PLVT11LL_CKT W=400n L=40.00n
XX1 net_0154 net0104 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
.ENDS LVT_LALHSV2
****Sub-Circuit for LVT_LALRNHSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_LALRNHSV1 D EN Q QN RDN VDD VSS
XX46 Q pm VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX44 net_0104 RDN VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX42 VSS RDN net_0119 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX30 cn c VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX27 c EN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX19 QN net_0154 VSS VPW NLVT11LL_CKT W=210n L=40.00n
XX12 net52 cn pm VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net_0119 net_0154 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 pm c net69 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX7 net69 D net_0104 VPW NLVT11LL_CKT W=285.00n L=40.00n
XX0 net_0154 pm VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX43 pm RDN VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX29 cn c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX28 c EN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX20 QN net_0154 VDD VNW PLVT11LL_CKT W=310n L=40.00n
XX47 Q pm VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX14 net117 c pm VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 VDD net_0154 net117 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX10 pm cn net128 VNW PLVT11LL_CKT W=400n L=40.00n
XX8 net128 D VDD VNW PLVT11LL_CKT W=400n L=40.00n
XX1 net_0154 pm VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
.ENDS LVT_LALRNHSV1
****Sub-Circuit for LVT_LALRNHSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_LALRNHSV2 D EN Q QN RDN VDD VSS
XX46 Q pm VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX44 net_0104 RDN VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX42 VSS RDN net_0119 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX30 cn c VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX27 c EN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX19 QN net_0154 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 net52 cn pm VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net_0119 net_0154 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 pm c net69 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX7 net69 D net_0104 VPW NLVT11LL_CKT W=285.00n L=40.00n
XX0 net_0154 pm VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX43 pm RDN VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX29 cn c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX28 c EN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX20 QN net_0154 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX47 Q pm VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX14 net117 c pm VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 VDD net_0154 net117 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX10 pm cn net128 VNW PLVT11LL_CKT W=400n L=40.00n
XX8 net128 D VDD VNW PLVT11LL_CKT W=400n L=40.00n
XX1 net_0154 pm VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
.ENDS LVT_LALRNHSV2
****Sub-Circuit for LVT_LALRSNHSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_LALRSNHSV1 D EN Q QN RDN SDN VDD VSS
XX2 m SDN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX6 net0156 RDN VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX46 Q net0152 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX21 net0152 m VSS VPW NLVT11LL_CKT W=170.00n L=40.00n
XX42 VSS RDN net_0119 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX30 cn c VSS VPW NLVT11LL_CKT W=315.00n L=40.00n
XX27 c EN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX19 QN net_0154 VSS VPW NLVT11LL_CKT W=210n L=40.00n
XX12 net52 cn net0152 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net_0119 net_0154 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net0152 c net69 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX7 net69 D net0156 VPW NLVT11LL_CKT W=285.00n L=40.00n
XX0 net_0154 net0152 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX3 m SDN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX18 net0152 RDN net0267 VNW PLVT11LL_CKT W=205.00n L=40.00n
XX4 net0267 m VDD VNW PLVT11LL_CKT W=205.00n L=40.00n
XX17 net0272 net_0154 net117 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX16 net128 D net0251 VNW PLVT11LL_CKT W=400n L=40.00n
XX29 cn c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX28 c EN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX20 QN net_0154 VDD VNW PLVT11LL_CKT W=310n L=40.00n
XX47 Q net0152 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX14 net117 c net0152 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 VDD m net0272 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX10 net0152 cn net128 VNW PLVT11LL_CKT W=400n L=40.00n
XX8 net0251 m VDD VNW PLVT11LL_CKT W=400n L=40.00n
XX1 net_0154 net0152 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
.ENDS LVT_LALRSNHSV1
****Sub-Circuit for LVT_LALRSNHSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_LALRSNHSV2 D EN Q QN RDN SDN VDD VSS
XX2 m SDN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX6 net0156 RDN VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX46 Q net0152 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX21 net0152 m VSS VPW NLVT11LL_CKT W=170.00n L=40.00n
XX42 VSS RDN net_0119 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX30 cn c VSS VPW NLVT11LL_CKT W=315.00n L=40.00n
XX27 c EN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX19 QN net_0154 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 net52 cn net0152 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net_0119 net_0154 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net0152 c net69 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX7 net69 D net0156 VPW NLVT11LL_CKT W=285.00n L=40.00n
XX0 net_0154 net0152 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX3 m SDN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX18 net0152 RDN net0267 VNW PLVT11LL_CKT W=205.00n L=40.00n
XX4 net0267 m VDD VNW PLVT11LL_CKT W=205.00n L=40.00n
XX17 net0272 net_0154 net117 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX16 net128 D net0251 VNW PLVT11LL_CKT W=400n L=40.00n
XX29 cn c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX28 c EN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX20 QN net_0154 VDD VNW PLVT11LL_CKT W=445.00n L=40.00n
XX47 Q net0152 VDD VNW PLVT11LL_CKT W=445.00n L=40.00n
XX14 net117 c net0152 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 VDD m net0272 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX10 net0152 cn net128 VNW PLVT11LL_CKT W=400n L=40.00n
XX8 net0251 m VDD VNW PLVT11LL_CKT W=400n L=40.00n
XX1 net_0154 net0152 VDD VNW PLVT11LL_CKT W=355.00n L=40.00n
.ENDS LVT_LALRSNHSV2
****Sub-Circuit for LVT_LALSNHSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_LALSNHSV1 D EN Q QN SDN VDD VSS
XX2 rn SDN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX46 Q net0129 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX44 net0129 rn VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX30 cn c VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX27 c EN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX19 QN net_0154 VSS VPW NLVT11LL_CKT W=210n L=40.00n
XX12 net52 cn net0129 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 VSS net_0154 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net0129 c net69 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX7 net69 D VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX0 net_0154 net0129 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX3 rn SDN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX4 net128 D net0143 VNW PLVT11LL_CKT W=400n L=40.00n
XX5 VDD rn net0189 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX29 cn c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX28 c EN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX20 QN net_0154 VDD VNW PLVT11LL_CKT W=310n L=40.00n
XX47 Q net0129 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX14 net117 c net0129 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 net0189 net_0154 net117 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX10 net0129 cn net128 VNW PLVT11LL_CKT W=400n L=40.00n
XX8 net0143 rn VDD VNW PLVT11LL_CKT W=400n L=40.00n
XX1 net_0154 net0129 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
.ENDS LVT_LALSNHSV1
****Sub-Circuit for LVT_LALSNHSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_LALSNHSV2 D EN Q QN SDN VDD VSS
XX46 Q net0119 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net0119 rn VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX3 rn SDN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX30 cn c VSS VPW NLVT11LL_CKT W=320.00n L=40.00n
XX27 c EN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX19 QN net_0154 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 net52 cn net0119 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 VSS net_0154 net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX9 net0119 c net69 VPW NLVT11LL_CKT W=190.00n L=40.00n
XX7 net69 D VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX0 net_0154 net0119 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX4 rn SDN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX5 net0171 rn VDD VNW PLVT11LL_CKT W=400n L=40.00n
XX6 VDD rn net0144 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX29 cn c VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX28 c EN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX20 QN net_0154 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX47 Q net0119 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX14 net117 c net0119 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 net0144 net_0154 net117 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX10 net0119 cn net128 VNW PLVT11LL_CKT W=400n L=40.00n
XX8 net128 D net0171 VNW PLVT11LL_CKT W=400n L=40.00n
XX1 net_0154 net0119 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
.ENDS LVT_LALSNHSV2
****Sub-Circuit for LVT_MAOI222HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MAOI222HSV1 A B C ZN VDD VSS
XX6 ZN B net4 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX10 net4 C VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 net5 B VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN C net6 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN A net5 VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net6 A VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 net2 C net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX11 ZN A net2 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX7 net1 C VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net1 A VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net2 B net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN B net2 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_MAOI222HSV1
****Sub-Circuit for LVT_MAOI222HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MAOI222HSV2 A B C ZN VDD VSS
XX6 ZN B net4 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX10 net4 C VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 net5 B VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN C net6 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN A net5 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net6 A VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 net2 C net1 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX11 ZN A net2 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX7 net1 C VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net1 A VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net2 B net1 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN B net2 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_MAOI222HSV2
****Sub-Circuit for LVT_MAOI22HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MAOI22HSV1 A1 A2 B1 B2 ZN VDD VSS
XX2 net039 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 ZN A2 net039 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 ZN net5 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 net5 B1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XXN1 net5 B2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 net063 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 ZN net5 net063 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX7 net1 B2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net063 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net5 B1 net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_MAOI22HSV1
****Sub-Circuit for LVT_MAOI22HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MAOI22HSV2 A1 A2 B1 B2 ZN VDD VSS
XX2 net039 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 ZN A2 net039 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 ZN net5 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 net5 B1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XXN1 net5 B2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 net063 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 ZN net5 net063 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX7 net1 B2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net063 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net5 B1 net1 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_MAOI22HSV2
****Sub-Circuit for LVT_MOAI22HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MOAI22HSV1 A1 A2 B1 B2 ZN VDD VSS
XX2 net039 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 ZN net1 net039 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 net039 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX10 net1 B1 net055 VPW NLVT11LL_CKT W=280.00n L=40.00n
XX9 net055 B2 VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX1 net063 A2 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX4 ZN A1 net063 VNW PLVT11LL_CKT W=430.00n L=40.00n
XX8 net1 B2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX11 ZN net1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX7 net1 B1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_MOAI22HSV1
****Sub-Circuit for LVT_MOAI22HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MOAI22HSV2 A1 A2 B1 B2 ZN VDD VSS
XX2 net039 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 ZN net1 net039 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 net039 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX10 net1 B1 net055 VPW NLVT11LL_CKT W=280.00n L=40.00n
XX9 net055 B2 VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX1 net063 A2 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX4 ZN A1 net063 VNW PLVT11LL_CKT W=430.00n L=40.00n
XX8 net1 B2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX11 ZN net1 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX7 net1 B1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_MOAI22HSV2
****Sub-Circuit for LVT_MUX2HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX2HSV1 I0 I1 S Z VDD VSS
XX47 net41 S net64 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX51 Z net64 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 net39 I0 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX31 net41 I1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX53 net43 S VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 net39 net43 net64 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 net39 I0 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX52 Z net64 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX48 net41 net43 net64 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX32 net41 I1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 net43 S VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX39 net39 S net64 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_MUX2HSV1
****Sub-Circuit for LVT_MUX2HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX2HSV2 I0 I1 S Z VDD VSS
XX47 net41 S net64 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX51 Z net64 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX49 net39 I0 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX31 net41 I1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX53 net43 S VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 net39 net43 net64 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 net39 I0 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX52 Z net64 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX48 net41 net43 net64 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX32 net41 I1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 net43 S VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX39 net39 S net64 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_MUX2HSV2
****Sub-Circuit for LVT_MUX2NHSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX2NHSV1 I0 I1 S ZN VDD VSS
XX47 net41 S ZN VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 net39 I0 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX31 net41 I1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX53 net43 S VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 net39 net43 ZN VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 net39 I0 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX48 net41 net43 ZN VNW PLVT11LL_CKT W=310.00n L=40.00n
XX32 net41 I1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 net43 S VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX39 net39 S ZN VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_MUX2NHSV1
****Sub-Circuit for LVT_MUX2NHSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX2NHSV2 I0 I1 S ZN VDD VSS
XX47 net41 S ZN VPW NLVT11LL_CKT W=310.00n L=40.00n
XX49 net39 I0 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX31 net41 I1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX53 net43 S VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 net39 net43 ZN VPW NLVT11LL_CKT W=310.00n L=40.00n
XX50 net39 I0 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX48 net41 net43 ZN VNW PLVT11LL_CKT W=365.00n L=40.00n
XX32 net41 I1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 net43 S VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX39 net39 S ZN VNW PLVT11LL_CKT W=365.00n L=40.00n
.ENDS LVT_MUX2NHSV2
****Sub-Circuit for LVT_MUX3HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX3HSV1 I0 I1 I2 S0 S1 Z VDD VSS
XX3 net_0205 I0 net_57 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net_57 sn VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX24 Z net_0201 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 net_0205 I1 net_77 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net_77 S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net0116 S1 net_0189 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX14 net0116 net_0205 net_0197 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net_0189 in VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX15 net_0197 s1n VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 s1n S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX26 net_0201 net0116 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX53 sn S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX22 in I2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX27 net_0201 net0116 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX23 in I2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX25 Z net_0201 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net_0205 S0 net_108 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net_108 sn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net_108 I0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net_0205 I1 net_108 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX13 s1n S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 net0116 in net_0268 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX54 sn S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX21 net0116 S1 net_0268 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX20 net_0268 s1n VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net_0268 net_0205 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_MUX3HSV1
****Sub-Circuit for LVT_MUX3HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX3HSV2 I0 I1 I2 S0 S1 Z VDD VSS
XX3 net_0205 I0 net_57 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net_57 sn VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX24 Z net_0201 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 net_0205 I1 net_77 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net_77 S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net0116 S1 net_0189 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX14 net0116 net_0205 net_0197 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net_0189 in VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX15 net_0197 s1n VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 s1n S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX26 net_0201 net0116 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX53 sn S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX22 in I2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX27 net_0201 net0116 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX23 in I2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX25 Z net_0201 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net_0205 S0 net_108 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net_108 sn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net_108 I0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net_0205 I1 net_108 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX13 s1n S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 net0116 in net_0268 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX54 sn S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX21 net0116 S1 net_0268 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX20 net_0268 s1n VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net_0268 net_0205 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_MUX3HSV2
****Sub-Circuit for LVT_MUX3NHSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX3NHSV1 I0 I1 I2 S0 S1 ZN VDD VSS
XX3 net_0205 I0 net_57 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net_57 sn VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX24 ZN net_0201 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 net_0205 I1 net_77 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net_77 S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net_0201 S1 net_0189 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX14 net_0201 net_0205 net_0197 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net_0189 in VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX15 net_0197 s1n VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 s1n S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX53 sn S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX22 in I2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX23 in I2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX25 ZN net_0201 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net_0205 S0 net_108 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net_108 sn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net_108 I0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net_0205 I1 net_108 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX13 s1n S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 net_0201 in net_0268 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX54 sn S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX21 net_0201 S1 net_0268 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX20 net_0268 s1n VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net_0268 net_0205 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_MUX3NHSV1
****Sub-Circuit for LVT_MUX3NHSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX3NHSV2 I0 I1 I2 S0 S1 ZN VDD VSS
XX3 net_0205 I0 net_57 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net_57 sn VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX24 ZN net_0201 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 net_0205 I1 net_77 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net_77 S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 net_0201 S1 net_0189 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX14 net_0201 net_0205 net_0197 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net_0189 in VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX15 net_0197 s1n VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 s1n S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX53 sn S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX22 in I2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX23 in I2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX25 ZN net_0201 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net_0205 S0 net_108 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net_108 sn VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net_108 I0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net_0205 I1 net_108 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX13 s1n S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 net_0201 in net_0268 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX54 sn S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX21 net_0201 S1 net_0268 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX20 net_0268 s1n VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net_0268 net_0205 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_MUX3NHSV2
****Sub-Circuit for LVT_MUX4HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX4HSV1 I0 I1 I2 I3 S0 S1 Z VDD VSS
XX28 net164 I3 net160 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX29 net160 S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX30 net164 s1n net152 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX31 net152 I1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net168 S0 net172 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net172 net164 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 net168 m net180 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net180 sn VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 m I0 net136 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX14 m I2 net140 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net136 s1n VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX15 net140 S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 s1n S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX38 Z net148 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 net148 net168 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX53 sn S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX32 net164 I1 net235 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX33 net235 I3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX34 net235 S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX35 net164 s1n net235 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net168 sn net239 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net239 net164 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX37 net148 net168 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net239 S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net168 m net239 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX13 s1n S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 m s1n net199 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX54 sn S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX39 Z net148 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX21 m I0 net199 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX20 net199 I2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net199 S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_MUX4HSV1
****Sub-Circuit for LVT_MUX4HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX4HSV2 I0 I1 I2 I3 S0 S1 Z VDD VSS
XX28 net164 I3 net160 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX29 net160 S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX30 net164 s1n net152 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX31 net152 I1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net168 S0 net172 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net172 net164 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 net168 m net180 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net180 sn VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 m I0 net136 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX14 m I2 net140 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net136 s1n VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX15 net140 S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 s1n S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX38 Z net148 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX36 net148 net168 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX53 sn S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX32 net164 I1 net235 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX33 net235 I3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX34 net235 S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX35 net164 s1n net235 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net168 sn net239 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net239 net164 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX37 net148 net168 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net239 S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net168 m net239 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX13 s1n S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 m s1n net199 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX54 sn S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX39 Z net148 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX21 m I0 net199 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX20 net199 I2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net199 S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_MUX4HSV2
****Sub-Circuit for LVT_MUX4NHSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX4NHSV1 I0 I1 I2 I3 S0 S1 ZN VDD VSS
XX28 net164 I3 net160 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX29 net160 S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX30 net164 s1n net152 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX31 net152 I1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net168 S0 net172 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net172 net164 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 net168 m net180 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net180 sn VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 m I0 net136 VPW NLVT11LL_CKT W=290.00n L=40.00n
XX14 m I2 net140 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net136 s1n VSS VPW NLVT11LL_CKT W=290.00n L=40.00n
XX15 net140 S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 s1n S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX38 ZN net168 VSS VPW NLVT11LL_CKT W=215.00n L=40.00n
XX53 sn S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX32 net164 I1 net235 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX33 net235 I3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX34 net235 S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX35 net164 s1n net235 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net168 sn net239 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net239 net164 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net239 S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net168 m net239 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX13 s1n S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 m s1n net199 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX54 sn S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX39 ZN net168 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX21 m I0 net199 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX20 net199 I2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net199 S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_MUX4NHSV1
****Sub-Circuit for LVT_MUX4NHSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_MUX4NHSV2 I0 I1 I2 I3 S0 S1 ZN VDD VSS
XX28 net164 I3 net160 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX29 net160 S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX30 net164 s1n net152 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX31 net152 I1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net168 S0 net172 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net172 net164 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX6 net168 m net180 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net180 sn VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 m I0 net136 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX14 m I2 net140 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net136 s1n VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX15 net140 S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 s1n S1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX38 ZN net168 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX53 sn S0 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX32 net164 I1 net235 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX33 net235 I3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX34 net235 S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX35 net164 s1n net235 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net168 sn net239 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net239 net164 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net239 S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 net168 m net239 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX13 s1n S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 m s1n net199 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX54 sn S0 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX39 ZN net168 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX21 m I0 net199 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX20 net199 I2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX19 net199 S1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_MUX4NHSV2
****Sub-Circuit for LVT_NAND2HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND2HSV1 A1 A2 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_NAND2HSV1
****Sub-Circuit for LVT_NAND2HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND2HSV2 A1 A2 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NAND2HSV2
****Sub-Circuit for LVT_NAND2HSV3, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND2HSV3 A1 A2 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=460.00n L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
.ENDS LVT_NAND2HSV3
****Sub-Circuit for LVT_NAND2HSV8, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND2HSV8 A1 A2 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=1.24u L=40.00n
XXN1 net18 A2 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
.ENDS LVT_NAND2HSV8
****Sub-Circuit for LVT_NAND3HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND3HSV1 A1 A2 A3 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net022 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net022 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 ZN A3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_NAND3HSV1
****Sub-Circuit for LVT_NAND3HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND3HSV2 A1 A2 A3 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net022 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net022 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 ZN A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NAND3HSV2
****Sub-Circuit for LVT_NAND3HSV3, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND3HSV3 A1 A2 A3 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=460.00n L=40.00n
XX3 net022 A3 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XXN1 net18 A2 net022 VPW NLVT11LL_CKT W=460.00n L=40.00n
XX2 ZN A3 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
.ENDS LVT_NAND3HSV3
****Sub-Circuit for LVT_NAND3HSV8, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND3HSV8 A1 A2 A3 ZN VDD VSS
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=1.24u L=40.00n
XX3 net022 A3 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XXN1 net18 A2 net022 VPW NLVT11LL_CKT W=1.24u L=40.00n
XX2 ZN A3 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
.ENDS LVT_NAND3HSV8
****Sub-Circuit for LVT_NAND4HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND4HSV1 A1 A2 A3 A4 ZN VDD VSS
XX4 net026 A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net022 A3 net026 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net022 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX5 ZN A4 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX2 ZN A3 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_NAND4HSV1
****Sub-Circuit for LVT_NAND4HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND4HSV2 A1 A2 A3 A4 ZN VDD VSS
XX4 net026 A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net022 A3 net026 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net022 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX5 ZN A4 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 ZN A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NAND4HSV2
****Sub-Circuit for LVT_NAND4HSV3, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND4HSV3 A1 A2 A3 A4 ZN VDD VSS
XX4 net026 A4 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=460.00n L=40.00n
XX3 net022 A3 net026 VPW NLVT11LL_CKT W=460.00n L=40.00n
XXN1 net18 A2 net022 VPW NLVT11LL_CKT W=460.00n L=40.00n
XX5 ZN A4 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
XX2 ZN A3 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
XX0 ZN A2 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
XXP1 ZN A1 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
.ENDS LVT_NAND4HSV3
****Sub-Circuit for LVT_NAND4HSV8, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NAND4HSV8 A1 A2 A3 A4 ZN VDD VSS
XX8 ZN net036 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX7 net036 net060 VSS VPW NLVT11LL_CKT W=620.00n L=40.00n
XX4 net026 A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net060 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net022 A3 net026 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net18 A2 net022 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 ZN net036 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX5 net060 A4 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net060 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX6 net036 net060 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
XX0 net060 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net060 A1 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NAND4HSV8
****Sub-Circuit for LVT_NOR2HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR2HSV1 A1 A2 ZN VDD VSS
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 net34 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net34 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NOR2HSV1
****Sub-Circuit for LVT_NOR2HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR2HSV2 A1 A2 ZN VDD VSS
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net34 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net34 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NOR2HSV2
****Sub-Circuit for LVT_NOR2HSV3, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR2HSV3 A1 A2 ZN VDD VSS
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX1 ZN A1 net34 VNW PLVT11LL_CKT W=700.00n L=40.00n
XXP1 net34 A2 VDD VNW PLVT11LL_CKT W=700.00n L=40.00n
.ENDS LVT_NOR2HSV3
****Sub-Circuit for LVT_NOR2HSV8, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR2HSV8 A1 A2 ZN VDD VSS
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=1.2u L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=1.2u L=40.00n
XX1 ZN A1 net34 VNW PLVT11LL_CKT W=1.8u L=40.00n
XXP1 net34 A2 VDD VNW PLVT11LL_CKT W=1.8u L=40.00n
.ENDS LVT_NOR2HSV8
****Sub-Circuit for LVT_NOR3HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR3HSV1 A1 A2 A3 ZN VDD VSS
XX3 ZN A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 net47 A3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net43 VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 net43 A2 net47 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_NOR3HSV1
****Sub-Circuit for LVT_NOR3HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR3HSV2 A1 A2 A3 ZN VDD VSS
XX3 ZN A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net47 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 ZN A1 net43 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net43 A2 net47 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NOR3HSV2
****Sub-Circuit for LVT_NOR3HSV3, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR3HSV3 A1 A2 A3 ZN VDD VSS
XX3 ZN A3 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX2 net47 A3 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
XX1 ZN A1 net43 VNW PLVT11LL_CKT W=680.00n L=40.00n
XXP1 net43 A2 net47 VNW PLVT11LL_CKT W=680.00n L=40.00n
.ENDS LVT_NOR3HSV3
****Sub-Circuit for LVT_NOR3HSV8, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR3HSV8 A1 A2 A3 ZN VDD VSS
XX3 ZN A3 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX2 net47 A3 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX1 ZN A1 net43 VNW PLVT11LL_CKT W=1.82u L=40.00n
XXP1 net43 A2 net47 VNW PLVT11LL_CKT W=1.82u L=40.00n
.ENDS LVT_NOR3HSV8
****Sub-Circuit for LVT_NOR4HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR4HSV1 A1 A2 A3 A4 ZN VDD VSS
XX4 ZN A4 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX3 ZN A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX5 net047 A4 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net47 A3 net047 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 ZN A1 net43 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net43 A2 net47 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NOR4HSV1
****Sub-Circuit for LVT_NOR4HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR4HSV2 A1 A2 A3 A4 ZN VDD VSS
XX4 ZN A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 ZN A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX5 net047 A4 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net47 A3 net047 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 ZN A1 net43 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net43 A2 net47 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NOR4HSV2
****Sub-Circuit for LVT_NOR4HSV3, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR4HSV3 A1 A2 A3 A4 ZN VDD VSS
XX4 ZN A4 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX3 ZN A3 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX0 ZN A2 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XXN1 ZN A1 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX5 net047 A4 VDD VNW PLVT11LL_CKT W=680.00n L=40.00n
XX2 net47 A3 net047 VNW PLVT11LL_CKT W=680.00n L=40.00n
XX1 ZN A1 net43 VNW PLVT11LL_CKT W=680.00n L=40.00n
XXP1 net43 A2 net47 VNW PLVT11LL_CKT W=680.00n L=40.00n
.ENDS LVT_NOR4HSV3
****Sub-Circuit for LVT_NOR4HSV8, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_NOR4HSV8 A1 A2 A3 A4 ZN VDD VSS
XX7 net033 net049 VSS VPW NLVT11LL_CKT W=620.00n L=40.00n
XX8 ZN net033 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XX4 net049 A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net049 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX0 net049 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net049 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 ZN net033 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX5 net047 A4 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX2 net47 A3 net047 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net049 A1 net43 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX6 net033 net049 VDD VNW PLVT11LL_CKT W=910.00n L=40.00n
XXP1 net43 A2 net47 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_NOR4HSV8
****Sub-Circuit for LVT_OAI211HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI211HSV1 A1 A2 B C ZN VDD VSS
XX2 ZN B net030 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX3 net030 C net027 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 net027 A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net027 A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN B VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 ZN C VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_OAI211HSV1
****Sub-Circuit for LVT_OAI211HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI211HSV2 A1 A2 B C ZN VDD VSS
XX2 ZN B net030 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net030 C net027 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net027 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net027 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 ZN C VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OAI211HSV2
****Sub-Circuit for LVT_OAI21HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI21HSV1 A1 A2 B ZN VDD VSS
XX2 ZN B net029 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 net029 A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net029 A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN B VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_OAI21HSV1
****Sub-Circuit for LVT_OAI21HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI21HSV2 A1 A2 B ZN VDD VSS
XX2 ZN B net029 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net029 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net029 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OAI21HSV2
****Sub-Circuit for LVT_OAI221HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI221HSV1 A1 A2 B1 B2 C ZN VDD VSS
XX9 net18 B2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 net18 B1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX3 ZN C net045 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 net045 A2 net18 VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net045 A1 net18 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 net071 B2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 ZN C VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_OAI221HSV1
****Sub-Circuit for LVT_OAI221HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI221HSV2 A1 A2 B1 B2 C ZN VDD VSS
XX9 net18 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net18 B1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 ZN C net045 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net045 A2 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net045 A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 net071 B2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 ZN C VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OAI221HSV2
****Sub-Circuit for LVT_OAI222HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI222HSV1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX12 net030 B2 VSS VPW NLVT11LL_CKT W=210n L=40.00n
XX9 net18 A2 net030 VPW NLVT11LL_CKT W=210n L=40.00n
XX2 net18 A1 net030 VPW NLVT11LL_CKT W=210n L=40.00n
XX3 net030 B1 VSS VPW NLVT11LL_CKT W=210n L=40.00n
XX1 ZN C1 net18 VPW NLVT11LL_CKT W=210n L=40.00n
XXN1 ZN C2 net18 VPW NLVT11LL_CKT W=210n L=40.00n
XX8 net071 B2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX10 net073 C2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX11 ZN C1 net073 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_OAI222HSV1
****Sub-Circuit for LVT_OAI222HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI222HSV2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
XX12 net030 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 net18 A2 net030 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net18 A1 net030 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net030 B1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN C1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN C2 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 net071 B2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX10 net073 C2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX11 ZN C1 net073 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OAI222HSV2
****Sub-Circuit for LVT_OAI22HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI22HSV1 A1 A2 B1 B2 ZN VDD VSS
XX9 net18 B2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 net18 B1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 ZN A2 net18 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 net071 B2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_OAI22HSV1
****Sub-Circuit for LVT_OAI22HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI22HSV2 A1 A2 B1 B2 ZN VDD VSS
XX9 net18 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net18 B1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN A2 net18 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX8 net071 B2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net067 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OAI22HSV2
****Sub-Circuit for LVT_OAI31HSV1, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI31HSV1 A1 A2 A3 B ZN VDD VSS
XX2 ZN B net064 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 net064 A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 net064 A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net064 A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN B VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX8 net065 A3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net067 A2 net065 VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_OAI31HSV1
****Sub-Circuit for LVT_OAI31HSV2, Wed Sep  5 13:54:27 CST 2012****
.SUBCKT LVT_OAI31HSV2 A1 A2 A3 B ZN VDD VSS
XX2 ZN B net064 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 net064 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net064 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net064 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net065 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net067 A2 net065 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OAI31HSV2
****Sub-Circuit for LVT_OAI32HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OAI32HSV1 A1 A2 A3 B1 B2 ZN VDD VSS
XX11 net041 B2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 net041 B1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 ZN A3 net041 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN A1 net041 VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 ZN A2 net041 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX8 net065 A3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX10 net071 B2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net067 A2 net065 VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_OAI32HSV1
****Sub-Circuit for LVT_OAI32HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OAI32HSV2 A1 A2 A3 B1 B2 ZN VDD VSS
XX11 net041 B2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net041 B1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 ZN A3 net041 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN A1 net041 VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN A2 net041 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net065 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX10 net071 B2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net067 A2 net065 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OAI32HSV2
****Sub-Circuit for LVT_OAI33HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OAI33HSV1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX11 net041 A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 net041 A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX9 ZN B3 net041 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 ZN B1 net041 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX13 net041 A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 ZN B2 net041 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX12 net076 B3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX8 net065 A3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX10 net071 B2 net076 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX0 net067 A2 net065 VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_OAI33HSV1
****Sub-Circuit for LVT_OAI33HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OAI33HSV2 A1 A2 A3 B1 B2 B3 ZN VDD VSS
XX11 net041 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 net041 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX9 ZN B3 net041 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 ZN B1 net041 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX13 net041 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 ZN B2 net041 VPW NLVT11LL_CKT W=310.00n L=40.00n
XX12 net076 B3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 ZN B1 net071 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net065 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX10 net071 B2 net076 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX0 net067 A2 net065 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 ZN A1 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OAI33HSV2
****Sub-Circuit for LVT_OR2HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OR2HSV1 A1 A2 Z VDD VSS
XX0 net31 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net31 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net31 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 net31 A1 net42 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX4 Z net31 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XXP1 net42 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_OR2HSV1
****Sub-Circuit for LVT_OR2HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OR2HSV2 A1 A2 Z VDD VSS
XX0 net31 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net31 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net31 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 net31 A1 net42 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX4 Z net31 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net42 A2 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_OR2HSV2
****Sub-Circuit for LVT_OR2HSV8, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OR2HSV8 A1 A2 Z VDD VSS
XX0 net31 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net31 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XXN1 net31 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net31 A1 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 Z net31 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XXP1 net42 A2 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OR2HSV8
****Sub-Circuit for LVT_OR3HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OR3HSV1 A1 A2 A3 Z VDD VSS
XX3 net31 A3 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 net31 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net31 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net31 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 net31 A1 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 Z net31 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net054 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net42 A2 net054 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OR3HSV1
****Sub-Circuit for LVT_OR3HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OR3HSV2 A1 A2 A3 Z VDD VSS
XX3 net31 A3 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 net31 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net31 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net31 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX1 net31 A1 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 Z net31 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net054 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net42 A2 net054 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OR3HSV2
****Sub-Circuit for LVT_OR3HSV8, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OR3HSV8 A1 A2 A3 Z VDD VSS
XX3 net31 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX0 net31 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net31 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XXN1 net31 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX1 net31 A1 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 Z net31 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX5 net054 A3 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net42 A2 net054 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OR3HSV8
****Sub-Circuit for LVT_OR4HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OR4HSV1 A1 A2 A3 A4 Z VDD VSS
XX6 net31 A4 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 net31 A3 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 net31 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net31 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXN1 net31 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX7 net067 A4 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net31 A1 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 Z net31 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net054 A3 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net42 A2 net054 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OR4HSV1
****Sub-Circuit for LVT_OR4HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OR4HSV2 A1 A2 A3 A4 Z VDD VSS
XX6 net31 A4 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 net31 A3 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 net31 A2 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 Z net31 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XXN1 net31 A1 VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX7 net067 A4 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net31 A1 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 Z net31 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX5 net054 A3 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net42 A2 net054 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OR4HSV2
****Sub-Circuit for LVT_OR4HSV8, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_OR4HSV8 A1 A2 A3 A4 Z VDD VSS
XX6 net31 A4 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX3 net31 A3 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX0 net31 A2 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 Z net31 VSS VPW NLVT11LL_CKT W=1.24u L=40.00n
XXN1 net31 A1 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX7 net067 A4 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX1 net31 A1 net42 VNW PLVT11LL_CKT W=455.00n L=40.00n
XX4 Z net31 VDD VNW PLVT11LL_CKT W=1.82u L=40.00n
XX5 net054 A3 net067 VNW PLVT11LL_CKT W=455.00n L=40.00n
XXP1 net42 A2 net054 VNW PLVT11LL_CKT W=455.00n L=40.00n
.ENDS LVT_OR4HSV8
****Sub-Circuit for LVT_PULLHS0, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_PULLHS0 Z VDD VSS
XXN1 Z net18 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XXP1 net18 net18 VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
.ENDS LVT_PULLHS0
****Sub-Circuit for LVT_PULLHS1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_PULLHS1 Z VDD VSS
XXN1 net14 net14 VSS VPW NLVT11LL_CKT W=140.0n L=40.00n
XXP1 Z net14 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_PULLHS1
****Sub-Circuit for LVT_SDHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDHSV1 CK D Q QN SE SI VDD VSS
XX13 VDD m net138 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=390.00n L=40.00n
XX10 QN ps VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX8 net174 SEN net177 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX44 net177 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX45 net177 SE VDD VNW PLVT11LL_CKT W=320.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX6 net174 D net177 VNW PLVT11LL_CKT W=320.00n L=40.00n
XX9 pm c net174 VNW PLVT11LL_CKT W=320.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net150 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net150 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net138 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX5 QN ps VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net202 D VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=300.00n L=40.00n
XX41 net258 SI net254 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net254 SE VSS VPW NLVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn net258 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=210.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net229 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net229 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX17 s ps VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net213 c pm VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS m net213 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX40 net258 SEN net202 VPW NLVT11LL_CKT W=140.00n L=40.00n
.ENDS LVT_SDHSV1
****Sub-Circuit for LVT_SDHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDHSV2 CK D Q QN SE SI VDD VSS
XX5 QN ps VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX41 net_0127 SI net_0123 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net_0123 SE VSS VPW NLVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn net_0127 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=210.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 s ps VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net52 c pm VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS m net52 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX40 net_0127 SEN net69 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX7 net69 D VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=300.00n L=40.00n
XX10 QN ps VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0226 SEN net_0202 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX44 net_0202 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0202 SE VDD VNW PLVT11LL_CKT W=320.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX6 net0226 D net_0202 VNW PLVT11LL_CKT W=320.00n L=40.00n
XX9 pm c net0226 VNW PLVT11LL_CKT W=320.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD m net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=390.00n L=40.00n
.ENDS LVT_SDHSV2
****Sub-Circuit for LVT_SDQHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDQHSV1 CK D Q SE SI VDD VSS
XX13 VDD m net128 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=345.00n L=40.00n
XX8 net164 SEN net167 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX44 net167 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX45 net167 SE VDD VNW PLVT11LL_CKT W=320.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX6 net164 D net167 VNW PLVT11LL_CKT W=320.00n L=40.00n
XX9 pm c net164 VNW PLVT11LL_CKT W=220.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net140 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net140 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net128 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX7 net188 D VSS VPW NLVT11LL_CKT W=160.00n L=40.00n
XX41 net244 SI net240 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net240 SE VSS VPW NLVT11LL_CKT W=120.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX2 pm cn net244 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=180.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net215 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net215 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX17 s ps VSS VPW NLVT11LL_CKT W=160.00n L=40.00n
XX12 net199 c pm VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS m net199 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX40 net244 SEN net188 VPW NLVT11LL_CKT W=160.00n L=40.00n
.ENDS LVT_SDQHSV1
****Sub-Circuit for LVT_SDQHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDQHSV2 CK D Q SE SI VDD VSS
XX41 net_0127 SI net_0123 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net_0123 SE VSS VPW NLVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn net_0127 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=180.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 s ps VSS VPW NLVT11LL_CKT W=160.00n L=40.00n
XX12 net52 c pm VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS m net52 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX40 net_0127 SEN net69 VPW NLVT11LL_CKT W=160.00n L=40.00n
XX7 net69 D VSS VPW NLVT11LL_CKT W=160.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX8 net0226 SEN net_0202 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX44 net_0202 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0202 SE VDD VNW PLVT11LL_CKT W=320.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX6 net0226 D net_0202 VNW PLVT11LL_CKT W=320.00n L=40.00n
XX9 pm c net0226 VNW PLVT11LL_CKT W=220.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD m net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=345.00n L=40.00n
.ENDS LVT_SDQHSV2
****Sub-Circuit for LVT_SDRNHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDRNHSV1 CK D Q QN RDN SE SI VDD VSS
XX13 VDD m net152 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX15 pm RDN VDD VNW PLVT11LL_CKT W=190.00n L=40.00n
XX32 QN ps VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX8 net192 SEN net195 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX44 net195 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX45 net195 SE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=190n L=40.00n
XX6 net192 D net195 VNW PLVT11LL_CKT W=240.00n L=40.00n
XX9 pm c net192 VNW PLVT11LL_CKT W=270.00n L=40.00n
XX22 s RDN VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net164 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net164 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net152 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX10 net283 RDN VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX7 net224 D net283 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX31 QN ps VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX16 VSS RDN net291 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX41 net284 SI net280 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net280 SE net283 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn net284 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=280.00n L=40.00n
XX21 s RDN net240 VPW NLVT11LL_CKT W=220.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net251 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net251 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX17 net240 ps VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net235 c pm VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net291 m net235 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX40 net284 SEN net224 VPW NLVT11LL_CKT W=140.00n L=40.00n
.ENDS LVT_SDRNHSV1
****Sub-Circuit for LVT_SDRNHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDRNHSV2 CK D Q QN RDN SE SI VDD VSS
XX10 net0159 RDN VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX31 QN ps VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX16 VSS RDN net0133 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX41 net_0127 SI net_0123 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net_0123 SE net0159 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn net_0127 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=280.00n L=40.00n
XX21 s RDN net0190 VPW NLVT11LL_CKT W=220.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net0190 ps VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net52 c pm VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 net0133 m net52 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX40 net_0127 SEN net69 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX7 net69 D net0159 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX15 pm RDN VDD VNW PLVT11LL_CKT W=190.00n L=40.00n
XX32 QN ps VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX8 net0226 SEN net_0202 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX44 net_0202 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0202 SE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=190n L=40.00n
XX6 net0226 D net_0202 VNW PLVT11LL_CKT W=240.00n L=40.00n
XX9 pm c net0226 VNW PLVT11LL_CKT W=270.00n L=40.00n
XX22 s RDN VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD m net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
.ENDS LVT_SDRNHSV2
****Sub-Circuit for LVT_SDRNQHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDRNQHSV1 CK D Q RDN SE SI VDD VSS
XX13 VDD m net140 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX15 pm RDN VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX8 net180 SEN net183 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX44 net183 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX45 net183 SE VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX6 net180 D net183 VNW PLVT11LL_CKT W=240.00n L=40.00n
XX9 pm c net180 VNW PLVT11LL_CKT W=240.00n L=40.00n
XX22 s RDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net152 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net152 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net140 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX7 net208 D net267 VPW NLVT11LL_CKT W=160.00n L=40.00n
XX10 net267 RDN VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX16 VSS RDN net275 VPW NLVT11LL_CKT W=130.00n L=40.00n
XX41 net268 SI net264 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net264 SE net267 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn net268 VPW NLVT11LL_CKT W=160.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=170.00n L=40.00n
XX21 s RDN net224 VPW NLVT11LL_CKT W=220.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net235 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net235 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX17 net224 ps VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net219 c pm VPW NLVT11LL_CKT W=130.00n L=40.00n
XX11 net275 m net219 VPW NLVT11LL_CKT W=130.00n L=40.00n
XX40 net268 SEN net208 VPW NLVT11LL_CKT W=160.00n L=40.00n
.ENDS LVT_SDRNQHSV1
****Sub-Circuit for LVT_SDRNQHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDRNQHSV2 CK D Q RDN SE SI VDD VSS
XX10 net0160 RDN VSS VPW NLVT11LL_CKT W=280.00n L=40.00n
XX16 VSS RDN net0133 VPW NLVT11LL_CKT W=130.00n L=40.00n
XX41 net_0127 SI net_0123 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net_0123 SE net0160 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn net_0127 VPW NLVT11LL_CKT W=160.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=170.00n L=40.00n
XX21 s RDN net0190 VPW NLVT11LL_CKT W=220.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 net0190 ps VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net52 c pm VPW NLVT11LL_CKT W=130.00n L=40.00n
XX11 net0133 m net52 VPW NLVT11LL_CKT W=130.00n L=40.00n
XX40 net_0127 SEN net69 VPW NLVT11LL_CKT W=160.00n L=40.00n
XX7 net69 D net0160 VPW NLVT11LL_CKT W=160.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX15 pm RDN VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX8 net0226 SEN net_0202 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX44 net_0202 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0202 SE VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX6 net0226 D net_0202 VNW PLVT11LL_CKT W=250.00n L=40.00n
XX9 pm c net0226 VNW PLVT11LL_CKT W=240.00n L=40.00n
XX22 s RDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD m net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
.ENDS LVT_SDRNQHSV2
****Sub-Circuit for LVT_SDRSNHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDRSNHSV1 CK D Q QN RDN SDN SE SI VDD VSS
XX25 net169 cn net305 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q net337 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX18 net161 net305 VDD VNW PLVT11LL_CKT W=395.00n L=40.00n
XX53 net337 net296 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX55 QN net296 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX39 net237 net337 net229 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX40 VDD rn net237 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX42 net229 c net296 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX54 VDD SDN net296 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX8 net177 SEN net180 VNW PLVT11LL_CKT W=215.00n L=40.00n
XX44 net180 SI VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX45 net180 SE VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX32 net161 SDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX9 net305 c net177 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 rn RDN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX33 net161 cn net296 VNW PLVT11LL_CKT W=265.00n L=40.00n
XX58 VDD RDN net305 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX31 net177 D net180 VNW PLVT11LL_CKT W=250.00n L=40.00n
XX26 VDD net161 net169 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX34 net313 SEN net249 VPW NLVT11LL_CKT W=180.00n L=40.00n
XX35 net249 D net312 VPW NLVT11LL_CKT W=180.00n L=40.00n
XX52 net337 net296 VSS VPW NLVT11LL_CKT W=315.00n L=40.00n
XX56 QN net296 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX48 net296 cn net325 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX49 net325 net337 net324 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX50 net296 rn net324 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX51 net324 SDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX41 net313 SI net309 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX43 net309 SE net312 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 net305 cn net313 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX16 rn RDN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX38 net161 c net296 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX57 VSS RDN net292 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=245.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net276 c net305 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX23 net292 net161 net276 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX19 Q net337 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX37 net161 SDN net261 VPW NLVT11LL_CKT W=285.00n L=40.00n
XX17 net261 net305 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX59 net312 RDN VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
.ENDS LVT_SDRSNHSV1
****Sub-Circuit for LVT_SDRSNHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDRSNHSV2 CK D Q QN RDN SDN SE SI VDD VSS
XX52 net205 net236 VSS VPW NLVT11LL_CKT W=315.00n L=40.00n
XX56 QN net236 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX48 net236 cn net193 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX49 net193 net205 net200 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX50 net236 rn net200 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX51 net200 SDN VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX41 net209 SI net213 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX43 net213 SE net0186 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX2 net0205 cn net209 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX16 rn RDN VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX38 net361 c net236 VPW NLVT11LL_CKT W=200.00n L=40.00n
XX57 VSS RDN net0220 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=245.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net252 c net0205 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX23 net0220 net361 net252 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX19 Q net205 VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX37 net361 SDN net257 VPW NLVT11LL_CKT W=285.00n L=40.00n
XX17 net257 net0205 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX59 net0186 RDN VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX34 net209 SEN net273 VPW NLVT11LL_CKT W=180.00n L=40.00n
XX35 net273 D net0186 VPW NLVT11LL_CKT W=180.00n L=40.00n
XX53 net205 net236 VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX55 QN net236 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX39 net289 net205 net297 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX40 VDD rn net289 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX42 net297 c net236 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX54 VDD SDN net236 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX8 net349 SEN net352 VNW PLVT11LL_CKT W=215.00n L=40.00n
XX44 net352 SI VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX45 net352 SE VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX32 net361 SDN VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX9 net0205 c net349 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX21 rn RDN VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX33 net361 cn net236 VNW PLVT11LL_CKT W=265.00n L=40.00n
XX58 VDD RDN net0205 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX31 net349 D net352 VNW PLVT11LL_CKT W=250.00n L=40.00n
XX26 VDD net361 net357 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net357 cn net0205 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q net205 VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 net361 net0205 VDD VNW PLVT11LL_CKT W=395.00n L=40.00n
.ENDS LVT_SDRSNHSV2
****Sub-Circuit for LVT_SDSNHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDSNHSV1 CK D Q QN SDN SE SI VDD VSS
XX49 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX43 net174 SDN VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX15 QN ps VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX33 net206 D net209 VNW PLVT11LL_CKT W=265.00n L=40.00n
XX8 net209 SE VDD VNW PLVT11LL_CKT W=320.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX6 net209 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX9 pm c net206 VNW PLVT11LL_CKT W=270.00n L=40.00n
XX50 VDD SDN ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX32 net206 SEN net209 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX4 net174 cn ps VNW PLVT11LL_CKT W=230.00n L=40.00n
XX44 net174 pm VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net158 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net158 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX14 net150 cn pm VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 VDD net174 net150 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX34 net290 D VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX41 net218 pm VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX45 VSS SDN net289 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX10 QN ps VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 pm cn net226 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX3 net174 c ps VPW NLVT11LL_CKT W=185.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX38 net258 SE VSS VPW NLVT11LL_CKT W=120.00n L=40.00n
XX24 net253 cn ps VPW NLVT11LL_CKT W=150.00n L=40.00n
XX23 net289 s net253 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX48 s ps VSS VPW NLVT11LL_CKT W=315.00n L=40.00n
XX12 net237 c pm VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS net174 net237 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX35 net226 SEN net290 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net226 SI net258 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX42 net174 SDN net218 VPW NLVT11LL_CKT W=285.00n L=40.00n
.ENDS LVT_SDSNHSV1
****Sub-Circuit for LVT_SDSNHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDSNHSV2 CK D Q QN SDN SE SI VDD VSS
XX34 net0150 D VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX45 VSS SDN net0333 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX10 QN ps VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX2 pm cn net_0127 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140n L=40.00n
XX3 net0266 c ps VPW NLVT11LL_CKT W=185.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX38 net_0162 SE VSS VPW NLVT11LL_CKT W=120.00n L=40.00n
XX24 net48 cn ps VPW NLVT11LL_CKT W=150.00n L=40.00n
XX23 net0333 s net48 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX48 s ps VSS VPW NLVT11LL_CKT W=315.00n L=40.00n
XX12 net52 c pm VPW NLVT11LL_CKT W=150.00n L=40.00n
XX11 VSS net0266 net52 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX35 net_0127 SEN net0150 VPW NLVT11LL_CKT W=150.00n L=40.00n
XX7 net_0127 SI net_0162 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX42 net0266 SDN net0206 VPW NLVT11LL_CKT W=290.00n L=40.00n
XX41 net0206 pm VSS VPW NLVT11LL_CKT W=290.00n L=40.00n
XX49 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX15 QN ps VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX33 net0224 D net0226 VNW PLVT11LL_CKT W=270.00n L=40.00n
XX8 net0226 SE VDD VNW PLVT11LL_CKT W=320.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210n L=40.00n
XX6 net0226 SI VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
XX9 pm c net0224 VNW PLVT11LL_CKT W=270.00n L=40.00n
XX50 VDD SDN ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX32 net0224 SEN net0226 VNW PLVT11LL_CKT W=140.00n L=40.00n
XX4 net0266 cn ps VNW PLVT11LL_CKT W=230.00n L=40.00n
XX44 net0266 pm VDD VNW PLVT11LL_CKT W=280.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX14 net117 cn pm VNW PLVT11LL_CKT W=150.00n L=40.00n
XX13 VDD net0266 net117 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX43 net0266 SDN VDD VNW PLVT11LL_CKT W=140.00n L=40.00n
.ENDS LVT_SDSNHSV2
****Sub-Circuit for LVT_SDXHSV1, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDXHSV1 CK DA DB Q QN SA SE SI VDD VSS
XX13 VDD m net169 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX10 QN ps VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX22 DA SAN net308 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX16 SAN SA VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX8 net205 SEN net208 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX32 DB SA net308 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX44 net208 SI VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX45 net208 SE VDD VNW PLVT11LL_CKT W=360.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX6 net205 net308 net208 VNW PLVT11LL_CKT W=340.00n L=40.00n
XX9 pm c net205 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net181 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net181 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net169 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX5 QN ps VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX7 net245 net308 VSS VPW NLVT11LL_CKT W=230.00n L=40.00n
XX21 DA SA net308 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX15 SAN SA VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX31 DB SAN net308 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX41 net249 SI net297 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net297 SE VSS VPW NLVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn net249 VPW NLVT11LL_CKT W=230.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=190.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net272 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net272 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX17 s ps VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net256 c pm VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS m net256 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX40 net249 SEN net245 VPW NLVT11LL_CKT W=230.00n L=40.00n
.ENDS LVT_SDXHSV1
****Sub-Circuit for LVT_SDXHSV2, Tue Sep 11 10:23:07 CST 2012****
.SUBCKT LVT_SDXHSV2 CK DA DB Q QN SA SE SI VDD VSS
XX5 QN ps VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX21 DA SA net0333 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX15 SAN SA VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX31 DB SAN net0333 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX41 net_0127 SI net_0123 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX43 net_0123 SE VSS VPW NLVT11LL_CKT W=120.00n L=40.00n
XX2 pm cn net_0127 VPW NLVT11LL_CKT W=230.00n L=40.00n
XX46 SEN SE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX3 m c ps VPW NLVT11LL_CKT W=190.00n L=40.00n
XX30 c cn VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 cn CK VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX24 net48 cn ps VPW NLVT11LL_CKT W=120.00n L=40.00n
XX23 VSS s net48 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX19 Q s VSS VPW NLVT11LL_CKT W=310.00n L=40.00n
XX17 s ps VSS VPW NLVT11LL_CKT W=220.00n L=40.00n
XX12 net52 c pm VPW NLVT11LL_CKT W=120.00n L=40.00n
XX11 VSS m net52 VPW NLVT11LL_CKT W=120.00n L=40.00n
XX40 net_0127 SEN net69 VPW NLVT11LL_CKT W=230.00n L=40.00n
XX7 net69 net0333 VSS VPW NLVT11LL_CKT W=230.00n L=40.00n
XX0 m pm VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX10 QN ps VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX22 DA SAN net0333 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX16 SAN SA VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX8 net0226 SEN net_0202 VNW PLVT11LL_CKT W=150.00n L=40.00n
XX32 DB SA net0333 VNW PLVT11LL_CKT W=210.00n L=40.00n
XX44 net_0202 SI VDD VNW PLVT11LL_CKT W=150.00n L=40.00n
XX45 net_0202 SE VDD VNW PLVT11LL_CKT W=360.00n L=40.00n
XX47 SEN SE VDD VNW PLVT11LL_CKT W=210.00n L=40.00n
XX6 net0226 net0333 net_0202 VNW PLVT11LL_CKT W=340.00n L=40.00n
XX9 pm c net0226 VNW PLVT11LL_CKT W=280.00n L=40.00n
XX4 m cn ps VNW PLVT11LL_CKT W=285.00n L=40.00n
XX29 c cn VDD VNW PLVT11LL_CKT W=380.00n L=40.00n
XX28 cn CK VDD VNW PLVT11LL_CKT W=130.00n L=40.00n
XX26 VDD s net109 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX25 net109 c ps VNW PLVT11LL_CKT W=120.00n L=40.00n
XX20 Q s VDD VNW PLVT11LL_CKT W=455.00n L=40.00n
XX18 s ps VDD VNW PLVT11LL_CKT W=370.00n L=40.00n
XX14 net117 cn pm VNW PLVT11LL_CKT W=120.00n L=40.00n
XX13 VDD m net117 VNW PLVT11LL_CKT W=120.00n L=40.00n
XX1 m pm VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
.ENDS LVT_SDXHSV2
****Sub-Circuit for LVT_TBUFHSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_TBUFHSV1 I OE Z VDD VSS
XX43 net080 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX44 net080 oen VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 oen OE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Z net080 VSS VPW NLVT11LL_CKT W=150.00n L=40.00n
XX36 net080 OE net_0163 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0163 OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX46 net_0163 I VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX28 oen OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX21 Z net_0163 VDD VNW PLVT11LL_CKT W=230.00n L=40.00n
XX39 net080 oen net_0163 VNW PLVT11LL_CKT W=200.00n L=40.00n
.ENDS LVT_TBUFHSV1
****Sub-Circuit for LVT_TBUFHSV12, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_TBUFHSV12 I OE Z VDD VSS
XX43 net080 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX44 net080 oen VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 oen OE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Z net080 VSS VPW NLVT11LL_CKT W=1.84u L=40.00n
XX36 net080 OE net_0163 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0163 OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX46 net_0163 I VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX28 oen OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX21 Z net_0163 VDD VNW PLVT11LL_CKT W=2.8u L=40.00n
XX39 net080 oen net_0163 VNW PLVT11LL_CKT W=200.00n L=40.00n
.ENDS LVT_TBUFHSV12
****Sub-Circuit for LVT_TBUFHSV16, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_TBUFHSV16 I OE Z VDD VSS
XX43 net080 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX44 net080 oen VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 oen OE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Z net080 VSS VPW NLVT11LL_CKT W=2.4u L=40.00n
XX36 net080 OE net_0163 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0163 OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX46 net_0163 I VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX28 oen OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX21 Z net_0163 VDD VNW PLVT11LL_CKT W=3.6u L=40.00n
XX39 net080 oen net_0163 VNW PLVT11LL_CKT W=200.00n L=40.00n
.ENDS LVT_TBUFHSV16
****Sub-Circuit for LVT_TBUFHSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_TBUFHSV2 I OE Z VDD VSS
XX43 net080 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX44 net080 oen VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 oen OE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Z net080 VSS VPW NLVT11LL_CKT W=300.00n L=40.00n
XX36 net080 OE net_0163 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0163 OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX46 net_0163 I VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX28 oen OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX21 Z net_0163 VDD VNW PLVT11LL_CKT W=460.00n L=40.00n
XX39 net080 oen net_0163 VNW PLVT11LL_CKT W=200.00n L=40.00n
.ENDS LVT_TBUFHSV2
****Sub-Circuit for LVT_TBUFHSV20, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_TBUFHSV20 I OE Z VDD VSS
XX43 net080 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX44 net080 oen VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 oen OE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Z net080 VSS VPW NLVT11LL_CKT W=2.99u L=40.00n
XX36 net080 OE net_0163 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0163 OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX46 net_0163 I VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX28 oen OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX21 Z net_0163 VDD VNW PLVT11LL_CKT W=4.55u L=40.00n
XX39 net080 oen net_0163 VNW PLVT11LL_CKT W=200.00n L=40.00n
.ENDS LVT_TBUFHSV20
****Sub-Circuit for LVT_TBUFHSV24, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_TBUFHSV24 I OE Z VDD VSS
XX43 net080 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX44 net080 oen VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 oen OE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Z net080 VSS VPW NLVT11LL_CKT W=3.68u L=40.00n
XX36 net080 OE net_0163 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0163 OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX46 net_0163 I VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX28 oen OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX21 Z net_0163 VDD VNW PLVT11LL_CKT W=5.6u L=40.00n
XX39 net080 oen net_0163 VNW PLVT11LL_CKT W=200.00n L=40.00n
.ENDS LVT_TBUFHSV24
****Sub-Circuit for LVT_TBUFHSV3, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_TBUFHSV3 I OE Z VDD VSS
XX43 net080 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX44 net080 oen VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 oen OE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Z net080 VSS VPW NLVT11LL_CKT W=460.00n L=40.00n
XX36 net080 OE net_0163 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0163 OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX46 net_0163 I VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX28 oen OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX21 Z net_0163 VDD VNW PLVT11LL_CKT W=700.00n L=40.00n
XX39 net080 oen net_0163 VNW PLVT11LL_CKT W=200.00n L=40.00n
.ENDS LVT_TBUFHSV3
****Sub-Circuit for LVT_TBUFHSV6, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_TBUFHSV6 I OE Z VDD VSS
XX43 net080 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX44 net080 oen VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 oen OE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Z net080 VSS VPW NLVT11LL_CKT W=920.00n L=40.00n
XX36 net080 OE net_0163 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0163 OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX46 net_0163 I VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX28 oen OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX21 Z net_0163 VDD VNW PLVT11LL_CKT W=1.4u L=40.00n
XX39 net080 oen net_0163 VNW PLVT11LL_CKT W=200.00n L=40.00n
.ENDS LVT_TBUFHSV6
****Sub-Circuit for LVT_TBUFHSV8, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_TBUFHSV8 I OE Z VDD VSS
XX43 net080 I VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX44 net080 oen VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX27 oen OE VSS VPW NLVT11LL_CKT W=140.00n L=40.00n
XX22 Z net080 VSS VPW NLVT11LL_CKT W=1.2u L=40.00n
XX36 net080 OE net_0163 VPW NLVT11LL_CKT W=140.00n L=40.00n
XX45 net_0163 OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX46 net_0163 I VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX28 oen OE VDD VNW PLVT11LL_CKT W=200.00n L=40.00n
XX21 Z net_0163 VDD VNW PLVT11LL_CKT W=1.8u L=40.00n
XX39 net080 oen net_0163 VNW PLVT11LL_CKT W=200.00n L=40.00n
.ENDS LVT_TBUFHSV8
****Sub-Circuit for LVT_XNOR2HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XNOR2HSV1 A1 A2 ZN VDD VSS
XX57 ZN xna1a2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX47 a2n A1 xna1a2 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX55 a2nn a2n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 a2nn a1n xna1a2 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX58 ZN xna1a2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX48 a2n a1n xna1a2 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX56 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX39 a2nn A1 xna1a2 VNW PLVT11LL_CKT W=300.00n L=40.00n
.ENDS LVT_XNOR2HSV1
****Sub-Circuit for LVT_XNOR2HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XNOR2HSV2 A1 A2 ZN VDD VSS
XX57 ZN xna1a2 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX47 a2n A1 xna1a2 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX55 a2nn a2n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 a2nn a1n xna1a2 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX58 ZN xna1a2 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX48 a2n a1n xna1a2 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX56 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX39 a2nn A1 xna1a2 VNW PLVT11LL_CKT W=300.00n L=40.00n
.ENDS LVT_XNOR2HSV2
****Sub-Circuit for LVT_XNOR3HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XNOR3HSV1 A1 A2 A3 ZN VDD VSS
XX47 net080 a3n xa1a2a3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 net080 net0107 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX60 a1nn A2 net0107 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX59 a1n a2n net0107 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX67 ZN xa1a2a3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX57 a3n A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX55 a1nn a1n VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 net0107 A3 xa1a2a3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=420.0n L=40.00n
XX58 a3n A3 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX62 a1nn a2n net0107 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX48 net080 A3 xa1a2a3 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX61 a1n A2 net0107 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX68 ZN xa1a2a3 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX56 a1nn a1n VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX1 net080 net0107 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX39 net0107 a3n xa1a2a3 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_XNOR3HSV1
****Sub-Circuit for LVT_XNOR3HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XNOR3HSV2 A1 A2 A3 ZN VDD VSS
XX47 net080 a3n xa1a2a3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 net080 net0107 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX60 a1nn A2 net0107 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX59 a1n a2n net0107 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX67 ZN xa1a2a3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX57 a3n A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX55 a1nn a1n VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 net0107 A3 xa1a2a3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=420.0n L=40.00n
XX58 a3n A3 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX62 a1nn a2n net0107 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX48 net080 A3 xa1a2a3 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX61 a1n A2 net0107 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX68 ZN xa1a2a3 VDD VNW PLVT11LL_CKT W=405.00n L=40.00n
XX56 a1nn a1n VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX1 net080 net0107 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX39 net0107 a3n xa1a2a3 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_XNOR3HSV2
****Sub-Circuit for LVT_XNOR4HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XNOR4HSV1 A1 A2 A3 A4 ZN VDD VSS
XX4 net0155 net0208 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX10 m net098 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX17 a3n A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX12 a4nn A3 net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX13 a4n a3n net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX20 a4n A4 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 a2nn a2n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX18 a4nn a4n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX23 net0148 net0155 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 n m VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX60 net0148 n net0109 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 ZN net0109 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX59 net0155 m net0109 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX65 a2nn A1 net0174 VPW NLVT11LL_CKT W=215.00n L=40.00n
XX66 a2n a1n net0174 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 net0208 net0174 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX22 a4n A4 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX15 a4n A3 net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX14 a4nn a3n net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX19 a3n A3 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX7 n m VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX24 net0148 net0155 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX21 a4nn a4n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX62 net0148 m net0109 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net0155 net0208 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX61 net0155 n net0109 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX63 a2nn a1n net0174 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX64 a2n A1 net0174 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX9 ZN net0109 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX3 net0208 net0174 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX11 m net098 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
.ENDS LVT_XNOR4HSV1
****Sub-Circuit for LVT_XNOR4HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XNOR4HSV2 A1 A2 A3 A4 ZN VDD VSS
XX4 net0155 net0208 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX10 m net098 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX17 a3n A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX12 a4nn A3 net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX13 a4n a3n net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX20 a4n A4 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 a2nn a2n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX18 a4nn a4n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX23 net0148 net0155 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 n m VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX60 net0148 n net0109 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 ZN net0109 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX59 net0155 m net0109 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX65 a2nn A1 net0174 VPW NLVT11LL_CKT W=215.00n L=40.00n
XX66 a2n a1n net0174 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 net0208 net0174 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX22 a4n A4 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX15 a4n A3 net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX14 a4nn a3n net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX19 a3n A3 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX7 n m VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX24 net0148 net0155 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX21 a4nn a4n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX62 net0148 m net0109 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net0155 net0208 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX61 net0155 n net0109 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX63 a2nn a1n net0174 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX64 a2n A1 net0174 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX9 ZN net0109 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX3 net0208 net0174 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX11 m net098 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
.ENDS LVT_XNOR4HSV2
****Sub-Circuit for LVT_XOR2HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XOR2HSV1 A1 A2 Z VDD VSS
XX57 Z xna1a2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX47 a2n a1n xna1a2 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX55 a2nn a2n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 a2nn A1 xna1a2 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX58 Z xna1a2 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX48 a2n A1 xna1a2 VNW PLVT11LL_CKT W=300.00n L=40.00n
XX56 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX39 a2nn a1n xna1a2 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_XOR2HSV1
****Sub-Circuit for LVT_XOR2HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XOR2HSV2 A1 A2 Z VDD VSS
XX57 Z xna1a2 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX47 a2n a1n xna1a2 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX55 a2nn a2n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 a2nn A1 xna1a2 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX58 Z xna1a2 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX48 a2n A1 xna1a2 VNW PLVT11LL_CKT W=300.00n L=40.00n
XX56 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX39 a2nn a1n xna1a2 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_XOR2HSV2
****Sub-Circuit for LVT_XOR3HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XOR3HSV1 A1 A2 A3 Z VDD VSS
XX47 net080 A3 xa1a2a3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 net080 net0107 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX60 a1nn A2 net0107 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX59 a1n a2n net0107 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX67 Z xa1a2a3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX57 a3n A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX55 a1nn a1n VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 net0107 a3n xa1a2a3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=420.0n L=40.00n
XX58 a3n A3 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX62 a1nn a2n net0107 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX48 net080 a3n xa1a2a3 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX61 a1n A2 net0107 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX68 Z xa1a2a3 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX56 a1nn a1n VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX1 net080 net0107 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX39 net0107 A3 xa1a2a3 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_XOR3HSV1
****Sub-Circuit for LVT_XOR3HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XOR3HSV2 A1 A2 A3 Z VDD VSS
XX47 net080 A3 xa1a2a3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 net080 net0107 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX60 a1nn A2 net0107 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX59 a1n a2n net0107 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX67 Z xa1a2a3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX57 a3n A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX55 a1nn a1n VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX36 net0107 a3n xa1a2a3 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=420.0n L=40.00n
XX58 a3n A3 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX62 a1nn a2n net0107 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX48 net080 a3n xa1a2a3 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX61 a1n A2 net0107 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX68 Z xa1a2a3 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX56 a1nn a1n VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX1 net080 net0107 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX39 net0107 A3 xa1a2a3 VNW PLVT11LL_CKT W=310.00n L=40.00n
.ENDS LVT_XOR3HSV2
****Sub-Circuit for LVT_XOR4HSV1, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XOR4HSV1 A1 A2 A3 A4 Z VDD VSS
XX4 net0155 net0208 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX10 m net098 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX17 a3n A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX12 a4n a3n net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX13 a4nn A3 net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX20 a4n A4 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 a2nn a2n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX18 a4nn a4n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX23 net0148 net0155 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 n m VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX60 net0148 m net0109 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 Z net0109 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX59 net0155 n net0109 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX65 a2nn A1 net0174 VPW NLVT11LL_CKT W=215.00n L=40.00n
XX66 a2n a1n net0174 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 net0208 net0174 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX22 a4n A4 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX15 a4nn a3n net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX14 a4n A3 net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX19 a3n A3 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX7 n m VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX24 net0148 net0155 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX21 a4nn a4n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX62 net0148 n net0109 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net0155 net0208 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX61 net0155 m net0109 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX63 a2nn a1n net0174 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX64 a2n A1 net0174 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX9 Z net0109 VDD VNW PLVT11LL_CKT W=315.00n L=40.00n
XX3 net0208 net0174 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX11 m net098 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
.ENDS LVT_XOR4HSV1
****Sub-Circuit for LVT_XOR4HSV2, Wed Sep  5 13:54:28 CST 2012****
.SUBCKT LVT_XOR4HSV2 A1 A2 A3 A4 Z VDD VSS
XX4 net0155 net0208 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX10 m net098 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX17 a3n A3 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX12 a4n a3n net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX13 a4nn A3 net098 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX20 a4n A4 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX0 a2nn a2n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX18 a4nn a4n VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX23 net0148 net0155 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX6 n m VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX49 a1n A1 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX60 net0148 m net0109 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX8 Z net0109 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX59 net0155 n net0109 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX65 a2nn A1 net0174 VPW NLVT11LL_CKT W=215.00n L=40.00n
XX66 a2n a1n net0174 VPW NLVT11LL_CKT W=210.00n L=40.00n
XX2 net0208 net0174 VSS VPW NLVT11LL_CKT W=285.00n L=40.00n
XX53 a2n A2 VSS VPW NLVT11LL_CKT W=210.00n L=40.00n
XX1 a2nn a2n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX22 a4n A4 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX15 a4nn a3n net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX14 a4n A3 net098 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX19 a3n A3 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX7 n m VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX24 net0148 net0155 VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX50 a1n A1 VDD VNW PLVT11LL_CKT W=250.00n L=40.00n
XX21 a4nn a4n VDD VNW PLVT11LL_CKT W=310.00n L=40.00n
XX62 net0148 n net0109 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX5 net0155 net0208 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX61 net0155 m net0109 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX63 a2nn a1n net0174 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX64 a2n A1 net0174 VNW PLVT11LL_CKT W=310.00n L=40.00n
XX54 a2n A2 VDD VNW PLVT11LL_CKT W=420.00n L=40.00n
XX9 Z net0109 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX3 net0208 net0174 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
XX11 m net098 VDD VNW PLVT11LL_CKT W=430.00n L=40.00n
.ENDS LVT_XOR4HSV2
