************************************************************************
* auCdl Netlist:
* 
* Library Name:  prima_sc180bcd_5v_9t_sch
* Top Cell Name: DFFSR_X1
* View Name:     schematic
* Netlisted on:  Apr 22 13:38:35 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    DFFSR_X1
* View Name:    schematic
************************************************************************

.SUBCKT DFFSR_X1 CLK D Q RN SN VDD VNW VPW VSS
*.PININFO CLK:I D:I RN:I SN:I Q:O VDD:B VNW:B VPW:B VSS:B
mNM13 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM39 net5 rnb net4 VPW nch5 mr=1 l=600n w=220n nf=1
mM19 Q net2 VSS VPW nch5 mr=1 l=600n w=1.15u nf=1
mM38 net4 SN VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM17 net1 clkn net5 VPW nch5 mr=1 l=600n w=220n nf=1
mM25 net7 net10 net8 VPW nch5 mr=1 l=600n w=220n nf=1
mM31 net7 D net12 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM28 net12 clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM22 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM34 rnb RN VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM7 net9 SN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM32 net10 clkp net1 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM9 net2 net1 VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM10 net10 rnb net9 VPW nch5 mr=1 l=600n w=735n nf=1
mNM3 net10 net7 net9 VPW nch5 mr=1 l=600n w=735n nf=1
mM24 net8 clkp VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM42 net5 net2 net4 VPW nch5 mr=1 l=600n w=220n nf=1
mM29 net6 clkp VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM43 net5 net2 net3 VNW pch5 mr=1 l=500n w=220n nf=1
mM27 net13 clkn VDD VNW pch5 mr=1 l=500n w=220n nf=1
mPM13 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM16 net1 clkp net5 VNW pch5 mr=1 l=500n w=220n nf=1
mM35 rnb RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM26 net7 net10 net13 VNW pch5 mr=1 l=500n w=220n nf=1
mM23 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM40 net5 SN VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM33 net10 clkn net1 VNW pch5 mr=1 l=500n w=1.03u nf=1
mM18 Q net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM6 net10 SN VDD VNW pch5 mr=1 l=500n w=1.01u nf=1
mPM3 net10 net7 net11 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM11 net11 rnb VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM30 net7 D net6 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM41 net3 rnb VDD VNW pch5 mr=1 l=500n w=220n nf=1
mPM9 net2 net1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
.ENDS

