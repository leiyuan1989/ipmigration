//* 
//* No part of this file can be released without the consent of SMIC.
//*
//******************************************************************************************
//* 0.18um Mixed Signal 1P6M with MIM Salicide 1.8V/3.3V RF SPICE Model (for SPECTRE only) *
//******************************************************************************************
//*
//* Release version    : 1.5
//*
//* Release date       : 12/22/2006
//*
//* Simulation tool    : Cadence spectre V6.0
//*
//*
//*  Inductor   :
//*
//*        *------------------------------* 
//*        | Inductor subckt |  ind_rf    |
//*        *------------------------------*
simulator lang=spectre  insensitive=yes
//*****************
//* 0.18um Inductor
//*****************
//* 1=port1(M6), 2=port2(M5)
//* R means inner redius; N means turns
//* Spacing is fixed at 1.5um and width is fixed at 8um
subckt ind_rf (1 2) 
parameters r=60u n=3.5 ls_rf=-1.7271-0.3612*n+0.2907*n*n+0.03256*r*1E6+0.000171*r*r*1E12 cf_rf=-25.41496+11.26813*n-1.25661*n*n+0.36097*r*1E6-0.0021636*r*r*1E12 rs_rf=-1.1605+0.66174*n+0.07719*n*n+0.02008*r*1E6+0.00011029*r*r*1E12
//* equivalent circuit
ls (1 4)      inductor    l=max(ls_rf*1E-9, 1E-12)
cf (1 3)      capacitor   c=max(cf_rf*1E-15, 1E-18)
rs (4 2)      resistor    r=max(rs_rf, 1E-6)
rsub1 (1  11) resistor    r=max(-481.30593+865.77248*ls_rf, 1E-6)
csub1 (11 12) capacitor   c=max((6.5234+1.4844*ls_rf)*1E-15, 1E-18)
lsub1 (12 10) inductor    l=max((0.44838+0.25562*ls_rf)*1E-9, 1E-15)
rsub2 (2  21) resistor    r=max(4.59004+142.22678*ls_rf, 1E-6)
csub2 (21 22) capacitor   c=max((6.12101+1.24623*ls_rf)*1E-15, 1E-18)
lsub2 (22 20) inductor    l=max((1.11853+0.04748*ls_rf)*1E-9, 1E-15)
rs2 (1 2)     resistor    r=max(7601.8+418.71024*ls_rf, 1E-6)
c11 (1 10)    capacitor   c=max((8.677+3.5886*ls_rf)*1E-15, 1E-18)
r11 (10 0)    resistor    r=max(66.08792+7.94856*ls_rf, 1E-6)
c22 (2 20)    capacitor   c=max((4.46577+3.65857*ls_rf)*1E-15, 1E-18)
r22 (20 0)    resistor    r=max(122.87152-5.8835*ls_rf, 1E-6)
r12 (3 2)     resistor    r=max(0.07804+0.00099619*ls_rf, 1E-6)
ends ind_rf
//*
