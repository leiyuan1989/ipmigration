* 
* No part of this file can be released without the consent of SMIC.
*
* Note: SMIC recommends that users set VNTOL=1E-9 at .option for more smooth convergence.
******************************************************************************************
* 0.18um Mixed Signal 1P6M with MIM Salicide 1.8V/3.3V RF SPICE Model (for HSPICE only)  *
******************************************************************************************
*
* Release version    : 1.5
*
* Release date       : 12/22/2006
*
* Simulation tool    : Synopsys Star-HSPICE version 2005.9
*
* Model type         :
*   MOSFET           : HSPICE Level 49(BSIM3V3.2)
*   Junction Diode   : HSPICE Level 3
* 
* Model and subcircuit name         :
*   MOSFET           :
*        *--------------------------------------*
*        |     MOSFET model   |  1.8V  |  3.3V  |
*        |======================================|
*        |        NMOS        | n18_rf | n33_rf |
*        *--------------------------------------*
*        |        PMOS        | p18_rf | p33_rf |
*        *--------------------------------------*
*
*        *----------------------------------------------*
*        |     MOSFET subckt  |    1.8V    |   3.3V     |
*        |==============================================|
*        |        NMOS        | n18_ckt_rf | n33_ckt_rf |
*        *----------------------------------------------*
*        |        PMOS        | p18_ckt_rf | p33_ckt_rf |
*        *----------------------------------------------*
*
*************************
* 1.8V RF NMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt n18_ckt_rf 1 2 3 4 lr=l wr=w nf=finger
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Rg_rf        = 'max((1542.7*lr*1e6+165.64)*pwr(wr*1e6,-0.9019*lr*1e6-0.5975)*pwr(nf,-0.9912*pwr(wr*1e6,-0.1348)), 1e-3)'
+Rsub1_rf     = 'max(341.64*pwr(nf,-0.5321), 1e-3)'
+Rsub2_rf     = 'max(341.64*pwr(nf,-0.5321), 1e-3)'
+Cgd_rf       = 'max(((8.85e-16*lr*lr*1e12-4.83e-16*lr*1e6+3.92e-16)*wr*1e6+2.95e-16)*nf+3.19e-16*pwr(wr*1e6,0.402), 1e-18)'
+Cgs_rf       = 'max(((4.82e-16*lr*1e6+9.58e-17)*pwr(wr*1e6,2.3513*lr*1e6-1.3178))*nf+1.34e-15*pwr(wr*1e6,-0.763), 1e-18)'
+Cds_rf       = 'max(((3.37e-17*pwr(lr*1e6,-1.38))*wr*1e6+1.89e-16)*nf+(-1.21e-14*lr*lr*1e12+9.83e-15*lr*1e6-9.86e-16)*pwr(wr*1e6,0.505), 1e-18)'
+Djdb_AREA_rf = '(nf/2*(0.8-2*0.07)*wr*1e6)*1e-12'
+Djdb_PJ_rf   = '(-0.048*log(wr*1e6)+1.1121)*(nf*wr)'
+Djsb_AREA_rf = '((nf/2-1)*(0.8-2*0.07)*wr*1e6+(0.8-0.07)*wr*1e6*2)*1e-12'
+Djsb_PJ_rf   = '(-0.0567*log(wr*1e6)+1.1608)*(nf*wr)'
+Rdc_n18      = 'max(17*(1/(pwr(wr*1e6,0.9))),1e-03)'
+Rsc_n18      = 'max(17*(1/(pwr(wr*1e6,0.9))),1e-03)'
+Cgdo_n18     = 'max((0+dcgdo_n18_rf), 0)'
+Cgso_n18     = 'max((0+dcgso_n18_rf), 0)'
+dt           = 'temper'
*****************************************
Lgate       2 20  1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 0.01
Ldrain       1 11 1p
Lsource      3 31 1p
*****************************************
Rjd   11 13 R='8.89e-09/Djdb_AREA_rf'
Djdb  12 13
+ ndio18_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
Cjdb  12 13 C='(9.68e-04+dcj_n18_rf)*(1+8.42e-04*(dt-25))*Djdb_AREA_rf*pwr((1+abs(V(13, 12))/0.7), -0.346)+(4.18e-10+dcjsw_n18_rf)*(1+6.69e-04*(dt-25))*Djdb_PJ_rf*pwr((1+abs(V(13, 12))/1), -0.538)' 
***
Rjs   31 33 R='8.89E-09/Djsb_AREA_rf'
Djsb  32 33
+ ndio18_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
Cjsb  32 33 C='(9.68e-04+dcj_n18_rf)*(1+8.42e-04*(dt-25))*Djsb_AREA_rf*pwr((1+abs(V(13, 12))/0.7), -0.346)+(4.18e-10+dcjsw_n18_rf)*(1+6.69e-04*(dt-25))*Djsb_PJ_rf*pwr((1+abs(V(13, 12))/1), -0.538)' 
*****************************************
Rsub1      41  4  Rsub1_rf
Rsub2      41  12 Rsub2_rf
Rsub3      41  32 12000
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 n18_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.MODEL n18_rf NMOS
+LEVEL = 49
*
* GENERAL PARAMETERS
*
+CALCACM  = 1
+LMIN     = 1.6E-7              LMAX     = 5.2E-7              WMIN     = 4.8E-7              
+WMAX     = 1.002E-5            TNOM     = 25.0                VERSION  = 3.2                 
+TOX      = '3.87E-09+DTOX_N18_RF' TOXM     = 3.87E-09            XJ       = 1.6000000E-07       
+NCH      = 3.8694000E+17       LLN      = 1.1205959           LWN      = 0.9200000           
+WLN      = 1.0599999           WWN      = 0.8768474           LINT     = 1.5757085E-08       
+LL       = 2.6352781E-16       LW       = -2.2625584E-16      LWL      = -2.0576711E-22      
+WINT     = -1.4450482E-09      WL       = -2.3664573E-16      WW       = -3.6409690E-14      
+WWL      = -4.0000000E-21      MOBMOD   = 1                   BINUNIT  = 2                   
+XL       = '1.8E-8+DXL_N18_RF'    XW       = '0.00+DXW_N18_RF'      DWG      = -5.9600000E-09      
+DWB      = 4.5000000E-09         
* DIODE PARAMETERS
+ACM      = 12                  LDIF     = 7.00E-08            HDIF     = 2.00E-07            
+RSH      = 7.08                RD       = 0                   RS       = 0                   
+RSC      = 'Rsc_n18'           RDC      = 'Rdc_n18'                 
*
* THRESHOLD VOLTAGE PARAMETERS
*
+VTH0     = '0.39+DVTH_N18_RF'     WVTH0    = -2.9709472E-08      PVTH0    = '5.0000000E-16+DPVTH0_N18_RF'       
+K1       = 0.6801043           WK1      = -2.4896840E-08      PK1      = 1.3000000E-15       
+K2       = -4.9977830E-02      K3       = 10.0000000          DVT0     = 1.3000000           
+DVT1     = 0.5771635           DVT2     = -0.1717554          DVT0W    = 0.00                
+DVT1W    = 0.00                DVT2W    = 0.00                NLX      = 7.5451030E-08       
+W0       = 5.5820150E-07       K3B      = -3.0000000                 
*
* MOBILITY PARAMETERS
*
+VSAT     = 8.2500000E+04       PVSAT    = -8.3000000E-10      UA       = -1.0300000E-09      
+LUA      = 7.7349790E-19       PUA      = -1.0000000E-24      UB       = 2.3666682E-18       
+UC       = 1.2000000E-10       PUC      = 1.5000000E-24       RDSW     = 55.5497200          
+PRWB     = -0.2400000          PRWG     = 0.4000000           WR       = 1.0000000           
+U0       = 3.4000000E-02       LU0      = 2.3057663E-11       WU0      = -3.1009695E-09      
+A0       = 0.8300000           KETA     = -3.0000000E-03      LKETA    = -1.7000000E-09      
+A1       = 0.00                A2       = 0.9900000           AGS      = 0.3200000           
+B0       = 6.0000000E-08       B1       = 0.00                
*
* SUBTHRESHOLD CURRENT PARAMETERS
*
+VOFF     = -0.1030000          LVOFF    = -3.3000000E-09      NFACTOR  = 1.2500000           
+LNFACTOR = 4.5000000E-08       CIT      = 0.00                CDSC     = 0.00                
+CDSCB    = 0.00                CDSCD    = 1.0000000E-04       ETA0     = 2.8000001E-02       
+ETAB     = -2.7000001E-02      DSUB     = 0.4000000           
*
* ROUT PARAMETERS
*
+PCLM     = 1.2000000           PPCLM    = 2.9999999E-15       PDIBLC1  = 2.5000000E-02       
+PDIBLC2  = 3.8000000E-03       PPDIBLC2 = 2.7000001E-16       PDIBLCB  = 0.00                
+DROUT    = 0.5600000           PSCBE1   = 3.4500000E+08       PSCBE2   = 1.0000000E-06       
+PVAG     = 0.00                DELTA    = 1.0000000E-02       ALPHA0   = 1.7753978E-08       
+ALPHA1   = 0.1764000           LALPHA1  = 7.6250000E-09       BETA0    = 11.1683940  
*
* TEMPERATURE EFFECTS PARAMETERS
*
+KT1      = -0.2572866          KT2      = -4.0000000E-02      AT       = 3.7000000E+04       
+PAT      = -7.5000000E-10      UTE      = -1.5500000          UA1      = 1.7600000E-09       
+LUA1     = 6.0000000E-18       WUA1     = -1.1000000E-16      PUA1     = -5.0000000E-25      
+UB1      = -2.4000000E-18      UC1      = -1.0000000E-10      LUC1     = 1.6999999E-17       
+PUC1     = -3.0000000E-24      KT1L     = -1.0000000E-09      PRT      = -55.0000000       
*
* CAPACITANCE PARAMETERS
*
+CJ       = 0                   MJ       = 0.346               PB       = 0.7                   
+CJSW     = 0                   MJSW     = 0.538               PBSW     = 1                 
+CJSWG    = 0                   MJSWG    = 0.538               PBSWG    = 1
+TCJ      = 8.42E-04            TCJSW    = 6.69E-04            TCJSWG   = 6.69E-04      
+TPB      = 1.47E-03            TPBSW    = 8.68E-04            TPBSWG   = 8.68E-04
+JS       = 3.52E-07            JSW      = 3.0E-13             NJ       = 1.0392 
+XTI      = 3.25                NQSMOD   = 0                   ELM      = 5
+CGDO     = 'Cgdo_n18'          CGSO     = 'Cgso_n18'          TLEVC    = 1            
+CAPMOD   = 3                   XPART    = 1                   CF       = 0.00                   
+ACDE     = 0.64                MOIN     = 24                  NOFF     = 1.2025                 
+DLC      = 8.5E-09             DWC      = 4.5E-08
+NLEV     = 3                   AF       = 0.85                KF       = 1.5E-24     
.model ndio18_rf D
+LEVEL    = 3                   JS       = 3.52e-07            JSW      = 1e-15            
+N        = 1.0233              IK       = 1.52e+05            
+IKR      = 2.78e+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.51e-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                             
+CJ       = 0                   CJSW     = 0                   RS       = 0
+MJ       = 0.346               PB       = 0.7                 MJSW     = 0.538               
+PHP      = 1                   CTA      = 0.000842            CTP      = 0.000669            
+TPB      = 0.00147             TPHP     = 0.000868            TLEV     = 1
+TLEVC    = 1                   FC       = 0                   FCS      = 0 
.ends n18_ckt_rf
*************************
* 1.8V RF PMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt p18_ckt_rf 1 2 3 4 lr=l wr=w nf=finger
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Rg_rf        = 'max((9852.3*lr*1e6-654.92)*pwr(wr*1e6,7.3896*lr*lr*1e12-5.4762*lr*1e6-0.0697)*pwr(nf,-1.0664*pwr(wr*1e6,2.8625*lr*lr*1e12-1.919*lr*1e6+0.2309)), 1e-3)'
+Rsub1_rf     = 'max(241.1*pwr(nf,-0.4726), 1e-3)'
+Rsub2_rf     = 'max(241.1*pwr(nf,-0.4726), 1e-3)'
+Cgd_rf       = 'max(((4.03e-16*lr*1e6+3.02e-16)*wr*1e6+3.06e-16)*nf+2.94e-16*pwr(wr*1e6,0.373), 1e-18)'
+Cgs_rf       = 'max((1.10e-15*pwr(wr*1e6,-0.367))*nf+(-1.06e-15*log(wr*1e6)+2.55e-15), 1e-18)'
+Cds_rf       = 'max((3.46e-16*wr*1e6+2.44e-16)*nf+(6.79e-17*wr*wr*1e12-3.13e-16*wr*1e6+1.17e-15), 1e-18)'
+Djdb_AREA_rf = '(nf/2*(0.8-2*0.07)*wr*1e6)*1e-12'
+Djdb_PJ_rf   = '(-0.0492*log(wr*1e6)+1.1146)*(nf*wr)'
+Djsb_AREA_rf = '((nf/2-1)*(0.8-2*0.07)*wr*1e6+(0.8-0.07)*wr*1e6*2)*1e-12'
+Djsb_PJ_rf   = '(-0.0582*log(wr*1e6)+1.1649)*(nf*wr)'
+Cgdo_p18     = 'max((0+dcgdo_p18_rf), 0)'
+Cgso_p18     = 'max((0+dcgso_p18_rf), 0)'
+dt           = 'temper'
*****************************************
Lgate       2 20  1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 0.01
Ldrain       1 11 1p
Lsource      3 31 1p
*****************************************
Rjd   11 13 R='8.77e-09/Djdb_AREA_rf'
Djdb  13 12
+ pdio18_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
Cjdb  13 12 C='(1.07E-03+dcj_p18_rf)*(1+8.76e-04*(dt-25))*Djdb_AREA_rf*pwr((1+abs(V(12, 13))/0.817), -0.415)+(5.07e-10+dcjsw_p18_rf)*(1+7.45e-04*(dt-25))*Djdb_PJ_rf*pwr((1+abs(V(12, 13))/1), -0.489)' 
***
Rjs   31 33 R='8.77e-09/Djsb_AREA_rf'
Djsb  33 32
+ pdio18_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
Cjsb  33 32 C='(1.07e-03+dcj_p18_rf)*(1+8.76e-04*(dt-25))*Djsb_AREA_rf*pwr((1+abs(V(12, 13))/0.817), -0.415)+(5.07e-10+dcjsw_p18_rf)*(1+7.45e-04*(dt-25))*Djsb_PJ_rf*pwr((1+abs(V(12, 13))/1), -0.489)' 
*****************************************
Rsub1      41  4  Rsub1_rf
Rsub2      41  12 Rsub2_rf
Rsub3      41  32 18000
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 p18_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.MODEL p18_rf PMOS
+LEVEL = 49
*
* GENERAL PARAMETERS
*
+CALCACM  = 1
+LMIN     = 1.6E-7              LMAX     = 5.2E-7              WMIN     = 4.8E-7              
+WMAX     = 1.002E-5            TNOM     = 25.0                VERSION  = 3.2                 
+TOX      = '3.74E-09+DTOX_P18_RF' TOXM     = 3.74E-09            XJ       = 1.7000001E-07       
+NCH      = 5.5000000E+17       LLN      = 1.0000000           LWN      = 1.0000000           
+WLN      = 1.0450000           WWN      = 1.0000000           LINT     = 1.0000000E-08       
+LL       = 3.4000000E-15       LW       = -3.3600000E-16      LWL      = 0.00                
+WINT     = 8.0000010E-09       WL       = 3.5904200E-15       WW       = -1.8999999E-15      
+WWL      = -1.1205000E-21      MOBMOD   = 1                   BINUNIT  = 2                   
+XL       = '-5.7E-09+DXL_P18_RF'  XW       = '0.00+DXW_P18_RF'      DWG      = -1.7361970E-08          
+DWB      = 2.0000000E-08       
* DIODE PARAMETERS
+ACM      = 12                  LDIF     = 7.00E-08            HDIF     = 2.00E-07            
+RSH      = 7.83                RD       = 0                   RS       = 0                   
+RSC      = 1.5                 RDC      = 1.5                 
*
* THRESHOLD VOLTAGE PARAMETERS
*
+VTH0     = '-0.402+DVTH_P18_RF'   WVTH0    = 1.2675420E-08       PVTH0    = '-1.2500000E-15+DPVTH0_P18_RF'      
+K1       = 0.5872390           LK1      = 3.5532110E-09       K2       = 7.0906860E-03       
+K3       = 2.5999999           DVT0     = 0.7194931           DVT1     = 0.2467441           
+DVT2     = 7.8089680E-02       DVT0W    = 0.00                DVT1W    = 8.0000000E+05       
+DVT2W    = 0.00                NLX      = 9.0000000E-08       W0       = 0.00                
+K3B      = 2.4862001           NGATE    = 3.1680000E+20               
*
* MOBILITY PARAMETERS
*
+VSAT     = 1.0000000E+05       UA       = 2.8500000E-10       LUA      = 5.5000000E-18       
+PUA      = -2.0000000E-24      UB       = 1.0000000E-18       UC       = -4.7700000E-11      
+WUC      = 3.1668000E-17       PUC      = -2.5000000E-24      RDSW     = 4.5500000E+02       
+PRWB     = -0.4000000          PRWG     = 0.00                WR       = 1.0000000           
+U0       = 8.6610000E-03       LU0      = -2.0000000E-11      WU0      = 1.3815350E-10       
+A0       = 1.0000000           KETA     = 2.0000000E-02       LKETA    = -8.5000000E-09      
+PKETA    = 5.0000000E-16       A1       = 0.00                A2       = 0.9900000           
+AGS      = 0.2000000           B0       = 6.3000000E-08       B1       = 0.00                
*
* SUBTHRESHOLD CURRENT PARAMETERS
*
+VOFF     = -9.5000000E-02      LVOFF    = -1.7000000E-09      WVOFF    = -1.9999999E-09      
+PVOFF    = -1.0000000E-16      NFACTOR  = 0.9000000           LNFACTOR = 1.0000000E-07       
+PNFACTOR = -5.0000000E-15      CIT      = 0.00                CDSC     = 0.00                
+CDSCB    = 0.00                CDSCD    = 0.00                ETA0     = 4.0000000E-02       
+ETAB     = -2.5000000E-02      DSUB     = 0.5600000           
*
* ROUT PARAMETERS
*
+PCLM     = 0.7000000           PDIBLC1  = 0.00                PDIBLC2  = 7.0000000E-03       
+PDIBLCB  = 0.00                DROUT    = 0.5600000           PSCBE1   = 4.0000000E+08       
+PSCBE2   = 1.0000000E-07       PVAG     = 0.00                DELTA    = 1.0000000E-02       
+ALPHA0   = 7.0000000E-08       ALPHA1   = 7.0491700           BETA0    = 22.8424000          
+LBETA0   = -7.5000000E-08         
*
* TEMPERATURE EFFECTS PARAMETERS
*
+KT1      = -0.2577007          KT2      = -3.0979900E-02      LKT2     = -3.0000000E-09      
+PKT2     = -6.5331750E-16      AT       = 1.0000000E+04       PAT      = -1.0000000E-09      
+UTE      = -1.2703574          UA1      = 5.3866300E-10       WUA1     = 1.1000000E-16       
+PUA1     = -2.3700001E-24      UB1      = -2.0709999E-18      UC1      = 2.0609721E-11       
+KT1L     = -8.0000000E-09      PRT      = 90.0000000          
*
* CAPACITANCE PARAMETERS
*
+CJ       = 0                   MJ       = 0.415               PB       = 0.817                   
+CJSW     = 0                   MJSW     = 0.489               PBSW     = 1               
+CJSWG    = 0                   MJSWG    = 0.489               PBSWG    = 1       
+TPB      = 0.00153             TPBSW    = 0.00117             TPBSWG   = 0.00117
+TCJ      = 0.000876            TCJSW    = 0.000745            TCJSWG   = 0.000745
+JS       = 1.66E-07            JSW      = 1.2E-13             NJ       = 1.0384   
+XTI      = 4.5                 NQSMOD   = 0                   ELM      = 5 
+CGDO     = 'Cgdo_p18'          CGSO     = 'Cgso_p18'          TLEVC    = 1            
+CAPMOD   = 3                   XPART    = 1                   CF       = 0.00                                    
+ACDE     = 0.8505076           MOIN     = 14.95341            NOFF     = 1.431824              
+DLC      = -1.5E-09
+NLEV     = 3                   AF       = 1.15                KF       = 3E-23        
.model pdio18_rf d
+LEVEL    = 3                   JS       = 1.66e-07            JSW      = 1e-15             
+N        = 1.0135              IK       = 4.03e+05            
+IKR      = 2.78e+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.78e-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                             
+CJ       = 0                   CJSW    = 0                    RS       = 0
+MJ       = 0.415               PB       = 0.817               MJSW     = 0.489               
+PHP      = 1                   CTA      = 0.000876            CTP      = 0.000745            
+TPB      = 0.00153             TPHP     = 0.00117             TLEV     = 1
+TLEVC    = 1                   FC       = 0                   FCS      = 0  
.ends p18_ckt_rf
*************************
* 3.3V RF NMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt n33_ckt_rf 1 2 3 4 lr=l wr=w nf=finger
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Rg_rf        = 'max((2182.1*lr*1e6+631.05)*pwr(nf,(-0.2332*lr*1e6-0.8064))*pwr((wr*1e6),((0.028*lr*1e6-0.003)*nf-0.385*lr*1e6-0.7245)),1e-3)'
+Cgd_rf       = 'max((((0.0583*lr*1e6+0.3367)*wr*1e6+(0.2972-0.0222*lr*1e6))*nf+0.4)*1E-15,1e-18)'
+Cgs_rf       = 'max((((2.4814*lr*1e6-0.1584)*log(wr*1e6)+(0.9772*lr*1e6+0.7258))*nf+(3.0576*lr*1e6+1.948))*1E-15,1e-18)'
+Cds_rf       = 'max((3.4-1.8*lr*1e6)*exp((0.047-0.038*lr*1e6)*nf*wr*1e6)*1E-15,1e-18)'
+Djdb_AREA_rf = '(nf/2*wr*1e6*(0.8-2*0.07))*1e-12'
+Djdb_PJ_rf   = '(1+4.0222e-6*wr*1e6+0.1771/(wr*1e6))*nf*wr'
+Djsb_AREA_rf = '(wr*1e6*(0.8-0.07)*2+(nf/2-1)*wr*1e6*(0.8-2*0.07))*1e-12'
+Djsb_PJ_rf   = '(1+4.0222e-6*wr*1e6+0.1771/(wr*1e6))*nf*wr'
+Rdc_n33      = 'max(50/(pwr(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.7)),1e-3)'
+Rsc_n33      = 'max(50/(pwr(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.7)),1e-3)'
+Cgdo_n33     = 'max((0+DCGDO_N33_RF),0)'
+Cgso_n33     = 'max((0+DCGSO_N33_RF),0)'
+dt           = 'temper'
*****************************************
Lgate       2 20 1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 1m
Ldrain      1 11 1p
Lsource     3 31 1p
*****************************************
Rjd   11 13 R='8.84E-09/Djdb_AREA_rf'
Djdb  12 13
+ ndio33_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
Cjdb  12 13 C='(0.000845+DCJ_N33_RF)*(1+0.000897*(dt-25))*Djdb_AREA_rf*pwr((1+abs(V(13, 12))/0.708), -0.321)+(3.41e-10+DCJSW_N33_RF)*(1+0.000695*(dt-25))*Djdb_PJ_rf*pwr((1+abs(V(13, 12))/1), -0.447)'
***
Rjs   31 33 R='8.84E-09/Djsb_AREA_rf'
Djsb  32 33
+ ndio33_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
Cjsb  32 33 C='(0.000845+DCJ_N33_RF)*(1+0.000897*(dt-25))*Djsb_AREA_rf*pwr((1+abs(V(33, 32))/0.708), -0.321)+(3.41e-10+DCJSW_N33_RF)*(1+0.000695*(dt-25))*Djsb_PJ_rf*pwr((1+abs(V(33, 32))/1), -0.447)'
*****************************************
Rsub1      41  4  150
Rsub2      41  12 500
Rsub3      41  32 500
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 n33_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.MODEL n33_rf NMOS
+LEVEL = 49
*
* GENERAL PARAMETERS
*
+CALCACM  = 1
+LMIN     = 3.3E-7              LMAX     = 5.2E-7              WMIN     = 4.8E-7              
+WMAX     = 1.002E-5            TNOM     = 25.0                VERSION  = 3.2                 
+TOX      = '6.65E-09+DTOX_N33_RF' TOXM     = 6.65E-09            XJ       = 1.6000000E-07       
+NCH      = 4.3441000E+17       LLN      = 1.0625758           LWN      = 1.0101005           
+WLN      = 0.9810000           WWN      = 0.9060000           LINT     = 6.3891300E-08       
+LL       = -2.3305548E-15      LW       = -2.4634918E-15      LWL      = 2.6243002E-24       
+WINT     = 3.5850000E-08       WL       = -1.8902563E-15      WW       = -1.3000000E-14      
+WWL      = -1.3027796E-20      MOBMOD   = 1                   BINUNIT  = 2                   
+XL       = '1E-8+DXL_N33_RF'   XW       = '0.00+DXW_N33_RF'   DWG      = -3.9100000E-09                  
+DWB      = 3.2000000E-09       
* DIODE PARAMETERS
+ACM      = 12                  LDIF     = 6.50E-08            HDIF     = 2.05E-07            
+RSH      = 7.08                RD       = 0                   RS       = 0                   
+RSC      = 'Rsc_n33'           RDC      = 'Rdc_n33'                 
*
* THRESHOLD VOLTAGE PARAMETERS
*
+VTH0     = '0.695+DVTH_N33_RF'    LVTH0    = 4.0100000E-10       WVTH0    = 1.0200000E-08       
+PVTH0    = '8.0000000E-16+DPVTH0_N33_RF'       K1       = 0.8451000           LK1      = 5.8182560E-10       
+WK1      = -6.2456240E-09      PK1      = 1.9938927E-15       K2       = 4.4575000E-02       
+K3       = -3.8500000          DVT0     = 9.4991400           LDVT0    = 8.0839730E-09       
+DVT1     = 0.6300000           LDVT1    = 5.5000000E-08       DVT2     = -0.1450000          
+DVT0W    = 0.00                DVT1W    = 0.1057000           DVT2W    = 0.00                
+NLX      = 2.0274594E-07       LNLX     = -2.8608589E-14      W0       = 0.00                
+K3B      = 0.5669292           NGATE    = 2.6812141E+21                 
*
* MOBILITY PARAMETERS
*
+VSAT     = 8.5000000E+04       LVSAT    = -1.7300000E-03      PVSAT    = 1.2000000E-10       
+UA       = -8.6001130E-10      UB       = 2.3000001E-18       UC       = 1.3100000E-10       
+PUC      = 5.0000000E-25       RDSW     = 2.4208382E+02       PRWB     = -8.5000000E-02      
+PRWG     = 3.8000000E-02       WR       = 1.0000000           U0       = 3.5000000E-02       
+LU0      = 5.0000000E-10       A0       = 1.0200000           LA0      = -1.2000000E-07      
+KETA     = 0.00                LKETA    = -1.4000000E-08      WKETA    = -1.9999999E-09      
+PKETA    = 1.0000000E-15       A1       = 0.00                A2       = 0.9900000           
+AGS      = 0.1700000           B0       = 1.0000000E-08       B1       = 0.00                
*
* SUBTHRESHOLD CURRENT PARAMETERS
*
+VOFF     = -0.1200000          NFACTOR  = 1.1000000           LNFACTOR = 4.0000000E-08       
+PNFACTOR = -1.4000000E-14      CIT      = 1.0000000E-04       CDSC     = 5.0000000E-04       
+CDSCB    = 0.00                CDSCD    = 0.00                ETA0     = 4.0000000E-02       
+PETA0    = 3.0000001E-16       ETAB     = -0.1000000          DSUB     = 0.6000000           
*
* ROUT PARAMETERS
*
+PCLM     = 0.8000000           LPCLM    = 5.0000000E-08       PPCLM    = 8.0000000E-15       
+PDIBLC1  = 9.0000000E-02       PDIBLC2  = 1.6000000E-03       PPDIBLC2 = -7.0000000E-17      
+PDIBLCB  = 0.00                DROUT    = 0.5987002           PSCBE1   = 3.4000000E+08       
+LPSCBE1  = 13.0000000          PSCBE2   = 3.8000000E-06       PVAG     = 0.00                
+DELTA    = 1.0000000E-02       ALPHA0   = -4.4760000E-08      ALPHA1   = 0.8998877           
+BETA0    = 18.8771250          LBETA0   = -5.7118000E-07
*
* TEMPERATURE EFFECTS PARAMETERS
*
+KT1      = -0.3250000          PKT1     = -2.3708420E-15      KT2      = -3.6844640E-02      
+AT       = 2.2000000E+04       UTE      = -1.4100000          UA1      = 2.0599999E-09       
+WUA1     = -1.2600000E-16      PUA1     = -1.0000000E-24      UB1      = -2.5000000E-18      
+WUB1     = 1.1000000E-25       UC1      = -1.1000000E-10      LUC1     = 1.6999999E-17       
+KT1L     = -5.0000000E-09      PRT      = 40.0000000          
*
* CAPACITANCE PARAMETERS
*
+CJ       = 0                   MJ       = 0.321               PB       = 0.708               
+CJSW     = 0                   MJSW     = 0.447               PBSW     = 1                   
+CJSWG    = 0                   MJSWG    = 0.447               PBSWG    = 1                   
+TPB      = 0.00166             TPBSW    = 0.00162             TPBSWG   = 0.00162     
+TCJ      = 0.000897            TCJSW    = 0.000695            TCJSWG   = 0.000695
+JS       = 3.65E-07            JSW      = 3.0E-13             NJ       = 1.04                 
+XTI      = 3.9                 NQSMOD   = 0                   ELM      = 5 
+CGDO     = 'Cgdo_n33'          CGSO     = 'Cgso_n33'          TLEVC    = 1 
+CAPMOD   = 3                   XPART    = 1                   CF       = 0.00                  
+ACDE     = 0.45                MOIN     = 24                  NOFF     = 2.3177            
+DLC      = 6.50E-08            NLEV     = 3                   AF       = 1
+KF       = 3E-23
.MODEL ndio33_rf D
+LEVEL    = 3                   JS       = 3.65E-07            JSW      = 1E-15            
+N        = 1.0203              RS       = 0                   IK       = 1.33E+05            
+IKR      = 2.78E+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.07E-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                 CJ       = 0                   MJ       = 0.321               
+PB       = 0.708               CJSW     = 0                   MJSW     = 0.447               
+PHP      = 1                   CTA      = 0.000897            CTP      = 0.000695            
+TPB      = 0.00166             TPHP     = 0.00162             TLEV     = 1
+TLEVC    = 1                   FC       = 0                   FCS      = 0
.ends n33_ckt_rf
*************************
* 3.3V RF PMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt p33_ckt_rf 1 2 3 4 lr=l wr=w nf=finger
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+Rg_rf        = 'max((6345.5*lr*1e6+389.25)*pwr(nf,(0.303*lr*1e6-1.1215))*pwr((wr*1e6),(-0.6785*lr*1e6-0.4944)),1e-3)'
+Cgd_rf       = 'max(((0.1595*lr*1e6+0.2682)*wr*1e6*nf+(0.255+0.058*lr*1e6)*nf+0.8393-1.1375*lr*1e6)*1e-15,1e-18)'
+Cgs_rf       = 'max((((0.3785-0.0165*lr*1e6)*wr*1e6+(0.9772*lr*1e6+0.1732))*nf+4)*1e-15,1e-18)'
+Cds_rf       = 'max(((0.8638-0.8045*lr*1e6)*wr*1e6+(1.9425*lr*1e6-0.7838))*nf*1e-15,1e-18)'
+Djdb_AREA_rf = '(nf/2*wr*1e6*(0.8-2*0.07))*1e-12'
+Djdb_PJ_rf   = '(1-6.0826e-6*wr*1e6+0.1854/wr*1e6)*nf*wr'
+Djsb_AREA_rf = '(wr*1e6*(0.8-0.07)*2+(nf/2-1)*wr*1e6*(0.8-2*0.07))*1e-12'
+Djsb_PJ_rf   = '(1-6.0826e-6*wr*1e6+0.1854/wr*1e6)*nf*wr'
+Rdc_p33      = 'max(81.5/(pwr(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.95)),1e-3)'
+Rsc_p33      = 'max(81.5/(pwr(((1-wr*1e6)/(wr*1e6)+wr*1e6),0.95)),1e-3)'
+Cgdo_p33     = 'max((0+DCGDO_P33_RF),0)'
+Cgso_p33     = 'max((0+DCGSO_P33_RF),0)'
+dt           = 'temper'
*****************************************
Lgate       2 20 1p
Rgate       20 21 Rg_rf
Cgd_ext     20 11 Cgd_rf
Cgs_ext     20 31 Cgs_rf
Cds_ext     15 31 Cds_rf
Rds         11 15 80.2
Ldrain      1 11 1p
Lsource     3 31 1p
*****************************************
Rjd   11 13 R='9.23E-09/Djdb_AREA_rf'
Djdb  12 13
+ pdio33_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
Cjdb  13 12 C='(0.00101+DCJ_P33_RF)*(1+0.000883*(dt-25))*Djdb_AREA_rf*pwr((1+abs(V(12, 13))/0.807), -0.401)+(3.19e-10+DCJSW_P33_RF)*(1+0.000709*(dt-25))*Djdb_PJ_rf*pwr((1+abs(V(12, 13))/1), -0.45)'
***
Rjs   31 33 R='9.23E-09/Djsb_AREA_rf'
Djsb  32 33
+ pdio33_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
Cjsb  33 32 C='(0.00101+DCJ_P33_RF)*(1+0.000883*(dt-25))*Djsb_AREA_rf*pwr((1+abs(V(32, 33))/0.807), -0.401)+(3.19e-10+DCJSW_P33_RF)*(1+0.000709*(dt-25))*Djsb_PJ_rf*pwr((1+abs(V(32, 33))/1), -0.45)'
*****************************************
Rsub1      41  4  10
Rsub2      41  12 50000
Rsub3      41  32 50000
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 p33_rf L=lr W=wr m=nf AD = 0 AS = 0 PD = 0 PS = 0
* MOS Model
.MODEL p33_rf PMOS
+LEVEL = 49
*
* GENERAL PARAMETERS
*
+CALCACM  = 1
+LMIN     = 2.8E-7              LMAX     = 5.2E-7              WMIN     = 4.8E-7              
+WMAX     = 1.002E-5            TNOM     = 25.0                VERSION  = 3.2                 
+TOX      = '6.62E-09+DTOX_P33_RF' TOXM     = 6.62E-09            XJ       = 1.7000001E-07       
+NCH      = 5.4852000E+17       LLN      = 1.0471729           LWN      = 0.9530895           
+WLN      = 1.0257638           WWN      = 0.9617700           LINT     = 3.5000000E-08       
+LL       = 5.5000000E-15       LW       = -4.7160380E-14      LWL      = 7.0054450E-22       
+WINT     = 1.3000000E-08       WL       = -3.1491245E-14      WW       = 2.3000000E-15       
+WWL      = -2.4167156E-22      MOBMOD   = 1                   BINUNIT  = 2                   
+XL       = '-1.70E-08+DXL_P33_RF' XW       = '0.00+DXW_P33_RF'      DWG      = 0.00                   
+DWB      = 8.6000000E-09                                 
* DIODE PARAMETERS
+ACM      = 12                  LDIF     = 6.50E-08            HDIF     = 2.05E-07            
+RSH      = 9.8                 RD       = 0                   RS       = 0                   
+RSC      = 'Rsc_p33'           RDC      = 'Rdc_p33'                   
*
* THRESHOLD VOLTAGE PARAMETERS
*
+VTH0     = '-0.672+DVTH_P33_RF'   WVTH0    = 4.0000000E-09       PVTH0    = '6.0000000E-15+DPVTH0_P33_RF'       
+K1       = 0.9145741           PK1      = -1.7000000E-14      K2       = 4.1276220E-02       
+K3       = 0.1293833           DVT0     = 1.8000000           DVT1     = 0.7100000           
+DVT2     = -7.0000000E-02      DVT0W    = 0.00                DVT1W    = 0.00                
+DVT2W    = 0.00                NLX      = 1.2000000E-08       W0       = 1.0021131E-09       
+K3B      = 0.4000000           NGATE    = 1.1600000E+20               
*
* MOBILITY PARAMETERS
*
+VSAT     = 8.5500000E+04       PVSAT    = -5.8000000E-09      UA       = 3.1500000E-10       
+LUA      = 1.5000001E-17       WUA      = -1.6763224E-16      PUA      = -1.1000000E-23      
+UB       = 1.0444180E-18       LUB      = -7.0000000E-27      UC       = -3.5000000E-11      
+LUC      = 4.0000000E-18       PUC      = 5.0000000E-24       RDSW     = 9.5000000E+02       
+PRWB     = 0.00                PRWG     = 6.3755660E-03       WR       = 1.0000000           
+U0       = 9.2500000E-03       LU0      = -4.1500680E-10      WU0      = -1.7001526E-12      
+PU0      = -3.7999640E-16      A0       = 0.8500000           KETA     = 1.5000000E-02       
+LKETA    = -1.0000000E-08      WKETA    = 1.0000000E-09       PKETA    = -6.0000000E-15      
+A1       = 0.00                A2       = 0.9900000           AGS      = 4.0000000E-02       
+B0       = 4.6000000E-08       B1       = 0.00                
*
* SUBTHRESHOLD CURRENT PARAMETERS
*
+VOFF     = -0.1000000          LVOFF    = 1.8000000E-09       PVOFF    = -2.9999999E-15      
+NFACTOR  = 1.1000000           PNFACTOR = -4.0000000E-14      CIT      = 1.9999999E-04       
+CDSC     = 4.5263850E-05       CDSCB    = 0.00                CDSCD    = 0.00                
+ETA0     = 5.0000000E-03       PETA0    = 7.0000000E-15       ETAB     = -1.5000000E-02      
+PETAB    = -2.0000000E-15      DSUB     = 0.5800000           
*
* ROUT PARAMETERS
*
+PCLM     = 0.6000000           PPCLM    = 1.3000000E-13       PDIBLC1  = 6.0000000E-03       
+PDIBLC2  = 2.5000001E-04       WPDIBLC2 = 8.0000000E-11       PDIBLCB  = 0.00                
+DROUT    = 0.5600000           PSCBE1   = 3.3000000E+08       PPSCBE1  = -7.0000000E-06      
+PSCBE2   = 2.0000000E-07       PVAG     = 0.00                DELTA    = 8.0000000E-03       
+PDELTA   = 4.0000000E-16       ALPHA0   = 1.3410400E-06       ALPHA1   = 5.6136910E-02       
+BETA0    = 27.5998000          
*
* TEMPERATURE EFFECTS PARAMETERS
*
+KT1      = -0.3840900          WKT1     = -9.4333370E-10      PKT1     = 4.9999980E-15       
+KT2      = -4.1563480E-02      AT       = -2.0000000E+03      PAT      = -7.5000000E-09      
+UTE      = -1.3236057          UA1      = 3.0000002E-10       WUA1     = 8.0000000E-18       
+PUA1     = 1.0000000E-23       UB1      = -2.0704662E-18      WUB1     = 1.4000000E-25       
+UC1      = -5.0000000E-11      KT1L     = -6.0000000E-09      PRT      = 1.3000000E+02
*
* CAPACITANCE PARAMETERS
*
+CJ       = 0                   MJ       = 0.401               PB       = 0.807
+CJSW     = 0                   MJSW     = 0.45                PBSW     = 1
+CJSWG    = 0                   MJSWG    = 0.45                PBSWG    = 1
+TPB      = 0.00157             TPBSW    = 0.00137             TPBSWG   = 0.00137
+TCJ      = 0.000883            TCJSW    = 0.000709            TCJSWG   = 0.000709
+JS       = 1.68E-07            JSW      = 4.0E-13             NJ       = 1.07
+XTI      = 3.0                 NQSMOD   = 0                   ELM      = 5
+CGDO     = 'Cgdo_p33'          CGSO     = 'Cgso_p33'          TLEVC    = 1
+CAPMOD   = 3                   XPART    = 1                   CF       = 0.00
+ACDE     = 0.55                MOIN     = 15                  NOFF     = 0.565
+DLC      = 7.0E-09             DWC      = 6.0E-8 
+NLEV     = 3                   AF       = 1.02                KF       = 3E-23
.MODEL pdio33_rf D
+LEVEL    = 3                   JS       = 1.68E-07            JSW      = 1E-15            
+N        = 1.0143              RS       = 0                   IK       = 4.07E+05            
+IKR      = 2.78E+05            BV       = 11.0                IBV      = 277.78              
+TRS      = 1.24E-03            EG       = 1.16                TREF     = 25.0                
+XTI      = 3.0                 CJ       = 0                   MJ       = 0.401               
+PB       = 0.807               CJSW     = 0                   MJSW     = 0.45                
+PHP      = 1                   CTA      = 0.000883            CTP      = 0.000709            
+TPB      = 0.00157             TPHP     = 0.00137             TLEV     = 1
+TLEVC    = 1                   FC       = 0                   FCS      = 0 
.ends p33_ckt_rf
