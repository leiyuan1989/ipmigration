.SUBCKT AOI222_X1 A1 A2 B1 B2 C1 C2 VDD VSS ZN
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:B VNW:B VPW:B VSS:B
mPM10 net2 B2 net1 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM9 net2 B1 net1 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM2 ZN A1 net2 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM1 ZN A2 net2 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM7 net1 C2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM6 net1 C1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mNM9 ZN C1 net4 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM3 ZN A1 net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM1 net6 A2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM8 ZN B1 net5 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM6 net5 B2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 net4 C2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    DLY_X1
* View Name:    schematic
************************************************************************

.SUBCKT DLY_X1 A VDD VSS Z
*.PININFO A:I Z:O VDD:B VNW:B VPW:B VSS:B
mM5 Z N0 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM9 N1 A VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM3 N0 N2 VSS VPW nch5 mr=1 l=1.74u w=610n nf=1
mM0 N2 N1 VSS VPW nch5 mr=1 l=930n w=610n nf=1
mM4 Z N0 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM9 N1 A VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM2 N0 N2 VDD VNW pch5 mr=1 l=1.74u w=870n nf=1
mM1 N2 N1 VDD VNW pch5 mr=1 l=930n w=870n nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    ADDF_X1
* View Name:    schematic
************************************************************************

.SUBCKT ADDF_X1 A B CI CO S VDD VSS
*.PININFO A:I B:I CI:I CO:O S:O VDD:B VNW:B VPW:B VSS:B
mM6 N0 B VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM0 N1 A VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM13 N2 B VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM3 N3 CI N1 VPW nch5 mr=1 l=600n w=610n nf=1
mM1 N1 B VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM19 N4 N3 N5 VPW nch5 mr=1 l=600n w=610n nf=1
mM17 N4 CI N6 VPW nch5 mr=1 l=600n w=610n nf=1
mM21 N5 CI VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM11 N5 A VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM23 S N4 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM10 N5 B VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM25 CO N3 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM4 N3 A N0 VPW nch5 mr=1 l=600n w=610n nf=1
mM15 N6 A N2 VPW nch5 mr=1 l=600n w=610n nf=1
mM26 CO N3 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM2 N3 CI N7 VNW pch5 mr=1 l=500n w=870n nf=1
mM12 N8 A VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM18 N4 CI N9 VNW pch5 mr=1 l=500n w=870n nf=1
mM16 N9 A N10 VNW pch5 mr=1 l=500n w=870n nf=1
mM14 N10 B VDD VNW pch5 mr=1 l=500n w=870n nf=1
mPM0 N7 A VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM22 N8 CI VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM20 N4 N3 N8 VNW pch5 mr=1 l=500n w=870n nf=1
mPM1 N7 B VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM24 S N4 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM7 N11 B VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM5 N3 A N11 VNW pch5 mr=1 l=500n w=870n nf=1
mM9 N8 B VDD VNW pch5 mr=1 l=500n w=870n nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    AO222_X1
* View Name:    schematic
************************************************************************

.SUBCKT AO222_X1 A1 A2 B1 B2 C1 C2 VDD VSS Z
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I Z:O VDD:B VNW:B VPW:B VSS:B
mPM6 net1 C1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM10 net2 B2 net1 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM9 net2 B1 net1 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM2 net7 A1 net2 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM1 net7 A2 net2 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM7 net1 C2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM5 Z net7 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mNM1 net6 A2 VSS VPW nch5 mr=1 l=600n w=1u nf=1
mNM3 net7 A1 net6 VPW nch5 mr=1 l=600n w=1u nf=1
mNM9 net7 C1 net4 VPW nch5 mr=1 l=600n w=1u nf=1
mNM6 net5 B2 VSS VPW nch5 mr=1 l=600n w=1u nf=1
mM0 net4 C2 VSS VPW nch5 mr=1 l=600n w=1u nf=1
mNM8 net7 B1 net5 VPW nch5 mr=1 l=600n w=1u nf=1
mNM4 Z net7 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    MUX4_X1
* View Name:    schematic
************************************************************************

.SUBCKT MUX4_X1 I0 I1 I2 I3 S0 S1 VDD VSS Z
*.PININFO I0:I I1:I I2:I I3:I S0:I S1:I Z:O VDD:B VNW:B VPW:B VSS:B
mM19 N0 I3 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM16 N1 S0 N0 VPW nch5 mr=1 l=600n w=610n nf=1
mM12 N2 I2 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM10 N3 I1 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM6 N4 N5 N6 VPW nch5 mr=1 l=600n w=610n nf=1
mM0 Z N7 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM4 N6 I0 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM8 N4 S0 N3 VPW nch5 mr=1 l=600n w=610n nf=1
mNM0 N8 S1 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM15 N1 N5 N2 VPW nch5 mr=1 l=600n w=610n nf=1
mM22 N7 S1 N1 VPW nch5 mr=1 l=600n w=610n nf=1
mNM12 N5 S0 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mM21 N7 N8 N4 VPW nch5 mr=1 l=600n w=610n nf=1
mM18 N1 N5 N9 VNW pch5 mr=1 l=500n w=870n nf=1
mM14 N1 S0 N10 VNW pch5 mr=1 l=500n w=870n nf=1
mM13 N10 I2 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM11 N11 I1 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM7 N4 S0 N12 VNW pch5 mr=1 l=500n w=870n nf=1
mM1 Z N7 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM5 N12 I0 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM9 N4 N5 N11 VNW pch5 mr=1 l=500n w=870n nf=1
mM23 N7 N8 N1 VNW pch5 mr=1 l=500n w=870n nf=1
mPM0 N8 S1 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM20 N9 I3 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mPM12 N5 S0 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mM24 N7 S1 N4 VNW pch5 mr=1 l=500n w=870n nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    NAND4_X1
* View Name:    schematic
************************************************************************

.SUBCKT NAND4_X1 A1 A2 A3 A4 VDD VSS ZN
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:B VNW:B VPW:B VSS:B
mPM1 ZN A4 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM3 ZN A2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM2 ZN A3 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM4 ZN A1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mNM2 ZN A1 net28 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM1 net28 A2 net27 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM3 net29 A4 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM0 net27 A3 net29 VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    AND4_X1
* View Name:    schematic
************************************************************************

.SUBCKT AND4_X1 A1 A2 A3 A4 VDD VSS Z
*.PININFO A1:I A2:I A3:I A4:I Z:O VDD:B VNW:B VPW:B VSS:B
mPM0 Z net6 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM1 net6 A4 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mPM2 net6 A3 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mPM3 net6 A2 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mPM4 net6 A1 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mNM2 net6 A1 net12 VPW nch5 mr=1 l=600n w=1u nf=1
mNM3 net10 A4 VSS VPW nch5 mr=1 l=600n w=1u nf=1
mNM4 Z net6 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM0 net11 A3 net10 VPW nch5 mr=1 l=600n w=1u nf=1
mNM1 net12 A2 net11 VPW nch5 mr=1 l=600n w=1u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    NOR4_X1
* View Name:    schematic
************************************************************************

.SUBCKT NOR4_X1 A1 A2 A3 A4 VDD VSS ZN
*.PININFO A1:I A2:I A3:I A4:I ZN:O VDD:B VNW:B VPW:B VSS:B
mNM4 ZN A1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM3 ZN A2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM1 ZN A4 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM0 ZN A3 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mPM4 net49 A1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM3 net48 A2 net49 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM1 net47 A3 net48 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM0 ZN A4 net47 VNW pch5 mr=1 l=500n w=1.74u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    OR4_X1
* View Name:    schematic
************************************************************************

.SUBCKT OR4_X1 A1 A2 A3 A4 VDD VSS Z
*.PININFO A1:I A2:I A3:I A4:I Z:O VDD:B VNW:B VPW:B VSS:B
mNM4 net27 A1 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mNM3 net27 A2 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mNM2 Z net27 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM1 net27 A4 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mNM0 net27 A3 VSS VPW nch5 mr=1 l=600n w=610n nf=1
mPM4 net36 A1 VDD VNW pch5 mr=1 l=500n w=870n nf=1
mPM3 net34 A2 net36 VNW pch5 mr=1 l=500n w=870n nf=1
mPM2 Z net27 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM1 net33 A3 net34 VNW pch5 mr=1 l=500n w=870n nf=1
mPM0 net27 A4 net33 VNW pch5 mr=1 l=500n w=870n nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    OAI33_X1
* View Name:    schematic
************************************************************************

.SUBCKT OAI33_X1 A1 A2 A3 B1 B2 B3 VDD VSS ZN
*.PININFO A1:I A2:I A3:I B1:I B2:I B3:I ZN:O VDD:B VNW:B VPW:B VSS:B
mM2 net40 A2 net41 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM1 ZN A3 net40 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM6 net42 B1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM10 net43 B2 net42 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM3 net41 A1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM7 ZN B3 net43 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM18 net6 A1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM17 net6 A3 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM11 ZN B3 net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM9 ZN B2 net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM8 ZN B1 net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM19 net6 A2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    BUF_X1
* View Name:    schematic
************************************************************************

.SUBCKT BUF_X1 A VDD VSS Z
*.PININFO A:I Z:O VDD:B VNW:B VPW:B VSS:B
mPM1 Z net08 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM0 net08 A VDD VNW pch5 mr=1 l=500n w=870n nf=1
mNM0 net08 A VSS VPW nch5 mr=1 l=600n w=610n nf=1
mNM1 Z net08 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    OA222_X1
* View Name:    schematic
************************************************************************

.SUBCKT OA222_X1 A1 A2 B1 B2 C1 C2 VDD VSS Z
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I Z:O VDD:B VNW:B VPW:B VSS:B
mM18 net5 A1 net7 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM16 Z net5 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM19 net7 A2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM11 net8 C2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM10 net5 C1 net8 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM9 net5 B1 net6 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM7 net6 B2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM13 net15 B1 net1 VPW nch5 mr=1 l=600n w=1u nf=1
mM12 net15 B2 net1 VPW nch5 mr=1 l=600n w=1u nf=1
mM17 net1 C2 VSS VPW nch5 mr=1 l=600n w=1u nf=1
mM20 net1 C1 VSS VPW nch5 mr=1 l=600n w=1u nf=1
mM8 net5 A1 net15 VPW nch5 mr=1 l=600n w=1u nf=1
mM6 net5 A2 net15 VPW nch5 mr=1 l=600n w=1u nf=1
mM15 Z net5 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    OAI222_X1
* View Name:    schematic
************************************************************************

.SUBCKT OAI222_X1 A1 A2 B1 B2 C1 C2 VDD VSS ZN
*.PININFO A1:I A2:I B1:I B2:I C1:I C2:I ZN:O VDD:B VNW:B VPW:B VSS:B
mM18 ZN A1 net4 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM19 net4 A2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM10 ZN C1 net3 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM11 net3 C2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM7 net1 B2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM9 ZN B1 net1 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM6 ZN A2 net119 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM12 net119 B2 net108 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM17 net108 C2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM20 net108 C1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM13 net119 B1 net108 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM8 ZN A1 net119 VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    XOR3_X1
* View Name:    schematic
************************************************************************

.SUBCKT XOR3_X1 A1 A2 A3 VDD VSS Z
*.PININFO A1:I A2:I A3:I Z:O VDD:B VNW:B VPW:B VSS:B
mM2 N0 A2 N1 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM8 N2 A1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM27 N0 N3 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM37 N3 A2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM30 N4 N2 N5 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM5 N1 A3 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM29 N5 N0 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM33 N4 A1 N0 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM14 N3 A3 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM36 Z N4 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM7 N2 A1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM25 N6 A2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM35 Z N4 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM32 N7 N0 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM26 N0 N3 N6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM31 N4 A1 N7 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM34 N4 N2 N0 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM24 N6 A3 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM13 N3 A3 N8 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM28 N8 A2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    DFFSR_X1
* View Name:    schematic
************************************************************************

.SUBCKT DFFSR_X1 CLK D Q RN SN VDD VSS
*.PININFO CLK:I D:I RN:I SN:I Q:O VDD:B VNW:B VPW:B VSS:B
mNM13 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM39 net5 rnb net4 VPW nch5 mr=1 l=600n w=220n nf=1
mM19 Q net2 VSS VPW nch5 mr=1 l=600n w=1.15u nf=1
mM38 net4 SN VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM17 net1 clkn net5 VPW nch5 mr=1 l=600n w=220n nf=1
mM25 net7 net10 net8 VPW nch5 mr=1 l=600n w=220n nf=1
mM31 net7 D net12 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM28 net12 clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM22 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM34 rnb RN VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM7 net9 SN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM32 net10 clkp net1 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM9 net2 net1 VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM10 net10 rnb net9 VPW nch5 mr=1 l=600n w=735n nf=1
mNM3 net10 net7 net9 VPW nch5 mr=1 l=600n w=735n nf=1
mM24 net8 clkp VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM42 net5 net2 net4 VPW nch5 mr=1 l=600n w=220n nf=1
mM29 net6 clkp VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM43 net5 net2 net3 VNW pch5 mr=1 l=500n w=220n nf=1
mM27 net13 clkn VDD VNW pch5 mr=1 l=500n w=220n nf=1
mPM13 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM16 net1 clkp net5 VNW pch5 mr=1 l=500n w=220n nf=1
mM35 rnb RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM26 net7 net10 net13 VNW pch5 mr=1 l=500n w=220n nf=1
mM23 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM40 net5 SN VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM33 net10 clkn net1 VNW pch5 mr=1 l=500n w=1.03u nf=1
mM18 Q net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM6 net10 SN VDD VNW pch5 mr=1 l=500n w=1.01u nf=1
mPM3 net10 net7 net11 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM11 net11 rnb VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM30 net7 D net6 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM41 net3 rnb VDD VNW pch5 mr=1 l=500n w=220n nf=1
mPM9 net2 net1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    EDFFR_X1
* View Name:    schematic
************************************************************************

.SUBCKT EDFFR_X1 CLK D E Q RN VDD VSS
*.PININFO CLK:I D:I E:I RN:I Q:O VDD:B VNW:B VPW:B VSS:B
mNM20 Q net2 VSS VPW nch5 mr=1 l=600n w=1.15u nf=1
mM22 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM16 net1 clkn VSS VPW nch5 mr=1 l=600n w=220n nf=1
mNM3 net11 D net12 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM17 net5 net6 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM13 net194 RN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM8 net10 E VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM5 net13 Q VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM4 net11 net10 net13 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM1 net2 net3 VSS VPW nch5 mr=1 l=600n w=780n nf=1
mNM2 net12 E VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM14 net7 net11 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM12 net5 clkp net3 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM9 net8 clkn net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM31 net9 clkp VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM30 net6 net5 net9 VPW nch5 mr=1 l=600n w=220n nf=1
mM12 net8 net7 net194 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM18 net3 net2 net1 VPW nch5 mr=1 l=600n w=220n nf=1
mNM15 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mPM20 Q net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM15 net7 net11 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM23 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM17 net14 clkp VDD VNW pch5 mr=1 l=500n w=300n nf=1
mPM5 net164 D VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM4 net164 E VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM2 net11 net10 net164 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM3 net11 Q net164 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM19 net3 net2 net14 VNW pch5 mr=1 l=500n w=300n nf=1
mPM15 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM17 net5 net6 VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mPM1 net2 net3 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM12 net5 clkn net3 VNW pch5 mr=1 l=500n w=1.68u nf=1
mPM9 net8 clkp net6 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM9 net10 E VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM10 net8 net7 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM11 net8 RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM28 net4 clkn VDD VNW pch5 mr=1 l=500n w=300n nf=1
mM29 net6 net5 net4 VNW pch5 mr=1 l=500n w=300n nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    CLKGTP_X1
* View Name:    schematic
************************************************************************

.SUBCKT CLKGTP_X1 CLK E GCLK VDD VSS
*.PININFO CLK:I E:I GCLK:O VDD:B VNW:B VPW:B VSS:B
mM22 net1 net10 net11 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM21 net10 net8 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM19 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM13 GCLK net1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM23 net11 clkp VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM7 net2 clkp net4 VNW pch5 mr=1 l=500n w=500n nf=1
mM6 net4 net8 VDD VNW pch5 mr=1 l=500n w=500n nf=1
mM1 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM3 net2 clkn net3 VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM1 net8 net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM2 net3 E VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM20 net10 net8 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM11 net1 clkp VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM18 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM12 GCLK net1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM10 net1 net10 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM9 net2 clkn net7 VPW nch5 mr=1 l=600n w=220n nf=1
mM8 net7 net8 VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM5 net2 clkp net9 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM4 net9 E VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM0 net8 net2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    LATSR_X1
* View Name:    schematic
************************************************************************

.SUBCKT LATSR_X1 D E Q RN SN VDD VSS
*.PININFO D:I E:I RN:I SN:I Q:O VDD:B VNW:B VPW:B VSS:B
mM11 net8 net2 net4 VPW nch5 mr=1 l=600n w=220n nf=1
mM10 net4 en VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM18 net1 net2 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM21 net2 rnb net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM7 net6 SN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM29 en E VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM25 net8 D net5 VPW nch5 mr=1 l=600n w=1.21u nf=1
mNM3 net2 net8 net6 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 Q net1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM34 rnb RN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM16 enb en VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM20 net5 enb VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM13 net3 enb VDD VNW pch5 mr=1 l=500n w=500n nf=1
mM12 net8 net2 net3 VNW pch5 mr=1 l=500n w=500n nf=1
mPM3 net2 net8 net10 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM22 net10 rnb VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM6 net2 SN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mPM29 en E VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM19 net1 net2 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM31 net8 D net7 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM17 enb en VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM35 rnb RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM1 Q net1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM33 net7 en VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    SDFFSR_X1
* View Name:    schematic
************************************************************************

.SUBCKT SDFFSR_X1 CLK D Q RN SE SI SN VDD VSS
*.PININFO CLK:I D:I RN:I SE:I SI:I SN:I Q:O VDD:B VNW:B VPW:B VSS:B
mM9 net4 SEN net11 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM7 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.68u nf=1
mM48 SEN SE VDD VNW pch5 mr=1 l=500n w=1.68u nf=1
mM11 net4 SE net14 VNW pch5 mr=1 l=500n w=1.68u nf=1
mM51 net2 SN VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM10 net14 D VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM50 net2 net6 net16 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM61 net1 net8 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM64 Q net1 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM59 net2 clkn net8 VNW pch5 mr=1 l=500n w=1.68u nf=1
mM56 net6 net2 net15 VNW pch5 mr=1 l=500n w=220n nf=1
mM8 net11 SI VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM69 net5 net1 net10 VNW pch5 mr=1 l=500n w=220n nf=1
mM42 net6 clkp net4 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM46 rnb RN VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM49 net16 rnb VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM68 net10 rnb VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM67 net5 SN VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM55 net15 clkn VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM66 net8 clkp net5 VNW pch5 mr=1 l=500n w=220n nf=1
mM5 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM62 net1 net8 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM47 SEN SE VSS VPW nch5 mr=1 l=600n w=1.15u nf=1
mM53 net2 rnb net3 VPW nch5 mr=1 l=600n w=1.15u nf=1
mM6 clkp clkn VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM15 net13 D VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM52 net2 net6 net3 VPW nch5 mr=1 l=600n w=780n nf=1
mM41 net6 clkn net9 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM14 net7 SI VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM16 net9 SEN net13 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM60 net2 clkp net8 VPW nch5 mr=1 l=600n w=780n nf=1
mM63 Q net1 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM54 net3 SN VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM4 clkn CLK VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 net9 SE net7 VPW nch5 mr=1 l=600n w=1.15u nf=1
mM57 net6 net2 net17 VPW nch5 mr=1 l=600n w=220n nf=1
mM45 rnb RN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM58 net17 clkp VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM71 net5 rnb net12 VPW nch5 mr=1 l=600n w=220n nf=1
mM70 net5 net1 net12 VPW nch5 mr=1 l=600n w=220n nf=1
mM72 net12 SN VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM65 net8 clkn net5 VPW nch5 mr=1 l=600n w=220n nf=1
.ENDS

************************************************************************
* Library Name: prima_sc180bcd_5v_9t_sch
* Cell Name:    SEDFFSR_X1
* View Name:    schematic
************************************************************************

.SUBCKT SEDFFSR_X1 CLK D E Q RN SE SI SN VDD VSS
*.PININFO CLK:I D:I E:I RN:I SE:I SI:I SN:I Q:O VDD:B VNW:B VPW:B VSS:B
mNM9 net010 clkn net013 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM14 seb SE VSS VPW nch5 mr=1 l=600n w=1.15u nf=1
mNM12 net12 clkp net15 VPW nch5 mr=1 l=600n w=1.15u nf=1
mM61 net060 RN net017 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM48 net060 seb net010 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM37 net15 clkn net26 VPW nch5 mr=1 l=600n w=220n nf=1
mM24 Q net20 VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM35 net013 clkp net28 VPW nch5 mr=1 l=600n w=220n nf=1
mM42 net12 net013 VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM36 net26 net20 VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM8 eb E VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM12 net010 SE net059 VPW nch5 mr=1 l=600n w=1.15u nf=1
mM44 net20 net15 VSS VPW nch5 mr=1 l=600n w=860n nf=1
mM49 net017 Q net047 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM3 net049 D VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM39 clkp clkn VSS VPW nch5 mr=1 l=600n w=780n nf=1
mNM1 clkn CLK VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM32 net28 net12 VSS VPW nch5 mr=1 l=600n w=220n nf=1
mM1 snb SN VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM4 net060 snb VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM50 net047 eb VSS VPW nch5 mr=1 l=600n w=1.21u nf=1
mM0 net017 E net049 VPW nch5 mr=1 l=600n w=1.21u nf=1
mM11 net059 SI VSS VPW nch5 mr=1 l=600n w=780n nf=1
mM62 net058 SI VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mPM9 net010 clkp net013 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM40 net15 clkp net25 VNW pch5 mr=1 l=500n w=220n nf=1
mM33 net013 clkn net27 VNW pch5 mr=1 l=500n w=220n nf=1
mM15 seb SE VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM65 net048 eb net1 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM58 net010 seb net058 VNW pch5 mr=1 l=500n w=1.25u nf=1
mM43 net12 net013 VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM31 clkn CLK VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM38 clkp clkn VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM60 net046 E net1 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM64 net060 RN net1 VNW pch5 mr=1 l=500n w=1.31u nf=1
mPM1 net20 net15 VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM18 net1 snb VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM54 net060 D net048 VNW pch5 mr=1 l=500n w=1.74u nf=1
mM9 eb E VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
mM63 net060 SE net010 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM66 net060 Q net046 VNW pch5 mr=1 l=500n w=1.68u nf=1
mPM12 net12 clkn net15 VNW pch5 mr=1 l=500n w=1.31u nf=1
mM41 net25 net20 VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM34 net27 net12 VDD VNW pch5 mr=1 l=500n w=220n nf=1
mM2 snb SN VDD VNW pch5 mr=1 l=500n w=1.31u nf=1
mM45 Q net20 VDD VNW pch5 mr=1 l=500n w=1.74u nf=1
.ENDS

