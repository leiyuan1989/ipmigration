*clk
.SUBCKT CLK1 CK VDD VSS C CN 
PM1 CN   CK  VDD VDD pmos l=1 w=1 n=1 ro=2 co=1
PM2 VDD  CN  C   VDD pmos l=1 w=1 n=1 ro=2 co=2
NM1 CN   CK  VSS VSS nmos l=1 w=1 n=1 ro=5 co=1
NM2 VSS  CN  C   VSS nmos l=1 w=1 n=1 ro=5 co=2  
.ends CLK1


.SUBCKT CLK2 CK VDD VSS C CN
PM1 nck   CK  VDD VDD pmos l=1 w=1 n=1 ro=1 co=1
NM1 nck   CK  VSS VSS nmos l=1 w=1 n=1 ro=1 co=1
PM2 VDD  nck  C   VDD pmos l=1 w=1 n=1 ro=1 co=2
NM2 VSS  nck  C   VSS nmos l=1 w=1 n=1 ro=1 co=2  
PM3 VDD  CK  net1 VDD pmos l=1 w=1 n=1 ro=1 co=3
NM3 VSS  CK  CN   VSS nmos l=1 w=1 n=1 ro=1 co=3
PM4 net1 C   CN   VDD pmos l=1 w=1 n=1 ro=1 co=4
.ends CLK2


******************INV************************

.SUBCKT INV IN1 VDD VSS OUT1
PM1 VDD  IN1  OUT1 VDD pmos l=1 w=1 n=1 ro=5 co=1
NM1 VSS  IN1  OUT1 VSS nmos l=1 w=1 n=1 ro=2 co=1
.ends INV



******************Logic 2************************
*Logic can be used to match clockgate output, D0 D1 and ...
.SUBCKT LOGIC2_AND2 IN1 IN2 VDD VSS OUT1
pmos_1 VDD  IN1  net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
nmos_1 net1 IN1  net2 VSS nmos l=1 w=1 n=1 ro=1 co=1
pmos_2 net1 IN2  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=2
nmos_2 net2 IN2  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=2
pmos_3 VDD  net1  OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=3
nmos_3 VSS  net1  OUT1  VSS nmos l=1 w=1 n=1 ro=1 co=3
.ends LOGIC2_AND2

.SUBCKT LOGIC2_AND2_2 IN1 IN2 VDD VSS OUT1
pmos_1 VDD  IN1  net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
pmos_2 net1 IN2  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=3
nmos_1 net1 IN1  net2 VSS nmos l=1 w=1 n=1 ro=1 co=1
nmos_3 net1 IN1  net3 VSS nmos l=1 w=1 n=1 ro=1 co=2
nmos_2 net2 IN2  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=3
nmos_4 net3 IN2  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=4
pmos_5 VDD  net1  OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=3
nmos_5 VSS  net1  OUT1  VSS nmos l=1 w=1 n=1 ro=1 co=3
.ends LOGIC2_AND2_2

.SUBCKT LOGIC2_OR2 IN1 IN2 VDD VSS OUT1
pmos_1 net1  IN1  net2 VDD pmos l=1 w=1 n=1 ro=1 co=1
nmos_1 VSS   IN1  net1 VSS nmos l=1 w=1 n=1 ro=1 co=1
pmos_2 net2  IN2  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=2
nmos_2 net1  IN2  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=2
pmos_3 VDD  net1  OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=3
nmos_3 VSS  net1  OUT1  VSS nmos l=1 w=1 n=1 ro=1 co=3
.ends LOGIC2_OR2

.SUBCKT LOGIC2_NAND2 IN1 IN2 VDD VSS OUT1
pmos_1 OUT1 IN2  VDD VDD pmos l=1 w=1 n=1 ro=1 co=1
nmos_1 OUT1 IN2  net1  VSS nmos l=1 w=1 n=1 ro=1 co=1
pmos_2 VDD  IN1  OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=2
nmos_2 net1 IN1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=2  
.ends LOGIC2_NAND2

.SUBCKT LOGIC2_NOR2 IN1 IN2 VDD VSS OUT1
PM1 VDD  IN1  net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
NM1 VSS  IN1  OUT1  VSS nmos l=1 w=1 n=1 ro=1 co=1
PM2 net1 IN2  OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=2
NM2 OUT1 IN2  VSS  VSS nmos l=1 w=1 n=1  ro=1 co=2
.ends LOGIC2_NOR2

******************Logic 3************************

******************Logic 4************************

******************Logic 5************************




******************Fully Cross************************
*FCROSS can be used to match D with E or CN/C with D
.SUBCKT FCROSS_1 D E E_N D1 VDD VSS OUT1 OUT2 
PM1 VDD   E_N net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 net1  D   OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 OUT1  D1  net2 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM4 net2  E   VDD  VDD pmos l=1 w=1 n=1 ro=1 co=4
NM1 VSS   E   net3 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 net3  D   OUT2 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 OUT2  D1  net4 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM4 net4  E_N VSS  VSS nmos l=1 w=1 n=1 ro=1 co=4
.ends FCROSS_1

.SUBCKT FCROSS_2  D E E_N D1 VDD VSS OUT1
PM1 VDD   E_N net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 net1  D   OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 OUT1  D1  net2 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM4 net2  E   VDD  VDD pmos l=1 w=1 n=1 ro=1 co=4
NM1 VSS   E   net3 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 net3  D   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 OUT1  D1  net4 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM4 net4  E_N VSS  VSS nmos l=1 w=1 n=1 ro=1 co=4
.ends FCROSS_2

.SUBCKT FCROSS_3  D E E_N D1 VDD VSS OUT1 OUT2
PM1 VDD   D   net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 net1  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM4 net2  D1  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=4

NM1 VSS   D   net3 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 net3  E   OUT2 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 OUT2  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM4 net4  D1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=4
.ends FCROSS_3

.SUBCKT FCROSS_4  D E E_N D1 VDD VSS OUT1
PM1 VDD   D   net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 net1  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM4 net2  D1  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=4
NM1 VSS   D   net3 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 net3  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM4 net4  D1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=4
.ends FCROSS_4

*2 D with 2 EN
.SUBCKT FCROSS_4_2  D E E_N D1 VDD VSS OUT1
PM0 OUT1  E_N net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM1 net1  D   VDD  VDD pmos l=1 w=1 n=1 ro=1 co=2
PM2 VDD   D   net2 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM3 net2  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=4
PM4 OUT1  E   net3 VDD pmos l=1 w=1 n=1 ro=1 co=5
PM5 net3  D1  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=6
NM0 OUT1  E   net4 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM1 net4  D   VSS  VSS nmos l=1 w=1 n=1 ro=1 co=2
NM2 VSS   D   net5 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM3 net5  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=4
NM4 OUT1  E_N net6 VSS nmos l=1 w=1 n=1 ro=1 co=5
NM5 net6  D1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=6
.ends FCROSS_4_2




******************PCROSS without D********************************
.SUBCKT PCROSS_1 IN1 IN2 D1 E_N E OUT1 VDD VSS 
PM1 IN1   E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 net2  D1  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=3
NM1 IN2   E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 net4  D1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=3
.ends PCROSS_1


.SUBCKT PCROSS_2 IN1 D1 E_N E OUT1 VDD VSS 
PM1 IN1   E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 net2  D1  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=3
NM1 IN1   E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 net4  D1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=3
.ends PCROSS_2







******************Asynchronous************************
*Cross with RN and SN
.SUBCKT FRSCROSS_1  D E E_N D1 RN NSN VDD VSS OUT1
PM1 nsnp  D   net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 net1  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM4 net2  D1  nsnp VDD pmos l=1 w=1 n=1 ro=1 co=4
NM1 rng   D   net3 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 net3  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM4 net4  D1  rng  VSS nmos l=1 w=1 n=1 ro=1 co=4

PM5 OUT1  RN  nsnp VDD pmos l=1 w=1 n=1 ro=1 co=6
NM5 rng   RN  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=6

PM6 nsnp  NSN VDD  VDD pmos l=1 w=1 n=1 ro=1 co=8
NM6 OUT1  NSN VSS  VSS nmos l=1 w=1 n=1 ro=1 co=8
.ends FRSCROSS_1

*net3 changed to net1
.SUBCKT FRSCROSS_1_2  D E E_N D1 RN NSN VDD VSS OUT1
PM1 nsnp  D   net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 net1  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM4 net2  D1  nsnp VDD pmos l=1 w=1 n=1 ro=1 co=4
NM1 rng   D   net1 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 net1  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM4 net4  D1  rng  VSS nmos l=1 w=1 n=1 ro=1 co=4

PM5 OUT1  RN  nsnp VDD pmos l=1 w=1 n=1 ro=1 co=6
NM5 rng   RN  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=6

PM6 nsnp  NSN VDD  VDD pmos l=1 w=1 n=1 ro=1 co=8
NM6 OUT1  NSN VSS  VSS nmos l=1 w=1 n=1 ro=1 co=8
.ends FRSCROSS_1_2


*Cross with RN 
.SUBCKT FRCROSS_1  D E E_N D1 RN VDD VSS OUT1
PM1 VDD   D   net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 net1  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM4 net2  D1  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=4
NM1 rng   D   net3 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 net3  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM4 net4  D1  rng  VSS nmos l=1 w=1 n=1 ro=1 co=4

PM5 OUT1  RN  VDD VDD pmos l=1 w=1 n=1 ro=1 co=6
NM5 rng   RN  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=6
.ends FRCROSS_1

*net3 changed to net1
.SUBCKT FRCROSS_1_2  D E E_N D1 RN VDD VSS OUT1
PM1 VDD   D   net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 net1  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM4 net2  D1  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=4
NM1 rng   D   net1 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 net1  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM4 net4  D1  rng  VSS nmos l=1 w=1 n=1 ro=1 co=4

PM5 OUT1  RN  VDD VDD pmos l=1 w=1 n=1 ro=1 co=6
NM5 rng   RN  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=6
.ends FRCROSS_1_2

*2 rng, maybe for layout, c110:LACHB0
.SUBCKT FRCROSS_1_3  D E E_N D1 RN VDD VSS OUT1
PM1 VDD   D   net1 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM2 net1  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM3 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=4
PM4 net2  D1  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=5

NM0 VSS   RN  rng1 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM1 rng1  D   net1 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM2 net1  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM3 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=4
NM4 net4  D1  rng2 VSS nmos l=1 w=1 n=1 ro=1 co=5

PM5 OUT1  RN  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=7
NM5 rng2  RN  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=7
.ends FRCROSS_1_3

*Cross with SN 
.SUBCKT FSCROSS_1  D E E_N D1 NSN VDD VSS OUT1
PM0 VDD   NSN nsnp VDD pmos l=1 w=1 n=1 ro=1 co=1
NM0 VSS   NSN OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=1

PM1 nsnp  D   net1 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM2 net1  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=4
PM3 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=5
PM4 net2  D1  nsnp VDD pmos l=1 w=1 n=1 ro=1 co=6
NM1 VSS   D   net3 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM2 net3  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=4
NM3 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=5
NM4 net4  D1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=6
.ends FSCROSS_1

*net3 changed to net1
.SUBCKT FSCROSS_1_2  D E E_N D1 NSN VDD VSS OUT1
PM0 VDD   NSN nsnp VDD pmos l=1 w=1 n=1 ro=1 co=1
NM0 VSS   NSN OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=1

PM1 nsnp  D   net1 VDD pmos l=1 w=1 n=1 ro=1 co=3
PM2 net1  E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=4
PM3 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=5
PM4 net2  D1  nsnp VDD pmos l=1 w=1 n=1 ro=1 co=6
NM1 VSS   D   net1 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM2 net1  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=4
NM3 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=5
NM4 net4  D1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=6
.ends FSCROSS_1_2

*2 nsnp, maybe for layout, c110:LAPHB0
.SUBCKT FSCROSS_1_3  D E E_N D1 NSN VDD VSS OUT1
PM0 VDD   NSN nsnp1 VDD pmos l=1 w=1 n=1 ro=1 co=1
NM0 VSS   NSN OUT1  VSS nmos l=1 w=1 n=1 ro=1 co=1

PM1 nsnp1 D   net1  VDD pmos l=1 w=1 n=1 ro=1 co=3
PM2 net1  E_N OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=4
PM3 OUT1  E   net2  VDD pmos l=1 w=1 n=1 ro=1 co=5
PM4 net2  D1  nsnp2 VDD pmos l=1 w=1 n=1 ro=1 co=6
PM5 nsnp2 NSN VDD   VDD pmos l=1 w=1 n=1 ro=1 co=7

NM1 VSS   D   net1 VSS nmos l=1 w=1 n=1 ro=1 co=3
NM2 net1  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=4
NM3 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=5
NM4 net4  D1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=6
.ends FSCROSS_1_3

*2 nsnp1 and 1 nsnp2,  c110:LAPLB3
.SUBCKT FSCROSS_1_3_2  D E E_N D1 NSN VDD VSS OUT1
PM1 net1  D   nsnp1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 nsnp1 NSN VDD   VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 VDD   NSN nsnp2 VDD pmos l=1 w=1 n=1 ro=1 co=3
NM1 VSS   NSN OUT1  VSS nmos l=1 w=1 n=1 ro=1 co=3

PM4 nsnp2 D   net1  VDD pmos l=1 w=1 n=1 ro=1 co=5
PM5 net1  E_N OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=6
PM6 OUT1  E   net2  VDD pmos l=1 w=1 n=1 ro=1 co=7
PM7 net2  D1  nsnp3 VDD pmos l=1 w=1 n=1 ro=1 co=8
PM8 nsnp3 NSN VDD   VDD pmos l=1 w=1 n=1 ro=1 co=9

NM2 VSS   D   net1 VSS nmos l=1 w=1 n=1 ro=1 co=5
NM3 net1  E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=6
NM4 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=7
NM5 net4  D1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=8
.ends FSCROSS_1_3_2





*
.SUBCKT PRCROSS_1 IN1 IN2 RN D1 E_N E OUT1 VDD VSS 
PM1 IN1   E_N OUT1 VDD pmos l=1 w=1 n=1 ro=1 co=1
PM2 OUT1  E   net2 VDD pmos l=1 w=1 n=1 ro=1 co=2
PM3 net2  D1  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=3
NM1 IN1   E   OUT1 VSS nmos l=1 w=1 n=1 ro=1 co=1
NM2 OUT1  E_N net4 VSS nmos l=1 w=1 n=1 ro=1 co=2
NM3 net4  D1  net5  VSS nmos l=1 w=1 n=1 ro=1 co=3
NM4 net5  RN  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=3
.ends PRCROSS_1












******************backtrack********************************
.SUBCKT BACKTRACK3_1  IN1 IN2 IN3 VDD VSS OUT1
PM1 VDD  IN1  NET3 VDD pmos  l=1 w=1 n=1 ro=1 co=1
PM2 NET3 IN2  OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=2
PM3 OUT1 IN3  VDD  VDD pmos  l=1 w=1 n=1 ro=1 co=3

NM1 NET4 IN1  OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=1
NM2 OUT1 IN2  NET4 VSS nmos  l=1 w=1 n=1 ro=1 co=2
NM3 NET4 IN3  VSS  VSS nmos  l=1 w=1 n=1 ro=1 co=3
.ends BACKTRACK3_1

.SUBCKT BACKTRACK3_2  IN1 IN2 IN3 VDD VSS OUT1
PM1 VDD  IN2 NET1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
PM2 NET1 IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=2
NM1 VSS  IN3 NET2 VSS nmos  l=1 w=1 n=1 ro=1 co=1
NM2 NET2 IN1 OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK3_2


*pull
.SUBCKT BACKTRACK3_3  IN1 IN2 IN3 VDD VSS OUT1
PM1 VDD  IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
PM2 IN1  IN2 VDD VDD pmos  l=1 w=1 n=1 ro=1 co=2
NM1 VSS  IN1 OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=2
NM2 IN1  IN3 VSS VSS nmos  l=1 w=1 n=1 ro=1 co=1
.ends BACKTRACK3_3

.SUBCKT BACKTRACK3_3_2  IN1 IN2 IN3 VDD VSS OUT1
PM1 VDD  IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
PM2 IN1 IN2 PDD  VDD pmos  l=1 w=1 n=1 ro=1 co=2
NM1 VSS  IN1 OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=1
NM2 IN1 IN3 VSS  VSS nmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK3_3_2

.SUBCKT BACKTRACK3_3_3  IN1 IN2 IN3 VDD VSS OUT1
PM1 VDD  IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
PM2 IN1 IN2 VDD  VDD pmos  l=1 w=1 n=1 ro=1 co=2
NM1 VSS  IN1 OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=1
NM2 IN1 IN3 PSS  VSS nmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK3_3_3

.SUBCKT BACKTRACK3_3_4  IN1 IN2 IN3 VDD VSS OUT1
PM1 VDD  IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
PM2 IN1 IN2 PDD  VDD pmos  l=1 w=1 n=1 ro=1 co=2
NM1 VSS  IN1 OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=1
NM2 IN1 IN3 PSS  VSS nmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK3_3_4


.SUBCKT BACKTRACK2_1  IN1 IN2 VDD VSS OUT1
PM1 VDD  IN2 NET1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
PM2 NET1 IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=2
NM2 VSS IN1 OUT1  VSS nmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK2_1

.SUBCKT BACKTRACK2_2  IN1 IN2 VDD VSS OUT1
PM1 VDD  IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
NM1 OUT1 IN1 NET1 VSS nmos  l=1 w=1 n=1 ro=1 co=2
NM2 NET1 IN2 VSS  VSS nmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK2_2



*pull
.SUBCKT BACKTRACK2_3  IN1 IN2  VDD VSS OUT1
PM1 VDD  IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
NM1 VSS  IN1 OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=1
PM2 IN1  IN2 VDD  VDD pmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK2_3

.SUBCKT BACKTRACK2_3_2  IN1 IN2  VDD VSS OUT1
PM1 VDD  IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
NM1 VSS  IN1 OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=1
PM2 IN1  IN2 PDD  VDD pmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK2_3_2

.SUBCKT BACKTRACK2_3_3  IN1 IN2  VDD VSS OUT1
PM1 VDD  IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
NM1 VSS  IN1 OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=1
NM2 IN1  IN2 VSS  VSS nmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK2_3_3

.SUBCKT BACKTRACK2_3_4  IN1 IN2  VDD VSS OUT1
PM1 VDD  IN1 OUT1 VDD pmos  l=1 w=1 n=1 ro=1 co=1
NM1 VSS  IN1 OUT1 VSS nmos  l=1 w=1 n=1 ro=1 co=1
NM2 IN1  IN2 PSS  VSS nmos  l=1 w=1 n=1 ro=1 co=2
.ends BACKTRACK2_3_4




