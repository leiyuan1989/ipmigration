* ---------------------------------------------------------------------------- 
* 
*     library Calibre-based CDL file 
* 
*     Date: Jan 31, 2012 7:10:22 PM IST 
* 
*     CellBuilder version 4.0.1 -- built on Nov 11, 2011 
*     Copyright (c) 2002-2011 ARM, Inc. 
*     The confidential and proprietary information contained in this file 
*     may only be used by a person authorised under and to the extent 
*     permitted by a subsisting licensing agreement from ARM Limited. 
*      
*     (C) COPYRIGHT 2004-2012 ARM Limited. 
*     ALL RIGHTS RESERVED 
*      
*     This entire notice must be reproduced on all copies of this file 
*     and copies of this file may only be made by a person if such person 
*     is permitted to do so under the terms of a subsisting license 
*     agreement from ARM Limited. 
* 
* ----------------------------------------------------------------------------

*.SCALE METER
*.OPTION SCALE 1e-6

.SUBCKT ADDFHX1MTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=130n w=530n
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=270n
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=6.3e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.9e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=6.3e-07
mXI5_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=3.9e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI11_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=3.7e-07
mXI12_MXNOE con xorab cin VPW n12 l=1.3e-07 w=3.7e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=3.7e-07
mXI10_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=3.7e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=7.7e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=7.7e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=7.7e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=5.8e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=7.7e-07
mXI5_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=6.8e-07
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI11_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=4.6e-07
mXI12_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=4.6e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=4.6e-07
mXI10_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=4.6e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT ADDFHX2MTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI15_MXNA1_2 ba na2 VSS VPW n12 l=1.3e-07 w=6e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=5.2e-07
mXI3_MXNOE_2 xnorab B ba VPW n12 l=1.3e-07 w=5.2e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNOE_2 xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=3.9e-07
mXI4_MXNOE_2 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI4_MXNOE_3 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI5_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=9.3e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI6_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI11_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=6.1e-07
mXI12_MXNOE con xorab cin VPW n12 l=1.3e-07 w=5.4e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI9_MXNOE_2 sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI10_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=5.5e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI7_MXNA1_2 cin CI VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI14_MXNA1_2 CO con VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI15_MXPA1_2 ba na2 VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=6.3e-07
mXI3_MXPOEN_2 xnorab nb ba VNW p12 l=1.3e-07 w=6.3e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPOEN_2 xnorab B na VNW p12 l=1.3e-07 w=5e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=6.3e-07
mXI4_MXPOEN_2 xorab nb na VNW p12 l=1.3e-07 w=6.3e-07
mXI5_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=1.22e-06
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI11_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=3.7e-07
mXI11_MXPOEN_2 con xorab nb VNW p12 l=1.3e-07 w=4.4e-07
mXI12_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=6e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=7.4e-07
mXI10_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=7.4e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=9.8e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI13_MXPA1_2 S sumn VDD VNW p12 l=1.3e-07 w=4.4e-07
.ends


.SUBCKT ADDFHX4MTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=8.6e-07
mXI15_MXNA1_2 ba na2 VSS VPW n12 l=1.3e-07 w=8.6e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=8.6e-07
mXI3_MXNOE_2 xnorab B ba VPW n12 l=1.3e-07 w=6.7e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNOE_2 xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=3.9e-07
mXI4_MXNOE_2 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI4_MXNOE_3 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI5_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=9.3e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=9.8e-07
mXI6_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=9.8e-07
mXI6_MXNA1_3 nb B VSS VPW n12 l=1.3e-07 w=9.8e-07
mXI11_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=6.1e-07
mXI12_MXNOE con xorab cin VPW n12 l=1.3e-07 w=5.4e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI9_MXNOE_2 sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI10_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=5.5e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI8_MXNA1_2 cib cin VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1_2 cin CI VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1_3 cin CI VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI14_MXNA1_2 CO con VSS VPW n12 l=1.3e-07 w=7e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI13_MXNA1_2 S sumn VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI15_MXPA1_2 ba na2 VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI15_MXPA1_3 ba na2 VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=6.7e-07
mXI3_MXPOEN_2 xnorab nb ba VNW p12 l=1.3e-07 w=6.7e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=5.5e-07
mXI1_MXPOEN_2 xnorab B na VNW p12 l=1.3e-07 w=5.5e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=8.6e-07
mXI4_MXPOEN_2 xorab nb na VNW p12 l=1.3e-07 w=1.01e-06
mXI5_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=1.2e-06
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI6_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_5 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_6 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_7 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI11_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=5.2e-07
mXI11_MXPOEN_2 con xorab nb VNW p12 l=1.3e-07 w=5.2e-07
mXI12_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=6e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=7.4e-07
mXI10_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=9.8e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=9.8e-07
mXI8_MXPA1_2 cib cin VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=9.8e-07
mXI7_MXPA1_2 cin CI VDD VNW p12 l=1.3e-07 w=9.8e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI14_MXPA1_2 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1_2 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT ADDFHX8MTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_4 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_5 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI2_MXNA1_2 na2 A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI2_MXNA1_3 na2 A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_2 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_3 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_4 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_5 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI15_MXNA1_6 ba na2 VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=6.9e-07
mXI3_MXNOE_2 xnorab B ba VPW n12 l=1.3e-07 w=6.7e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNOE_2 xnorab nb na VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=3.7e-07
mXI4_MXNOE_2 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI4_MXNOE_3 xorab B na VPW n12 l=1.3e-07 w=3.2e-07
mXI5_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=6.7e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=9.9e-07
mXI6_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=9.9e-07
mXI11_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=6.1e-07
mXI12_MXNOE con xorab cin VPW n12 l=1.3e-07 w=5.4e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI9_MXNOE_2 sumn xnorab cin VPW n12 l=1.3e-07 w=2.4e-07
mXI10_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=5.5e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=5.5e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI7_MXNA1_2 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI7_MXNA1_3 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI7_MXNA1_4 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI7_MXNA1_5 cin CI VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI14_MXNA1_2 CO con VSS VPW n12 l=1.3e-07 w=6.7e-07
mXI14_MXNA1_3 CO con VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI14_MXNA1_4 CO con VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNA1_2 S sumn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNA1_3 S sumn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI13_MXNA1_4 S sumn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_4 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_5 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_6 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI2_MXPA1_2 na2 A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI2_MXPA1_3 na2 A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_2 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_3 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_4 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_5 ba na2 VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI15_MXPA1_6 ba na2 VDD VNW p12 l=1.3e-07 w=6.7e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=6.7e-07
mXI3_MXPOEN_2 xnorab nb ba VNW p12 l=1.3e-07 w=6.7e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=5.5e-07
mXI1_MXPOEN_2 xnorab B na VNW p12 l=1.3e-07 w=5.5e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=8.6e-07
mXI4_MXPOEN_2 xorab nb na VNW p12 l=1.3e-07 w=1.01e-06
mXI5_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=1.22e-06
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI11_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=5.3e-07
mXI11_MXPOEN_2 con xorab nb VNW p12 l=1.3e-07 w=5.3e-07
mXI12_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=6e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=9.8e-07
mXI10_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=9.8e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI7_MXPA1_2 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI7_MXPA1_3 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI7_MXPA1_4 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI7_MXPA1_5 cin CI VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI14_MXPA1_2 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI14_MXPA1_3 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI14_MXPA1_4 CO con VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI13_MXPA1_2 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1_3 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI13_MXPA1_4 S sumn VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT ADDFHXLMTR CO S VDD VNW VPW VSS A B CI
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI2_MXNA1 na2 A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 ba na2 VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI3_MXNOE xnorab B ba VPW n12 l=1.3e-07 w=3.5e-07
mXI1_MXNOE xnorab nb na VPW n12 l=1.3e-07 w=3.5e-07
mXI4_MXNOE xorab B na VPW n12 l=1.3e-07 w=3.5e-07
mXI25_MXNOE xorab nb ba VPW n12 l=1.3e-07 w=3.5e-07
mXI6_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI23_MXNOE con xnorab nb VPW n12 l=1.3e-07 w=2.1e-07
mXI24_MXNOE con xorab cin VPW n12 l=1.3e-07 w=2.1e-07
mXI9_MXNOE sumn xnorab cin VPW n12 l=1.3e-07 w=2.1e-07
mXI22_MXNOE sumn xorab cib VPW n12 l=1.3e-07 w=2.1e-07
mXI8_MXNA1 cib cin VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI7_MXNA1 cin CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI14_MXNA1 CO con VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 S sumn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=4.3e-07
mXI2_MXPA1 na2 A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 ba na2 VDD VNW p12 l=1.3e-07 w=4.3e-07
mXI3_MXPOEN xnorab nb ba VNW p12 l=1.3e-07 w=4.3e-07
mXI1_MXPOEN xnorab B na VNW p12 l=1.3e-07 w=4.3e-07
mXI4_MXPOEN xorab nb na VNW p12 l=1.3e-07 w=4.3e-07
mXI25_MXPOEN xorab B ba VNW p12 l=1.3e-07 w=4.3e-07
mXI6_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI6_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=3e-07
mXI23_MXPOEN con xorab nb VNW p12 l=1.3e-07 w=2.5e-07
mXI24_MXPOEN con xnorab cin VNW p12 l=1.3e-07 w=2.5e-07
mXI9_MXPOEN sumn xorab cin VNW p12 l=1.3e-07 w=2.5e-07
mXI22_MXPOEN sumn xnorab cib VNW p12 l=1.3e-07 w=2.5e-07
mXI8_MXPA1 cib cin VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI7_MXPA1 cin CI VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI14_MXPA1 CO con VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI13_MXPA1 S sumn VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT ADDFX1MTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT ADDFX2MTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.5e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.8e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDFX4MTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.5e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDFX8MTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 CO nco VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_3 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 S ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.5e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 S ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDFXLMTR CO S VDD VNW VPW VSS A B CI
mX_g4_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5e-07
MXN0 xo na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE xo bb na VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE xn nb na VPW n12 l=1.3e-07 w=3e-07
MX_t8 xn na nb VPW n12 l=1.3e-07 w=4.5e-07
mXI7_MXNOE nco xn nb VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE nci xo nco VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nci CI VSS VPW n12 l=1.3e-07 w=3e-07
mXI10_MXNOE ns CI xo VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE ns nci xn VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 S ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t9 bb na xn VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN xn bb na VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN xo nb na VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nb na xo VNW p12 l=1.3e-07 w=5.5e-07
mXI7_MXPOEN nco xo nb VNW p12 l=1.3e-07 w=3.7e-07
mXI8_MXPOEN nci xn nco VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nci CI VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI10_MXPOEN ns nci xo VNW p12 l=1.3e-07 w=3.7e-07
mXI9_MXPOEN ns CI xn VNW p12 l=1.3e-07 w=3.7e-07
mX_g1_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 S ns VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT ADDHX1MTR CO S VDD VNW VPW VSS A B
mX_g3_MXNA1 ba na VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNOE S nb ba VPW n12 l=1.3e-07 w=3e-07
mXI9_MXNOE S B na VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 na A VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g2_MXNA2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g2_MXNA1 nco B X_g2_n1 VPW n12 l=1.3e-07 w=2.3e-07
mX_g0_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 ba na VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPOEN S B ba VNW p12 l=1.3e-07 w=3.8e-07
mXI9_MXPOEN S nb na VNW p12 l=1.3e-07 w=3.8e-07
mX_g4_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g2_MXPA2 nco A VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 nco B VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT ADDHX2MTR CO S VDD VNW VPW VSS A B
mX_g1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g3_MXNA1 ba na VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI10_MXNOE S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE S B na VPW n12 l=1.3e-07 w=6e-07
mX_g2_MXNA1 nco B X_g2_n1 VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g4_MXNA1 na A VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g4_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g4_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=5.9e-07
mX_g0_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g3_MXPA1 ba na VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI10_MXPOEN S B ba VNW p12 l=1.3e-07 w=7.5e-07
mXI9_MXPOEN S nb na VNW p12 l=1.3e-07 w=7.5e-07
mX_g2_MXPA1 nco B VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA2 nco A VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g4_MXPA1 na A VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g4_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDHX4MTR CO S VDD VNW VPW VSS A B
mX_g3_MXNA1 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI10_MXNOE S nb ba VPW n12 l=1.3e-07 w=5.9e-07
mXI10_MXNOE_2 S nb ba VPW n12 l=1.3e-07 w=5.9e-07
mXI9_MXNOE S B na VPW n12 l=1.3e-07 w=5.9e-07
mXI9_MXNOE_2 S B na VPW n12 l=1.3e-07 w=5.9e-07
mX_g2_MXNA1 nco B X_g2_n1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1_4 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1_5 na A VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g0_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI10_MXPOEN S B ba VNW p12 l=1.3e-07 w=7.6e-07
mXI10_MXPOEN_2 S B ba VNW p12 l=1.3e-07 w=7.6e-07
mXI9_MXPOEN S nb na VNW p12 l=1.3e-07 w=7.6e-07
mXI9_MXPOEN_2 S nb na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 nco B VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g2_MXPA2 nco A VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g4_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g4_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g4_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g4_MXPA1_4 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g4_MXPA1_5 na A VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g0_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT ADDHX8MTR CO S VDD VNW VPW VSS A B
mX_g3_MXNA1 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_2 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_3 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXNA1_4 ba na VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=5.7e-07
mX_g1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI10_MXNOE S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI10_MXNOE_2 S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI10_MXNOE_3 S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI10_MXNOE_4 S nb ba VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE S B na VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE_2 S B na VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE_3 S B na VPW n12 l=1.3e-07 w=6e-07
mXI9_MXNOE_4 S B na VPW n12 l=1.3e-07 w=6e-07
mX_g2_MXNA1 nco B X_g2_n1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nco B X_g2_n1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA2_2 X_g2_n1 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g4_MXNA1 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_3 na A VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g4_MXNA1_4 na A VSS VPW n12 l=1.3e-07 w=7e-07
mX_g4_MXNA1_5 na A VSS VPW n12 l=1.3e-07 w=7e-07
mX_g4_MXNA1_6 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_7 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_8 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_9 na A VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g4_MXNA1_10 na A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 CO nco VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_2 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 ba na VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI10_MXPOEN S B ba VNW p12 l=1.3e-07 w=6.1e-07
mXI10_MXPOEN_2 S B ba VNW p12 l=1.3e-07 w=6.1e-07
mXI10_MXPOEN_3 S B ba VNW p12 l=1.3e-07 w=6.1e-07
mXI10_MXPOEN_4 S B ba VNW p12 l=1.3e-07 w=6.1e-07
mXI9_MXPOEN S nb na VNW p12 l=1.3e-07 w=5.8e-07
mXI9_MXPOEN_2 S nb na VNW p12 l=1.3e-07 w=8.2e-07
mXI9_MXPOEN_3 S nb na VNW p12 l=1.3e-07 w=8.2e-07
mXI9_MXPOEN_4 S nb na VNW p12 l=1.3e-07 w=8.2e-07
mX_g2_MXPA1 nco B VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g2_MXPA1_2 nco B VDD VNW p12 l=1.3e-07 w=7.5e-07
mX_g2_MXPA2 nco A VDD VNW p12 l=1.3e-07 w=7.5e-07
mX_g2_MXPA2_2 nco A VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g4_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_3 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_4 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_5 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_6 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_7 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_8 na A VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g4_MXPA1_9 na A VDD VNW p12 l=1.3e-07 w=8.6e-07
mX_g4_MXPA1_10 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 CO nco VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND2X12MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA2_2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA2_3 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1_2 ny A XI0_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1_3 ny A XI0_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=6e-07
.ends


.SUBCKT AND2X1MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.1e-07
.ends


.SUBCKT AND2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=5.9e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND3X12MTR Y VDD VNW VPW VSS A B C
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A XI0_n2__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n2__3 B XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n1__3 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA3_3 ny C VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=5.9e-07
.ends


.SUBCKT AND3X1MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AND3X2MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=4.5e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND3X4MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND3X6MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_2 ny A XI0_n2__2 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND3X8MTR Y VDD VNW VPW VSS A B C
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 ny A XI0_n2__2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 ny A XI0_n2__3 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_3 XI0_n2__3 B XI0_n1__3 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3_3 XI0_n1__3 C VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3_3 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
.ends


.SUBCKT AND3XLMTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AND4X12MTR Y VDD VNW VPW VSS A B C D
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 ny A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA4_2 ny D VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA4_3 ny D VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA4_4 ny D VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA3_3 ny C VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA3_4 ny C VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA2_4 ny B VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=5e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=5e-07
.ends


.SUBCKT AND4X1MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=3.3e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=3.3e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=3.3e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AND4X2MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND4X4MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4_2 XI0_n1__2 D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3_2 XI0_n2__2 C XI0_n1__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_2 XI0_n3__2 B XI0_n2__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 ny A XI0_n3__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA4_2 ny D VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND4X6MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=6.5e-07
mXI0_MXNA1_2 ny A XI0_n3 VPW n12 l=1.3e-07 w=6.5e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA4_2 ny D VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AND4X8MTR Y VDD VNW VPW VSS A B C D
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 ny A XI0_n3 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 ny A XI0_n3 VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA4_2 ny D VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA4_3 ny D VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3_2 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA3_3 ny C VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
.ends


.SUBCKT AND4XLMTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA1 ny A XI0_n3 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA3 ny C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA4 ny D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends




.SUBCKT AO21X1MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AO21X2MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO21X4MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO21X8MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 ny A0 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 ny B0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO21XLMTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 ny A0 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 ny B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny B0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.4e-07
.ends


.SUBCKT AO22X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.1e-07
.ends


.SUBCKT AO22X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=4.4e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=4.4e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=4.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO22X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO22X8MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2_2 XI0_n1B__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 ny B0 XI0_n1B__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1A__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A0 XI0_n1A__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO22XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 ny B0 XI0_n1B VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 ny A0 XI0_n1A VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 ny A1 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AO2B2BX1MTR Y VDD VNW VPW VSS A0 A1N B0 B1N
mXI2_MXNA1 b1 B1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN6 net34 b1 VSS VPW n12 l=1.3e-07 w=2.3e-07
MXNB0 ny B0 net34 VPW n12 l=1.3e-07 w=2.3e-07
MXN4 ny A0 net40 VPW n12 l=1.3e-07 w=2.3e-07
MXN5 net40 a1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI2_MXPA1 b1 B1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net46 b1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXPB0 net46 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 ny A0 net46 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 ny a1 net46 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AO2B2BX2MTR Y VDD VNW VPW VSS A0 A1N B0 B1N
mXI2_MXNA1 b1 B1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN9 net34 b1 VSS VPW n12 l=1.3e-07 w=3.7e-07
MXNB0 ny B0 net34 VPW n12 l=1.3e-07 w=3.7e-07
MXN7 ny A0 net40 VPW n12 l=1.3e-07 w=3.7e-07
MXN8 net40 a1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 b1 B1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net46 b1 VDD VNW p12 l=1.3e-07 w=4.4e-07
MXPB0 net46 B0 VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP7 ny A0 net46 VNW p12 l=1.3e-07 w=4.4e-07
MXP9 ny a1 net46 VNW p12 l=1.3e-07 w=4.4e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO2B2BX4MTR Y VDD VNW VPW VSS A0 A1N B0 B1N
mXI2_MXNA1 b1 B1N VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN12 net34 b1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 ny B0 net34 VPW n12 l=1.3e-07 w=7.1e-07
MXN10 ny A0 net40 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 net40 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 b1 B1N VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP10 net46 b1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPB0 net46 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12 ny A0 net46 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 ny a1 net46 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO2B2BXLMTR Y VDD VNW VPW VSS A0 A1N B0 B1N
mXI2_MXNA1 b1 B1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN15 net34 b1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNB0 ny B0 net34 VPW n12 l=1.3e-07 w=1.8e-07
MXN13 ny A0 net40 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net40 a1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXPA1 b1 B1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 net46 b1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 net46 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 ny A0 net46 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 ny a1 net46 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AO2B2X1MTR Y VDD VNW VPW VSS A0 A1N B0 B1
MXN8 net051 B1 VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN5 ny B0 net051 VPW n12 l=1.3e-07 w=2.3e-07
MXN6 ny A0 net35 VPW n12 l=1.3e-07 w=2.3e-07
MXN7 net35 a1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP5 net41 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net41 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 ny A0 net41 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 ny a1 net41 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AO2B2X2MTR Y VDD VNW VPW VSS A0 A1N B0 B1
MXN12 net051 B1 VSS VPW n12 l=1.3e-07 w=3.7e-07
MXN13 ny B0 net051 VPW n12 l=1.3e-07 w=3.7e-07
MXN10 ny A0 net35 VPW n12 l=1.3e-07 w=3.7e-07
MXN11 net35 a1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP9 net41 B1 VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP10 net41 B0 VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP11 ny A0 net41 VNW p12 l=1.3e-07 w=4.4e-07
MXP12 ny a1 net41 VNW p12 l=1.3e-07 w=4.4e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO2B2X4MTR Y VDD VNW VPW VSS A0 A1N B0 B1
MXN2 net051 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 ny B0 net051 VPW n12 l=1.3e-07 w=7.1e-07
MXN0 ny A0 net35 VPW n12 l=1.3e-07 w=7.1e-07
MXN1 net35 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP14 net41 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 net41 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16 ny A0 net41 VNW p12 l=1.3e-07 w=8.7e-07
MXP17 ny a1 net41 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AO2B2XLMTR Y VDD VNW VPW VSS A0 A1N B0 B1
MXN7 net051 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 ny B0 net051 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 ny A0 net35 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net35 a1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP19 net41 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP20 net41 B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP21 ny A0 net41 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 ny a1 net41 VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI211X1MTR Y VDD VNW VPW VSS A0 A1 B0 C0
MXN5 Y A0 net17 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 net17 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN4 Y C0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNC0 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP6 p1 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXPA1 p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 net045 C0 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 Y B0 net045 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI211X2MTR Y VDD VNW VPW VSS A0 A1 B0 C0
MXN8 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y C0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNC0 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP9 p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA1 p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net045 C0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 Y B0 net045 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI211X4MTR Y VDD VNW VPW VSS A0 A1 B0 C0
MXN12_2 net17__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y A0 net17__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 Y C0 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN13 Y B0 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN13_2 Y B0 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN10_2 Y C0 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXPA1 p1 A1 VDD VNW p12 l=1.3e-07 w=8e-07
MXP12 p1 A0 VDD VNW p12 l=1.3e-07 w=8e-07
MXP12_2 p1 A0 VDD VNW p12 l=1.3e-07 w=8e-07
MXPA1_2 p1 A1 VDD VNW p12 l=1.3e-07 w=8e-07
MXP13_2 net045__2 C0 p1 VNW p12 l=1.3e-07 w=8e-07
MXP14_2 Y B0 net045__2 VNW p12 l=1.3e-07 w=8e-07
MXP14 Y B0 net045 VNW p12 l=1.3e-07 w=8e-07
MXP13 net045 C0 p1 VNW p12 l=1.3e-07 w=8e-07
.ends


.SUBCKT AOI211XLMTR Y VDD VNW VPW VSS A0 A1 B0 C0
MXN8 Y A0 net17 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net17 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 Y C0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNC0 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP9 p1 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXPA1 p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP10 net045 C0 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP11 Y B0 net045 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI21BX1MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=3e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI21BX2MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21BX4MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=3.4e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI2_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21BX8MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI1_MXNA2_2 XI1_n1__2 B0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 ny a0a1 XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1_2 ny a0a1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2_2 ny B0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI2_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI2_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI2_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21BXLMTR Y VDD VNW VPW VSS A0 A1 B0N
mXI0_MXNA2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI0_MXNA1 a0a1 A1 XI0_n1 VPW n12 l=1.3e-07 w=2.1e-07
mXI1_MXNA1 ny a0a1 XI1_n1 VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 XI1_n1 B0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI2_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 a0a1 A0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 a0a1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 ny a0a1 VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA2 ny B0N VDD VNW p12 l=1.3e-07 w=3e-07
mXI2_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI21X1MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI21X2MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21X3MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB1_2 Y A0 XI0_n1__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT AOI21X4MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 Y A0 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21X6MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB1_2 Y A0 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_3 XI0_n1__3 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 Y A0 XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_3 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_3 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21X8MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2_2 XI0_n1__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 Y A0 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 Y A0 XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_3 XI0_n1__3 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_4 XI0_n1__4 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_4 Y A0 XI0_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_3 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_3 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_4 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_4 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI21XLMTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 Y A0 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI221X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN7 Y B0 net26 VPW n12 l=1.3e-07 w=3.6e-07
MXN10 net26 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN9 net17 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN8 Y A0 net17 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y C0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP5 p1 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP6 p1 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 p2 A1 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP9 p2 A0 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 Y C0 p2 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI221X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN14 net26 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B0 net26 VPW n12 l=1.3e-07 w=7.1e-07
MXN12 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXN13 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP10 p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5 p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12 p2 A0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 p2 A1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 Y C0 p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI221X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN18_2 net26__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 Y B0 net26__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN15 Y B0 net26 VPW n12 l=1.3e-07 w=7.1e-07
MXN18 net26 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN17_2 net17__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN16_2 Y A0 net17__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN16 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXN17 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y C0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP14 p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5 p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP14_2 p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 p2 A1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP16 p2 A0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 p2 A0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP15_2 p2 A1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP17 Y C0 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 Y C0 p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI221XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN12 Y B0 net26 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net26 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net17 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 Y A0 net17 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 Y C0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP10 p1 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP11 p1 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP12 p2 A1 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP13 p2 A0 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP14 Y C0 p2 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI222X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN6 Y C0 net29 VPW n12 l=1.3e-07 w=3.6e-07
MXN4 net29 C1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net26 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y B0 net26 VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y A0 net17 VPW n12 l=1.3e-07 w=3.6e-07
MXN2 net17 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP5 p1 C0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP6 p1 C1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP7 p2 B1 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 p2 B0 p1 VNW p12 l=1.3e-07 w=6.2e-07
MXP9 Y A0 p2 VNW p12 l=1.3e-07 w=6.2e-07
MXP10 Y A1 p2 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI222X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN10 net29 C1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 Y C0 net29 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y B0 net26 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net26 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXP11 p1 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12 p1 C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP13 p2 B0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 p2 B1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP15 Y A1 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP16 Y A0 p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI222X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN11_2 Y C0 net29__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN16_2 net29__2 C1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN16 net29 C1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y C0 net29 VPW n12 l=1.3e-07 w=7.1e-07
MXN12_2 Y B0 net26__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 net26__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15 net26 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 Y B0 net26 VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 Y A0 net17__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 net17__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14 net17 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13 Y A0 net17 VPW n12 l=1.3e-07 w=7.1e-07
MXP5 p1 C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17 p1 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 p1 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 p1 C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP18 p2 B0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP19 p2 B1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_2 p2 B1 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 p2 B0 p1 VNW p12 l=1.3e-07 w=8.7e-07
MXP21 Y A0 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP20 Y A1 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 Y A1 p2 VNW p12 l=1.3e-07 w=8.7e-07
MXP21_2 Y A0 p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI222XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN11 Y C0 net29 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net29 C1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net26 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 Y B0 net26 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 Y A0 net17 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net17 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP12 p1 C0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP11 p1 C1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP14 p2 B1 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP13 p2 B0 p1 VNW p12 l=1.3e-07 w=3.6e-07
MXP16 Y A0 p2 VNW p12 l=1.3e-07 w=3.6e-07
MXP15 Y A1 p2 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI22X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 Y B0 XI0_n1B VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A0 XI0_n1A VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI22X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y B0 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI22X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB1_2 Y B0 XI0_n1B__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1B__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y B0 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A0 XI0_n1A__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1A__2 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI22XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1
mXI0_MXNB2 XI0_n1B B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 Y B0 XI0_n1B VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A0 XI0_n1A VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1A A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 XI0_p1 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y A1 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI2B1X1MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN3 net022 a1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=3.6e-07
MXN4 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net36 a1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP5 Y B0 net36 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI2B1X2MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=3e-07
MXN5 net022 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP8 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2B1X4MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN7_2 net022__2 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_2 Y A0 net022__2 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=7.1e-07
MXN7 net022 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP8 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0_2 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
MXP9_2 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2B1X8MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 net022__2 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_2 Y A0 net022__2 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_3 Y A0 net022__3 VPW n12 l=1.3e-07 w=7.1e-07
MXN9_3 net022__3 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_4 net022__4 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_4 Y A0 net022__4 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net022 a1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10_3 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10_4 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0_2 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10_2 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10_3 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0_3 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA0_4 net36 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10_4 net36 a1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP11 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
MXP11_2 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
MXP11_3 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
MXP11_4 Y B0 net36 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2B1XLMTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 a1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN5 net022 a1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNA0 Y A0 net022 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 net36 a1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXPA0 net36 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP7 Y B0 net36 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI2BB1X1MTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI2BB1X2MTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB1X4MTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA2_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2_2 XI24_p1__2 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_2 Y nmin XI24_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB1X8MTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNA1_2 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI23_MXNA2_2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA2_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA2_3 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI24_MXNA2_4 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI23_MXPA2_2 XI23_p1__2 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI23_MXPA1_2 nmin A0N XI23_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2_2 XI24_p1__2 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_2 Y nmin XI24_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_3 Y nmin XI24_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2_3 XI24_p1__3 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2_4 XI24_p1__4 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1_4 Y nmin XI24_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB1XLMTR Y VDD VNW VPW VSS A0N A1N B0
mXI23_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA2 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI24_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI23_MXPA1 nmin A0N XI23_p1 VNW p12 l=1.3e-07 w=3e-07
mXI23_MXPA2 XI23_p1 A1N VDD VNW p12 l=1.3e-07 w=3e-07
mXI24_MXPA2 XI24_p1 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI24_MXPA1 Y nmin XI24_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI2BB2X1MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI2BB2X2MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB2X4MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2_2 XI27_n1__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1_2 Y B0 XI27_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1_2 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1_2 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2_2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB2X8MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI28_MXNA2_2 nmin A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI28_MXNA1_2 nmin A0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2_2 XI27_n1__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1_2 Y B0 XI27_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1_3 Y B0 XI27_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2_3 XI27_n1__3 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2_4 XI27_n1__4 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1_4 Y B0 XI27_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI28_MXPA1_2 nmin A0N XI28_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI28_MXPA2_2 XI28_p1__2 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1_2 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1_3 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPA1_4 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1_2 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2_2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2_3 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1_3 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB1_4 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI27_MXPB2_4 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI2BB2XLMTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI28_MXNA2 nmin A1N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI28_MXNA1 nmin A0N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI27_MXNB2 XI27_n1 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI27_MXNB1 Y B0 XI27_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI27_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI28_MXPA2 XI28_p1 A1N VDD VNW p12 l=1.3e-07 w=3e-07
mXI28_MXPA1 nmin A0N XI28_p1 VNW p12 l=1.3e-07 w=3e-07
mXI27_MXPB2 XI27_p1 B1 VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI27_MXPB1 XI27_p1 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI27_MXPA1 Y nmin XI27_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI31X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0
mXI0_MXNB3 XI0_n1 A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB2 XI0_n2 A1 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 Y A0 XI0_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI31X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0
mXI0_MXNB3 XI0_n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n2 A1 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI31X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0
mXI0_MXNB1_2 Y A0 XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n2__2 A1 XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB3_2 XI0_n1__2 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB3 XI0_n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n2 A1 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB3_2 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI31XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0
mXI0_MXNB3 XI0_n1 A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB2 XI0_n2 A1 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 Y A0 XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI32X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
mXI0_MXNB3 XI0_n1B A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB2 XI0_n2B A1 XI0_n1B VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 Y A0 XI0_n2B VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 XI0_n1A VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 XI0_n1A B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI32X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
mXI0_MXNB3 XI0_n1B A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n2B A1 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n2B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI32X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
mXI0_MXNB1_2 Y A0 XI0_n2B__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n2B__2 A1 XI0_n1B__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB3_2 XI0_n1B__2 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB3 XI0_n1B A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2 XI0_n2B A1 XI0_n1B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 Y A0 XI0_n2B VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n1A__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1A__2 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1A B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1A VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB3_2 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI32XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
mXI0_MXNB3 XI0_n1B A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB2 XI0_n2B A1 XI0_n1B VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 Y A0 XI0_n2B VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 XI0_n1A VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1A B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB3 XI0_p1 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 XI0_p1 A0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y B1 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT AOI33X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN8 net55 B2 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN7 net49 B1 net55 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y B0 net49 VPW n12 l=1.3e-07 w=3.6e-07
MXNA0 Y A0 net43 VPW n12 l=1.3e-07 w=3.6e-07
MXN9 net43 A1 net40 VPW n12 l=1.3e-07 w=3.6e-07
MXN10 net40 A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP12 net057 B2 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP11 net057 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXPB0 net057 B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP15 Y A0 net057 VNW p12 l=1.3e-07 w=6.2e-07
MXP14 Y A1 net057 VNW p12 l=1.3e-07 w=6.2e-07
MXP13 Y A2 net057 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT AOI33X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN13 net55 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net49 B1 net55 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B0 net49 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net43 VPW n12 l=1.3e-07 w=7.1e-07
MXN15 net43 A1 net40 VPW n12 l=1.3e-07 w=7.1e-07
MXN14 net40 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP12 net057 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP11 net057 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPB0 net057 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 Y A0 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 Y A1 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 Y A2 net057 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI33X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN16_2 Y B0 net49__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN17_2 net49__2 B1 net55__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN18_2 net55__2 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN18 net55 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN17 net49 B1 net55 VPW n12 l=1.3e-07 w=7.1e-07
MXN16 Y B0 net49 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0_2 Y A0 net43__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN20_2 net43__2 A1 net40__2 VPW n12 l=1.3e-07 w=7.1e-07
MXN19_2 net40__2 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN19 net40 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN20 net43 A1 net40 VPW n12 l=1.3e-07 w=7.1e-07
MXNA0 Y A0 net43 VPW n12 l=1.3e-07 w=7.1e-07
MXPB0 net057 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16 net057 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17 net057 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net057 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 net057 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPB0_2 net057 B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP20 Y A0 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP19 Y A1 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP18 Y A2 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A2 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_2 Y A1 net057 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 Y A0 net057 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT AOI33XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN13 net55 B2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 net49 B1 net55 VPW n12 l=1.3e-07 w=1.8e-07
MXN11 Y B0 net49 VPW n12 l=1.3e-07 w=1.8e-07
MXNA0 Y A0 net43 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net43 A1 net40 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net40 A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP17 net057 B2 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP16 net057 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXPB0 net057 B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP20 Y A0 net057 VNW p12 l=1.3e-07 w=3.6e-07
MXP19 Y A1 net057 VNW p12 l=1.3e-07 w=3.6e-07
MXP18 Y A2 net057 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT BUFX10MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT BUFX12MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT BUFX14MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT BUFX16MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX18MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT BUFX20MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT BUFX24MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_5 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_11 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_12 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_5 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_11 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_12 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX2MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX32MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_5 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_6 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXNA1_7 ny A VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_11 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_12 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_13 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_14 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_15 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_16 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_5 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_6 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI0_MXPA1_7 ny A VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_11 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_12 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_13 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_14 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_15 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_16 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX3MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=7.2e-07
.ends


.SUBCKT BUFX4MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX5MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3.8e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=4.6e-07
.ends


.SUBCKT BUFX6MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.5e-07
.ends


.SUBCKT BUFX8MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKAND2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1_3 ny A XI0_n1__3 VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=1.05e-06
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=1.05e-06
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=1.05e-06
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=1.05e-06
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X16MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1_3 ny A XI0_n1__3 VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=4.7e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=5.55e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=5.55e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=5.55e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=5.55e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI0_MXPA2_3 ny B VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=9.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.32e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=3.5e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=3.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X3MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKAND2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=4e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=3.05e-07
mXI0_MXNA1_2 ny A XI0_n1__2 VPW n12 l=1.3e-07 w=3.05e-07
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=3.05e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3.05e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=1.04e-06
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=1.04e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKAND2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=5.45e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=5.45e-07
mXI0_MXPA2 ny B VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2_2 ny B VDD VNW p12 l=1.3e-07 w=7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX12MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX16MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=4e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.02e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX1MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=5.1e-07
.ends


.SUBCKT CLKBUFX20MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=1.12e-06
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX24MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=1.03e-06
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=1.03e-06
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKBUFX2MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX32MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_11 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_11 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_12 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX3MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT CLKBUFX40MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1_4 ny A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_8 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_9 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_10 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_11 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_12 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_13 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI1_MXNA1_14 Y ny VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI0_MXPA1_3 ny A VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI0_MXPA1_4 ny A VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI0_MXPA1_5 ny A VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_8 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_9 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_10 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_11 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_12 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_13 Y ny VDD VNW p12 l=1.3e-07 w=1.14e-06
mXI1_MXPA1_14 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX4MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKBUFX6MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=2.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=8.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKBUFX8MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI0_MXPA1_2 ny A VDD VNW p12 l=1.3e-07 w=5.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT CLKINVX12MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.9e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX16MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX1MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=2.55e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=5e-07
.ends


.SUBCKT CLKINVX20MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=1.01e-06
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX24MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=5.6e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=5.6e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=9.2e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=9.2e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=9.2e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=9.2e-07
.ends


.SUBCKT CLKINVX2MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX32MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=1.005e-06
mXI0_MXPA1_11 Y A VDD VNW p12 l=1.3e-07 w=1.005e-06
mXI0_MXPA1_12 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX3MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.4e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT CLKINVX40MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_10 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_11 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_12 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_13 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_14 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_15 Y A VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA1_16 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_17 Y A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_11 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_12 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_13 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_14 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_15 Y A VDD VNW p12 l=1.3e-07 w=1.06e-06
mXI0_MXPA1_16 Y A VDD VNW p12 l=1.3e-07 w=8.65e-07
mXI0_MXPA1_17 Y A VDD VNW p12 l=1.3e-07 w=8.65e-07
.ends


.SUBCKT CLKINVX4MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.85e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.85e-07
.ends


.SUBCKT CLKINVX6MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKINVX8MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7.25e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.25e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7.25e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=7.25e-07
.ends


.SUBCKT CLKMX2X12MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g0_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g0_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g0_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X16MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1_7 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=6.8e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=1.22e-06
mX_g0_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X2MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=2.5e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=7e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X3MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=4.5e-07
.ends


.SUBCKT CLKMX2X4MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X6MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.8e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKMX2X8MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 ns0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI7_MXNOE ny S0 nb VPW n12 l=1.3e-07 w=3.1e-07
mXI6_MXNOE ny ns0 na VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 ns0 S0 VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI7_MXPOEN ny ns0 nb VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN ny S0 na VNW p12 l=1.3e-07 w=7.6e-07
mX_g2_MXPA1 na A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT CLKNAND2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=6.5e-07
.ends


.SUBCKT CLKNAND2X16MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA2_4 XI0_n1__4 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_4 Y A XI0_n1__4 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_5 Y A XI0_n1__5 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_5 XI0_n1__5 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_6 XI0_n1__6 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_6 Y A XI0_n1__6 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_7 Y A XI0_n1__7 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_7 XI0_n1__7 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_8 XI0_n1__8 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_8 Y A XI0_n1__8 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_7 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=7.15e-07
mXI0_MXPA2_8 Y B VDD VNW p12 l=1.3e-07 w=7.15e-07
.ends


.SUBCKT CLKNAND2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8e-07
.ends


.SUBCKT CLKNAND2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.2e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.2e-07
.ends


.SUBCKT CLKNAND2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=7e-07
.ends


.SUBCKT CLKXOR2X12MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g3_MXNA1_2 nB B VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g3_MXNA1_3 nB B VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g2_MXNA1_2 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g2_MXNA1_3 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=3.8e-07
mXI6_MXNOE_2 ny A bB VPW n12 l=1.3e-07 w=3.8e-07
mXI6_MXNOE_3 ny A bB VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=3.8e-07
mXI5_MXNOE_2 ny nA nB VPW n12 l=1.3e-07 w=3.8e-07
mXI5_MXNOE_3 ny nA nB VPW n12 l=1.3e-07 w=4e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.65e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=3e-07
mX_g0_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g3_MXPA1_2 nB B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_3 nB B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_4 nB B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g3_MXPA1_5 nB B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=1.09e-06
mX_g2_MXPA1_2 bB nB VDD VNW p12 l=1.3e-07 w=1.09e-06
mX_g2_MXPA1_3 bB nB VDD VNW p12 l=1.3e-07 w=1.09e-06
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=8.1e-07
mXI6_MXPOEN_2 ny nA bB VNW p12 l=1.3e-07 w=8.3e-07
mXI6_MXPOEN_3 ny nA bB VNW p12 l=1.3e-07 w=8.3e-07
mXI6_MXPOEN_4 ny nA bB VNW p12 l=1.3e-07 w=8.3e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=8.3e-07
mXI5_MXPOEN_2 ny A nB VNW p12 l=1.3e-07 w=8.3e-07
mXI5_MXPOEN_3 ny A nB VNW p12 l=1.3e-07 w=8.3e-07
mXI5_MXPOEN_4 ny A nB VNW p12 l=1.3e-07 w=8.1e-07
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=1.04e-06
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=1.05e-06
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=1.05e-06
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=1.05e-06
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=3.4e-07
.ends


.SUBCKT CLKXOR2X16MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g3_MXNA1_2 nB B VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g3_MXNA1_3 nB B VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g3_MXNA1_4 nB B VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=5e-07
mX_g2_MXNA1_2 bB nB VSS VPW n12 l=1.3e-07 w=5e-07
mX_g2_MXNA1_3 bB nB VSS VPW n12 l=1.3e-07 w=5e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=5.2e-07
mXI6_MXNOE_2 ny A bB VPW n12 l=1.3e-07 w=5.2e-07
mXI6_MXNOE_3 ny A bB VPW n12 l=1.3e-07 w=5.2e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE_2 ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE_3 ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE_4 ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=1.6e-07
mX_g1_MXNA1_2 nA A VSS VPW n12 l=1.3e-07 w=1.6e-07
mX_g1_MXNA1_3 nA A VSS VPW n12 l=1.3e-07 w=1.6e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=5.45e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=5.45e-07
mX_g0_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g0_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g0_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g3_MXPA1_2 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_3 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_4 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_5 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_6 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g3_MXPA1_7 nB B VDD VNW p12 l=1.3e-07 w=8.3e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=1.08e-06
mX_g2_MXPA1_2 bB nB VDD VNW p12 l=1.3e-07 w=1.08e-06
mX_g2_MXPA1_3 bB nB VDD VNW p12 l=1.3e-07 w=1.08e-06
mX_g2_MXPA1_4 bB nB VDD VNW p12 l=1.3e-07 w=1.08e-06
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=8.9e-07
mXI6_MXPOEN_2 ny nA bB VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN_3 ny nA bB VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN_4 ny nA bB VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN_5 ny nA bB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN_2 ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN_3 ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN_4 ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mXI5_MXPOEN_5 ny A nB VNW p12 l=1.3e-07 w=8.8e-07
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=1.33e-06
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=9.55e-07
mX_g0_MXPA1_7 Y ny VDD VNW p12 l=1.3e-07 w=8.55e-07
.ends


.SUBCKT CLKXOR2X2MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=1.9e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.55e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=5.5e-07
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=4.5e-07
.ends


.SUBCKT CLKXOR2X4MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=5.9e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g3_MXPA1_2 nB B VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g2_MXPA1_2 bB nB VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=5.5e-07
mXI6_MXPOEN_2 ny nA bB VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=5.5e-07
mXI5_MXPOEN_2 ny A nB VNW p12 l=1.3e-07 w=5.5e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=4.5e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=4.5e-07
.ends


.SUBCKT CLKXOR2X8MTR Y VDD VNW VPW VSS A B
mX_g3_MXNA1 nB B VSS VPW n12 l=1.3e-07 w=7e-07
mX_g3_MXNA1_2 nB B VSS VPW n12 l=1.3e-07 w=7e-07
mX_g2_MXNA1 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g2_MXNA1_2 bB nB VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g1_MXNA1 nA A VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI6_MXNOE ny A bB VPW n12 l=1.3e-07 w=3.9e-07
mXI6_MXNOE_2 ny A bB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE_2 ny nA nB VPW n12 l=1.3e-07 w=3.9e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=4e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=4e-07
mX_g3_MXPA1 nB B VDD VNW p12 l=1.3e-07 w=6.85e-07
mX_g3_MXPA1_2 nB B VDD VNW p12 l=1.3e-07 w=6.85e-07
mX_g3_MXPA1_3 nB B VDD VNW p12 l=1.3e-07 w=6.85e-07
mX_g3_MXPA1_4 nB B VDD VNW p12 l=1.3e-07 w=6.85e-07
mX_g2_MXPA1 bB nB VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g2_MXPA1_2 bB nB VDD VNW p12 l=1.3e-07 w=1.1e-06
mX_g1_MXPA1 nA A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI6_MXPOEN ny nA bB VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN_2 ny nA bB VNW p12 l=1.3e-07 w=7.3e-07
mXI6_MXPOEN_3 ny nA bB VNW p12 l=1.3e-07 w=7.3e-07
mXI5_MXPOEN ny A nB VNW p12 l=1.3e-07 w=7.3e-07
mXI5_MXPOEN_2 ny A nB VNW p12 l=1.3e-07 w=7.3e-07
mXI5_MXPOEN_3 ny A nB VNW p12 l=1.3e-07 w=7.3e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=9.2e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.8e-07
.ends



.SUBCKT DLY1X1MTR Y VDD VNW VPW VSS A
mX_g1_MXNA1 nmin A VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 nmin1 nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 ny nmin1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 nmin A VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 nmin1 nmin VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 ny nmin1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=5.1e-07
.ends


.SUBCKT DLY1X4MTR Y VDD VNW VPW VSS A
mX_g1_MXNA1 nmin A VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN1 nmin1 nmin VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN3 ny nmin1 VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 nmin A VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP2 nmin1 nmin VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP3 ny nmin1 VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DLY2X1MTR Y VDD VNW VPW VSS A
mXI0_MXNOE ny A XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 A VSS VPW n12 l=1.3e-07 w=1.5e-07
MXN0 VSS ny VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN ny A XI0_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI0_MXPA1 XI0_p1 A VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP0 VDD ny VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DLY2X4MTR Y VDD VNW VPW VSS A
mXI0_MXNOE ny A XI0_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI0_MXNA1 XI0_n1 A VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN0 VSS ny VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPOEN ny A XI0_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI0_MXPA1 XI0_p1 A VDD VNW p12 l=1.3e-07 w=6.5e-07
MXP0 VDD ny VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DLY3X1MTR Y VDD VNW VPW VSS A
mX_g1_MXNA1 nmin A VSS VPW n12 l=1.3e-07 w=1.5e-07
MXN6 net64 nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net70 nmin net64 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 nmin1 nmin net70 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 ny nmin1 net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net67 nmin1 net61 VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net61 nmin1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXPA1 nmin A VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP2 net51 nmin VDD VNW p12 l=1.3e-07 w=3.15e-07
MXP0 net36 nmin net51 VNW p12 l=1.3e-07 w=3.15e-07
MXP1 nmin1 nmin net36 VNW p12 l=1.3e-07 w=3.15e-07
MXP5 ny nmin1 net39 VNW p12 l=1.3e-07 w=3.15e-07
MXP4 net39 nmin1 net48 VNW p12 l=1.3e-07 w=3.15e-07
MXP3 net48 nmin1 VDD VNW p12 l=1.3e-07 w=3.15e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DLY3X4MTR Y VDD VNW VPW VSS A
mX_g1_MXNA1 nmin A VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN6 net64 nmin VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN0 net70 nmin net64 VPW n12 l=1.3e-07 w=4.2e-07
MXN1 nmin1 nmin net70 VPW n12 l=1.3e-07 w=4.2e-07
MXN3 ny nmin1 net67 VPW n12 l=1.3e-07 w=4.2e-07
MXN4 net67 nmin1 net61 VPW n12 l=1.3e-07 w=4.2e-07
MXN5 net61 nmin1 VSS VPW n12 l=1.3e-07 w=4.2e-07
mX_g0_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmin A VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP2 net51 nmin VDD VNW p12 l=1.3e-07 w=7.2e-07
MXP0 net36 nmin net51 VNW p12 l=1.3e-07 w=7.2e-07
MXP1 nmin1 nmin net36 VNW p12 l=1.3e-07 w=7.2e-07
MXP5 ny nmin1 net39 VNW p12 l=1.3e-07 w=7.2e-07
MXP4 net39 nmin1 net48 VNW p12 l=1.3e-07 w=7.2e-07
MXP3 net48 nmin1 VDD VNW p12 l=1.3e-07 w=7.2e-07
mX_g0_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DLY4X1MTR Y VDD VNW VPW VSS A
mXI0_MXNOE na A XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 A VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 na VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNOE ba na XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNOE nba ba XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 ba VSS VPW n12 l=1.3e-07 w=1.5e-07
MXN0 VSS nba VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI3_MXNA1 Y nba VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPOEN na A XI0_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI0_MXPA1 XI0_p1 A VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 na VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPOEN ba na XI1_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI2_MXPOEN nba ba XI2_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI2_MXPA1 XI2_p1 ba VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP0 VDD nba VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI3_MXPA1 Y nba VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DLY4X4MTR Y VDD VNW VPW VSS A
mXI0_MXNOE na A XI0_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 XI0_n1 A VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 na VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI1_MXNOE ba na XI1_n1 VPW n12 l=1.3e-07 w=2.2e-07
mXI2_MXNOE nba ba XI2_n1 VPW n12 l=1.3e-07 w=5.3e-07
mXI2_MXNA1 XI2_n1 ba VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN0 VSS nba VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI3_MXNA1 Y nba VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 Y nba VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPOEN na A XI0_p1 VNW p12 l=1.3e-07 w=2.6e-07
mXI0_MXPA1 XI0_p1 A VDD VNW p12 l=1.3e-07 w=2.6e-07
mXI1_MXPA1 XI1_p1 na VDD VNW p12 l=1.3e-07 w=3.75e-07
mXI1_MXPOEN ba na XI1_p1 VNW p12 l=1.3e-07 w=3.75e-07
mXI2_MXPOEN nba ba XI2_p1 VNW p12 l=1.3e-07 w=6.5e-07
mXI2_MXPA1 XI2_p1 ba VDD VNW p12 l=1.3e-07 w=6.5e-07
MXP0 VDD nba VDD VNW p12 l=1.3e-07 w=6.5e-07
mXI3_MXPA1 Y nba VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 Y nba VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX10MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX12MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX14MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX16MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX18MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX1MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT INVX20MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_10 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX24MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_10 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_11 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_12 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_11 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_12 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX2MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX32MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_8 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_9 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_10 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_11 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_12 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_13 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_14 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_15 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_16 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_7 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_8 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_9 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_10 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_11 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_12 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_13 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_14 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_15 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_16 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX3MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT INVX4MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX5MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT INVX6MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVX8MTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT INVXLMTR Y VDD VNW VPW VSS A
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends



.SUBCKT MX2X12MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=7.1e-07
MXN3 nmin nmsel net42 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_5 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_6 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=8.7e-07
MXP1 net42 S0 nmin VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_5 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2X1MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=3.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=3.7e-07
MXN0 nmin nmsel net38 VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 net38 A VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=4.6e-07
MXP0 net38 S0 nmin VNW p12 l=1.3e-07 w=4.6e-07
mX_g2_MXPA1 net38 A VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT MX2X2MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=4.1e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=5.9e-07
MXN0 nmin nmsel net38 VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1 net38 A VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=5.7e-07
MXP0 net38 S0 nmin VNW p12 l=1.3e-07 w=7.4e-07
mX_g2_MXPA1 net38 A VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2X3MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=6.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=6.7e-07
MXN1 nmin nmsel net42 VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net42 S0 nmin VNW p12 l=1.3e-07 w=8.6e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=6.3e-07
.ends


.SUBCKT MX2X4MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=6.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=6.7e-07
MXN1 nmin nmsel net42 VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net42 S0 nmin VNW p12 l=1.3e-07 w=8.6e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2X6MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=6.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=6.7e-07
MXN1 nmin nmsel net42 VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net42 S0 nmin VNW p12 l=1.3e-07 w=8.6e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2X8MTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=6.7e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=6.7e-07
MXN1 nmin nmsel net42 VPW n12 l=1.3e-07 w=6.7e-07
mX_g2_MXNA1 net42 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net42 S0 nmin VNW p12 l=1.3e-07 w=8.6e-07
mX_g2_MXPA1 net42 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX2XLMTR Y VDD VNW VPW VSS A B S0
mX_g1_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net36 B VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t2 nmin S0 net36 VPW n12 l=1.3e-07 w=2.1e-07
MXN1 nmin nmsel net38 VPW n12 l=1.3e-07 w=2.1e-07
mX_g2_MXNA1 net38 A VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g0_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 net36 B VDD VNW p12 l=1.3e-07 w=2.5e-07
MX_t3 net36 nmsel nmin VNW p12 l=1.3e-07 w=2.5e-07
MXP1 net38 S0 nmin VNW p12 l=1.3e-07 w=2.5e-07
mX_g2_MXPA1 net38 A VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g0_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MX3X1MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=4.1e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=4.7e-07
MX_t4 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=5.6e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=1.9e-07
MX_t0 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=4.5e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=3.7e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
MX_t5 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=6.8e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=2.4e-07
MX_t1 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=6.7e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=4.6e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MX3X2MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=5.8e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=6.4e-07
MX_t4 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=6.6e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t0 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=6.5e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=5.9e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=8.7e-07
MX_t5 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=8.8e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=3.4e-07
MX_t1 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=8.8e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=6.9e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX3X4MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=5.8e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=6.4e-07
MX_t4 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=6.6e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t0 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=6.6e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=6.6e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=8.7e-07
MX_t5 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=8.8e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MX_t1 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=8.8e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=7e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=7.6e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX3X8MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=5e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=6.4e-07
MX_t4 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=6.4e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=6.8e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t0 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=6.6e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=5.3e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y net66 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=7.8e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=7.8e-07
MX_t5 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.6e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=8.6e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP0 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=8.6e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=8.6e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y net66 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX3XLMTR Y VDD VNW VPW VSS A B C S0 S1
mX_g2_MXNA1 net73 S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g4_MXNA1 net69 B VSS VPW n12 l=1.3e-07 w=3.1e-07
MX_t6 nmin0in1 S0 net69 VPW n12 l=1.3e-07 w=3.1e-07
MXN0 nmin0in1 net73 net71 VPW n12 l=1.3e-07 w=3.1e-07
mX_g3_MXNA1 net71 A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g1_MXNA1 net75 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net66 net75 nmin0in1 VPW n12 l=1.3e-07 w=3.1e-07
MX_t2 net66 S1 nmin2 VPW n12 l=1.3e-07 w=3e-07
mX_g5_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=3e-07
mX_g0_MXNA1 Y net66 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXPA1 net73 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 net69 B VDD VNW p12 l=1.3e-07 w=3.8e-07
MX_t7 net69 net73 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 net71 S0 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
mX_g3_MXPA1 net71 A VDD VNW p12 l=1.3e-07 w=3.8e-07
mX_g1_MXPA1 net75 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 nmin0in1 S1 net66 VNW p12 l=1.3e-07 w=3.8e-07
MX_t3 nmin2 net75 net66 VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=3e-07
mX_g0_MXPA1 Y net66 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MX4X1MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI17_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=5.6e-07
MXN0 nmin2in3 nmsel0 net100 VPW n12 l=1.3e-07 w=5.6e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=5.6e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g2_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI18_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=5.6e-07
MXN1 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=5.6e-07
MXN2 nmin0in1 nmsel0 net104 VPW n12 l=1.3e-07 w=5.6e-07
mXI19_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=5.6e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN4 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=5.6e-07
MXN3 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=5.6e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI17_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t9 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=5.9e-07
MX_t11 net98 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=6.8e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g2_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=5.8e-07
mXI18_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=6.8e-07
MX_t7 net102 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=6.1e-07
MXP0 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=6.8e-07
mXI19_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=2.9e-07
MXP2 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=6.8e-07
MXP1 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=6.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MX4X2MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI17_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0 nmin2in3 nmsel0 net100 VPW n12 l=1.3e-07 w=7.1e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=6.8e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN1 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=6.8e-07
MXN2 nmin0in1 nmsel0 net104 VPW n12 l=1.3e-07 w=6.9e-07
mXI19_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MXN6 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=6.9e-07
MXN7 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI17_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t9 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=8.6e-07
MX_t11 net98 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI18_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t7 net102 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
MXP3 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.6e-07
mXI19_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP4 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=8.6e-07
MXP1 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=8.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX4X4MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI17_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0 nmin2in3 nmsel0 net100 VPW n12 l=1.3e-07 w=7.1e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=6.8e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN1 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=6.8e-07
MXN2 nmin0in1 nmsel0 net104 VPW n12 l=1.3e-07 w=6.9e-07
mXI19_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MXN7 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI17_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t9 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=8.6e-07
MX_t11 net98 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI18_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t7 net102 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
MXP3 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.6e-07
mXI19_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP4 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=8.6e-07
MXP1 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=8.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX4X8MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI17_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0 nmin2in3 nmsel0 net100 VPW n12 l=1.3e-07 w=7.1e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=6.8e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN1 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=6.8e-07
MXN2 nmin0in1 nmsel0 net104 VPW n12 l=1.3e-07 w=6.9e-07
mXI19_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
MXN7 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y net97 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI17_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t9 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=8.6e-07
MX_t11 net98 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=8.7e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI18_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t7 net102 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=8.8e-07
MXP3 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=8.6e-07
mXI19_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP4 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=8.6e-07
MXP1 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=8.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y net97 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MX4XLMTR Y VDD VNW VPW VSS A B C D S0 S1
mXI20_MXNA1 net100 C VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN5 nmin2in3 net0110 net100 VPW n12 l=1.3e-07 w=3.1e-07
MX_t10 nmin2in3 S0 net98 VPW n12 l=1.3e-07 w=3.1e-07
mX_g6_MXNA1 net98 D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g2_MXNA1 net0110 S0 VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI21_MXNA1 net102 B VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN6 nmin0in1 S0 net102 VPW n12 l=1.3e-07 w=3.1e-07
MXN7 nmin0in1 net0110 net104 VPW n12 l=1.3e-07 w=3.1e-07
mXI22_MXNA1 net104 A VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net97 nmsel1 nmin0in1 VPW n12 l=1.3e-07 w=3.1e-07
MXN8 net97 S1 nmin2in3 VPW n12 l=1.3e-07 w=3.1e-07
mX_g0_MXNA1 Y net97 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI20_MXPA1 net100 C VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net100 S0 nmin2in3 VNW p12 l=1.3e-07 w=3.8e-07
MX_t11 net98 net0110 nmin2in3 VNW p12 l=1.3e-07 w=3.8e-07
mX_g6_MXPA1 net98 D VDD VNW p12 l=1.3e-07 w=3.8e-07
mX_g2_MXPA1 net0110 S0 VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI21_MXPA1 net102 B VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP4 net102 net0110 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
MXP5 net104 S0 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
mXI22_MXPA1 net104 A VDD VNW p12 l=1.3e-07 w=3.8e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 nmin0in1 S1 net97 VNW p12 l=1.3e-07 w=3.8e-07
MXP6 nmin2in3 nmsel1 net97 VNW p12 l=1.3e-07 w=3.8e-07
mX_g0_MXPA1 Y net97 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MXI2DX1MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=1.9e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=3.7e-07
MXN0 nmin nmsel A VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=4.6e-07
MXP0 A net31 nmin VNW p12 l=1.3e-07 w=4.6e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MXI2DX2MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=2.6e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MXN1 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=4.5e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=3.1e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MXP0 A net31 nmin VNW p12 l=1.3e-07 w=7.4e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2DX4MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=5.2e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MX_t2_2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MXN2 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
MXN2_2 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MX_t3_2 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MXP0 A net31 nmin VNW p12 l=1.3e-07 w=7.1e-07
MXP0_2 A net31 nmin VNW p12 l=1.3e-07 w=7.8e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2DX8MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 nmsel S0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g1_MXNA1_2 net31 nmsel VSS VPW n12 l=1.3e-07 w=5.7e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MX_t2_2 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MX_t2_3 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MX_t2_4 nmin net31 B VPW n12 l=1.3e-07 w=6.1e-07
MXN3 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
MXN3_2 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
MXN3_3 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
MXN3_4 nmin nmsel A VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_3 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_4 Y nmin VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 nmsel S0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g1_MXPA1_2 net31 nmsel VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MX_t3_2 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MX_t3_3 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MX_t3_4 B nmsel nmin VNW p12 l=1.3e-07 w=6.6e-07
MXP0 A net31 nmin VNW p12 l=1.3e-07 w=7.2e-07
MXP0_2 A net31 nmin VNW p12 l=1.3e-07 w=7.7e-07
MXP0_3 A net31 nmin VNW p12 l=1.3e-07 w=7.7e-07
MXP0_4 A net31 nmin VNW p12 l=1.3e-07 w=7.3e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_3 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2DXLMTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 net31 nmsel VSS VPW n12 l=1.3e-07 w=1.9e-07
MX_t2 nmin net31 B VPW n12 l=1.3e-07 w=3e-07
MXN1 nmin nmsel A VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 Y nmin VSS VPW n12 l=1.3e-07 w=3e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 net31 nmsel VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t3 B nmsel nmin VNW p12 l=1.3e-07 w=3e-07
MXP1 A net31 nmin VNW p12 l=1.3e-07 w=3e-07
mX_g2_MXPA1 Y nmin VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MXI2X12MTR Y VDD VNW VPW VSS A B S0
mXI16_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_3 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_4 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_5 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXNA1_6 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=6.7e-07
mX_g0_MXNA1_2 nmsel S0 VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g0_MXNA1_3 nmsel S0 VSS VPW n12 l=1.3e-07 w=5.8e-07
MXN5 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_3 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_4 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_5 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN5_6 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_3 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_4 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_5 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_6 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_3 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_4 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_5 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_6 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI16_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_3 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_4 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_5 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI16_MXPA1_6 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g0_MXPA1_2 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g0_MXPA1_3 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.5e-07
MXP4 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_3 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_4 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_5 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4_6 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_4 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_5 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_6 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_3 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_4 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_5 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_6 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2X1MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y nmsel nmin0 VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=5.3e-07
MX_t1 nmin0 S0 Y VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MXI2X2MTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7e-07
MXN0 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
mXI11_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.6e-07
MX_t1 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
mXI11_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2X3MTR Y VDD VNW VPW VSS A B S0
mXI12_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI12_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN1 Y nmsel nmin0 VPW n12 l=1.3e-07 w=5.4e-07
MXN1_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=5.4e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=5.4e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=5.4e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=4.7e-07
mXI12_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI12_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=5.6e-07
MXP0 nmin0 S0 Y VNW p12 l=1.3e-07 w=6.6e-07
MXP0_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=6.6e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=5.3e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=7.9e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=6.9e-07
.ends


.SUBCKT MXI2X4MTR Y VDD VNW VPW VSS A B S0
mXI13_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI13_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=6e-07
MXN2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN2_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI13_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI13_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP1 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP1_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2X6MTR Y VDD VNW VPW VSS A B S0
mXI14_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXNA1_3 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g0_MXNA1_2 nmsel S0 VSS VPW n12 l=1.3e-07 w=4.4e-07
MXN3 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN3_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN3_3 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_3 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_3 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI14_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI14_MXPA1_3 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g0_MXPA1_2 nmsel S0 VDD VNW p12 l=1.3e-07 w=5.6e-07
MXP2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP2_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP2_3 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_3 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2X8MTR Y VDD VNW VPW VSS A B S0
mXI15_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI15_MXNA1_2 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI15_MXNA1_3 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI15_MXNA1_4 nmin0 A VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=6.4e-07
mX_g0_MXNA1_2 nmsel S0 VSS VPW n12 l=1.3e-07 w=5.8e-07
MXN4 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN4_3 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MXN4_4 Y nmsel nmin0 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_2 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_3 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
MX_t2_4 Y S0 nmin1 VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_2 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_3 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1_4 nmin1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI15_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI15_MXPA1_2 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI15_MXPA1_3 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI15_MXPA1_4 nmin0 A VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.8e-07
mX_g0_MXPA1_2 nmsel S0 VDD VNW p12 l=1.3e-07 w=7.1e-07
MXP3 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP3_3 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP3_4 nmin0 S0 Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_2 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
MX_t3_4 nmin1 nmsel Y VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_2 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_3 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g2_MXPA1_4 nmin1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI2XLMTR Y VDD VNW VPW VSS A B S0
mX_g0_MXNA1 nmsel S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 nmin1 B VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 Y S0 nmin1 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 Y nmsel nmin0 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 nmin0 A VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXPA1 nmsel S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 nmin1 B VDD VNW p12 l=1.3e-07 w=3.6e-07
MX_t3 nmin1 nmsel Y VNW p12 l=1.3e-07 w=3.6e-07
MXP0 nmin0 S0 Y VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPA1 nmin0 A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT MXI3X1MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=2.9e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=3.2e-07
MXN4 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=3.2e-07
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=3.7e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=3.7e-07
MXN5 net115 net104 net98 VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=3.9e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=3.8e-07
MXP1 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=3.9e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=3.9e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=4.6e-07
MXP3 net98 S1 net115 VNW p12 l=1.3e-07 w=4.6e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT MXI3X2MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=4.7e-07
MXN0 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=5.1e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=4.7e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=6.1e-07
MXN1 net115 net104 net98 VPW n12 l=1.3e-07 w=4.1e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t5 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=6.2e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=2.7e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=7.2e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=7.2e-07
MXP0 net98 S1 net115 VNW p12 l=1.3e-07 w=7e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=3.2e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=6e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI3X4MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=4.7e-07
MXN0 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=6.1e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=4.7e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=6.1e-07
MXN1 net115 net104 net98 VPW n12 l=1.3e-07 w=4.1e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=4.7e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t5 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=7.4e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=8.1e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=8.1e-07
MXP0 net98 S1 net115 VNW p12 l=1.3e-07 w=7e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI3X8MTR Y VDD VNW VPW VSS A B C S0 S1
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=4.7e-07
MXN0 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=6.1e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=4.7e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=3e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=6.1e-07
MXN1 net115 net104 net98 VPW n12 l=1.3e-07 w=4.3e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y net115 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t5 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=7.4e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=8.2e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=7.1e-07
MXP0 net98 S1 net115 VNW p12 l=1.3e-07 w=7e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y net115 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI3XLMTR Y VDD VNW VPW VSS A B C S0 S1
mX_g4_MXNA1 net86 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g6_MXNA1 net74 B VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t6 nmin0in1 S0 net74 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 nmin0in1 net86 net80 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 net80 A VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 Y net115 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 nmin2 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net92 nmin2 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t2 net115 S1 net92 VPW n12 l=1.3e-07 w=2.1e-07
MXN3 net115 net104 net98 VPW n12 l=1.3e-07 w=2.1e-07
mX_g2_MXNA1 net98 nmin0in1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g1_MXNA1 net104 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXPA1 net86 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g6_MXPA1 net74 B VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t7 net74 net86 nmin0in1 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net80 S0 nmin0in1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 net80 A VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 Y net115 VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g7_MXPA1 nmin2 C VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPA1 net92 nmin2 VDD VNW p12 l=1.3e-07 w=2.5e-07
MX_t3 net92 net104 net115 VNW p12 l=1.3e-07 w=2.5e-07
MXP2 net98 S1 net115 VNW p12 l=1.3e-07 w=2.5e-07
mX_g2_MXPA1 net98 nmin0in1 VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g1_MXPA1 net104 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT MXI4X1MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=3.2e-07
MXN2 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=3.2e-07
MXN1 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=3.2e-07
mXI18_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g4_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=3.2e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=3.2e-07
MXN0 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=3.2e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=3.7e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=3.7e-07
MXN3 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=3.7e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=3.9e-07
MXP2 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=3.9e-07
MXP1 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=3.9e-07
mXI18_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=3.9e-07
mX_g4_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=3.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=3.9e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=3.9e-07
MXP0 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=3.9e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=3.9e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=4.6e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=4.6e-07
MXP3 net112 S1 net99 VNW p12 l=1.3e-07 w=4.6e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=4.6e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MXI4X2MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=5.1e-07
MXN2 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=5.1e-07
MXN1 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=4.2e-07
mXI18_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=4.4e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=4e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=4.9e-07
MXN0 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=5.2e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=4.8e-07
MXN3 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=4.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP2 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=6.3e-07
MXP4 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mXI18_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g4_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=5.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=5.7e-07
MXP0 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=6.3e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=7.4e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=7.4e-07
MXP5 net112 S1 net99 VNW p12 l=1.3e-07 w=7.4e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI4X4MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN5 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=6.1e-07
MXN4 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=4e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=6.1e-07
MXN0 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=6.1e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=5e-07
MXN3 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=4.4e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP7 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=7.4e-07
MXP6 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mXI18_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=5.7e-07
MXP0 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=7.4e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=8.4e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=8.4e-07
MXP5 net112 S1 net99 VNW p12 l=1.3e-07 w=8.3e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI4X8MTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN5 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=6.1e-07
MXN4 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=6.1e-07
mXI18_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=4e-07
mX_g4_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=5.2e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=4e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=6.1e-07
MXN0 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=6.1e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=6.1e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=5e-07
MXN3 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=4.4e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=3e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_3 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_4 Y net99 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP7 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=7.4e-07
MXP6 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=5.7e-07
mXI18_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g4_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=5.7e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=5.7e-07
MXP0 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=7.4e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=7.4e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=8.4e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=8.4e-07
MXP5 net112 S1 net99 VNW p12 l=1.3e-07 w=8.3e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_3 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_4 Y net99 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MXI4XLMTR Y VDD VNW VPW VSS A B C D S0 S1
mXI19_MXNA1 net106 A VSS VPW n12 l=1.3e-07 w=3e-07
MXN6 nmin0in1 nmsel0 net106 VPW n12 l=1.3e-07 w=3e-07
MXN5 nmin0in1 S0 net104 VPW n12 l=1.3e-07 w=1.8e-07
mXI21_MXNA1 net104 B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI22_MXNA1 nmsel0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 net100 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t10 nmin2in3 S0 net100 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 nmin2in3 nmsel0 net102 VPW n12 l=1.3e-07 w=1.8e-07
mXI17_MXNA1 net102 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNA1 net110 nmin2in3 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t2 net99 S1 net110 VPW n12 l=1.3e-07 w=2.1e-07
MXN7 net99 nmsel1 net112 VPW n12 l=1.3e-07 w=2.1e-07
mX_g1_MXNA1 nmsel1 S1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI20_MXNA1 net112 nmin0in1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g0_MXNA1 Y net99 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXPA1 net106 A VDD VNW p12 l=1.3e-07 w=3e-07
MXP6 net106 S0 nmin0in1 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 net104 nmsel0 nmin0in1 VNW p12 l=1.3e-07 w=2.3e-07
mXI21_MXPA1 net104 B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI22_MXPA1 nmsel0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g8_MXPA1 net100 D VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t11 net100 nmsel0 nmin2in3 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net102 S0 nmin2in3 VNW p12 l=1.3e-07 w=2.3e-07
mXI17_MXPA1 net102 C VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPA1 net110 nmin2in3 VDD VNW p12 l=1.3e-07 w=3e-07
MX_t3 net110 nmsel1 net99 VNW p12 l=1.3e-07 w=2.5e-07
MXP7 net112 S1 net99 VNW p12 l=1.3e-07 w=2.5e-07
mX_g1_MXPA1 nmsel1 S1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI20_MXPA1 net112 nmin0in1 VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g0_MXPA1 Y net99 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND2BX12MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_3 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2_2 XI1_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y a XI1_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 XI1_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 XI1_n1__4 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y a XI1_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y a XI1_n1__5 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_5 XI1_n1__5 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_6 XI1_n1__6 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y a XI1_n1__6 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_2 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_3 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2BX1MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND2BX2MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2BX4MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2_2 XI1_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2BX8MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2_2 XI1_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y a XI1_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 XI1_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 XI1_n1__4 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y a XI1_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_2 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2BXLMTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 XI1_n1 B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y a XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n1__4 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A XI0_n1__5 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 XI0_n1__5 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_6 XI0_n1__6 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A XI0_n1__6 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2X1MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2X3MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=4.4e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT NAND2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2X5MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_3 XI0_n1 B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 Y A XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 Y A XI0_n1 VPW n12 l=1.3e-07 w=6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=7.3e-07
.ends


.SUBCKT NAND2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2_2 XI0_n1__2 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n1__3 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n1__4 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n1__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND2XLMTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 XI0_n1 B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND3BX1MTR Y VDD VNW VPW VSS AN B C
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA3 XI1_n1 C VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA2 XI1_n2 B XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y a XI1_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND3BX2MTR Y VDD VNW VPW VSS AN B C
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA3 XI1_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n2 B XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3BX4MTR Y VDD VNW VPW VSS AN B C
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA3_2 XI1_n1__2 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 XI1_n2__2 B XI1_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n2 B XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA3 XI1_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3BXLMTR Y VDD VNW VPW VSS AN B C
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA3 XI1_n1 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n2 B XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y a XI1_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND3X12MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_5 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_6 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_6 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_4 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_5 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_6 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3X1MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND3X2MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3X3MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y A XI0_n2__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT NAND3X4MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3X6MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n2__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n2__3 B XI0_n1__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n1__3 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND3X8MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3_2 XI0_n1__2 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_2 XI0_n2__2 B XI0_n1__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y A XI0_n2__2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_3 Y A XI0_n2__3 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_3 XI0_n2__3 B XI0_n1__3 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3_3 XI0_n1__3 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3_4 XI0_n1__4 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_4 XI0_n2__4 B XI0_n1__4 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_4 Y A XI0_n2__4 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA3_4 Y C VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT NAND3XLMTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 XI0_n1 C VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n2 B XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND4BBX1MTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net43 D VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net47 C net43 VPW n12 l=1.3e-07 w=3.6e-07
MXN0 net51 B net47 VPW n12 l=1.3e-07 w=3.6e-07
MXNA Y A net51 VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 Y D VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP1 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
MXPA Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT NAND4BBX2MTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=3e-07
MXN7 net43 D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN6 net47 C net43 VPW n12 l=1.3e-07 w=7.1e-07
MXN5 net51 B net47 VPW n12 l=1.3e-07 w=7.1e-07
MXNA Y A net51 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP5 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=3.7e-07
.ends


.SUBCKT NAND4BBX4MTR Y VDD VNW VPW VSS AN BN C D
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN11 net43 D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 net43 D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 net47 C net43 VPW n12 l=1.3e-07 w=7.1e-07
MXN10_2 net47 C net43 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net51 B net47 VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 net51 B net47 VPW n12 l=1.3e-07 w=7.1e-07
MXNA Y A net51 VPW n12 l=1.3e-07 w=7.1e-07
MXNA_2 Y A net51 VPW n12 l=1.3e-07 w=7.2e-07
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP5 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A VDD VNW p12 l=1.3e-07 w=8e-07
MXPA_2 Y A VDD VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT NAND4BBXLMTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN12 net43 D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 net47 C net43 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net51 B net47 VPW n12 l=1.3e-07 w=1.8e-07
MXNA Y A net51 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP10 Y D VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP9 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP8 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
MXPA Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT NAND4BX1MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA4 XI1_n1 D VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA3 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y a XI1_n3 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND4BX2MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA4 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA3 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4BX4MTR Y VDD VNW VPW VSS AN B C D
mXI1_MXNA4 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA4_2 XI1_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA3 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA3_2 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a XI1_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a XI1_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT NAND4BXLMTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA4 XI1_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA3 XI1_n2 C XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n3 B XI1_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y a XI1_n3 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y a VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NAND4X12MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_5 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_6 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_5 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_6 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_6 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_3 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_5 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_6 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_4 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_5 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_6 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_6 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4X1MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NAND4X2MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4X4MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4_2 XI0_n1__2 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2__2 C XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3__2 B XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n3__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4X6MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_3 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4X8MTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_2 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_3 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA4_4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A XI0_n3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_2 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_3 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA4_4 Y D VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_4 Y C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 Y B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NAND4XLMTR Y VDD VNW VPW VSS A B C D
mXI0_MXNA4 XI0_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA3 XI0_n2 C XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n3 B XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A XI0_n3 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA4 Y D VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA3 Y C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 Y B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR2BX12MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_3 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_5 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_6 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_2 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_3 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPA2_2 XI1_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y a XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y a XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y a XI1_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_5 XI1_p1__5 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_6 XI1_p1__6 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y a XI1_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2BX1MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NOR2BX2MTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2BX4MTR Y VDD VNW VPW VSS AN B
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPA2_2 XI1_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT NOR2BX8MTR Y VDD VNW VPW VSS AN B
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y a VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 a AN VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPA2_2 XI1_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y a XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y a XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_3 XI1_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_4 XI1_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y a XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA1_2 a AN VDD VNW p12 l=1.3e-07 w=7.5e-07
.ends


.SUBCKT NOR2BXLMTR Y VDD VNW VPW VSS AN B
mXI0_MXNA1 a AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y a VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 a AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1 B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y a XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_6 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 XI0_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y A XI0_p1__5 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 XI0_p1__5 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_6 XI0_p1__6 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y A XI0_p1__6 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2X1MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NOR2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2X3MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT NOR2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2X5MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=6e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1_3 Y A XI0_p1__3 VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=7.3e-07
.ends


.SUBCKT NOR2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 XI0_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y A XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR2XLMTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR3BX1MTR Y VDD VNW VPW VSS AN B C
mX_g0_MXNA1 net38 AN VSS VPW n12 l=1.3e-07 w=1.9e-07
MX_t5 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y net38 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 net38 AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t0 VDD C net33 VNW p12 l=1.3e-07 w=6.2e-07
MXP0 net33 B net30 VNW p12 l=1.3e-07 w=6.2e-07
MXP1 net30 net38 Y VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NOR3BX2MTR Y VDD VNW VPW VSS AN B C
mX_g0_MXNA1 net38 AN VSS VPW n12 l=1.3e-07 w=3e-07
MX_t5 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN3 Y net38 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 net38 AN VDD VNW p12 l=1.3e-07 w=3.7e-07
MX_t0 VDD C net33 VNW p12 l=1.3e-07 w=8.7e-07
MXP2 net33 B net30 VNW p12 l=1.3e-07 w=8.7e-07
MXP3 net30 net38 Y VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3BX4MTR Y VDD VNW VPW VSS AN B C
mX_g0_MXNA1 net38 AN VSS VPW n12 l=1.3e-07 w=6.1e-07
MX_t5 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 Y net38 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5_2 Y net38 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MX_t5_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 net38 AN VDD VNW p12 l=1.3e-07 w=7.4e-07
MX_t0_2 VDD C net33__2 VNW p12 l=1.3e-07 w=8.1e-07
MXP4_2 net33__2 B net30__2 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_2 net30__2 net38 Y VNW p12 l=1.3e-07 w=8.1e-07
MXP5 net30 net38 Y VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net33 B net30 VNW p12 l=1.3e-07 w=8.7e-07
MX_t0 VDD C net33 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3BXLMTR Y VDD VNW VPW VSS AN B C
mX_g0_MXNA1 net38 AN VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t5 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN6 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 Y net38 VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXPA1 net38 AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t0 VDD C net33 VNW p12 l=1.3e-07 w=3.6e-07
MXP4 net33 B net30 VNW p12 l=1.3e-07 w=3.6e-07
MXP5 net30 net38 Y VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR3X12MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_5 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_5 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y A VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA2_6 Y B VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXNA3_6 Y C VSS VPW n12 l=1.3e-07 w=6.8e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_2 Y A XI0_p2__2 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_3 Y A XI0_p2__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_3 XI0_p2__3 B XI0_p1__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_3 XI0_p1__3 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_4 XI0_p1__4 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_4 XI0_p2__4 B XI0_p1__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_4 Y A XI0_p2__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_5 Y A XI0_p2__5 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2_5 XI0_p2__5 B XI0_p1__5 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3_5 XI0_p1__5 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_6 XI0_p1__6 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_6 XI0_p2__6 B XI0_p1__6 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_6 Y A XI0_p2__6 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3X1MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT NOR3X2MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3X4MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p2__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3X6MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y A XI0_p2__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y A XI0_p2__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_3 XI0_p2__3 B XI0_p1__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_3 XI0_p1__3 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.1e-07
.ends


.SUBCKT NOR3X8MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_4 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3_4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_2 Y A XI0_p2__2 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_3 Y A XI0_p2__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_3 XI0_p2__3 B XI0_p1__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_3 XI0_p1__3 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA3_4 XI0_p1__4 C VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA2_4 XI0_p2__4 B XI0_p1__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_4 Y A XI0_p2__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR3XLMTR Y VDD VNW VPW VSS A B C
mXI0_MXNA3 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y A XI0_p2 VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT NOR4BBX1MTR Y VDD VNW VPW VSS AN BN C D
MXN2 Y D VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=2.5e-07
MXPD net90 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0 net86 C net90 VNW p12 l=1.3e-07 w=8.7e-07
MXP1 net068 B net86 VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y A net068 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=3e-07
.ends


.SUBCKT NOR4BBX2MTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=4.9e-07
MXN5 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=6e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=6e-07
MXP5_2 Y A net068__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_2 net068__2 B net86__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 net86__2 C net90__2 VNW p12 l=1.3e-07 w=8.7e-07
MXPD_2 net90__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXPD net90 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP3 net86 C net90 VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net068 B net86 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y A net068 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BBX4MTR Y VDD VNW VPW VSS AN BN C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_2 A AN VSS VPW n12 l=1.3e-07 w=5e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=5e-07
mXI1_MXNA1_2 B BN VSS VPW n12 l=1.3e-07 w=5e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN9 Y D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN9_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI0_MXPA1_2 A AN VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI1_MXPA1_2 B BN VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP5_2 Y A net068__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_2 net068__2 B net86__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP6_2 net86__2 C net90__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP7_2 net90__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7_3 net90__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6_3 net86__3 C net90__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_3 net068__3 B net86__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_3 Y A net068__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_4 Y A net068__4 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_4 net068__4 B net86__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP6_4 net86__4 C net90__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_4 net90__4 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7 net90 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6 net86 C net90 VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net068 B net86 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y A net068 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BBXLMTR Y VDD VNW VPW VSS AN BN C D
MXN5 Y D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 B BN VSS VPW n12 l=1.3e-07 w=1.9e-07
MXP5 net90 D VDD VNW p12 l=1.3e-07 w=4.7e-07
MXP4 net86 C net90 VNW p12 l=1.3e-07 w=4.7e-07
MXP3 net068 B net86 VNW p12 l=1.3e-07 w=4.7e-07
MXP2 Y A net068 VNW p12 l=1.3e-07 w=4.7e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 B BN VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT NOR4BX1MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=2.5e-07
MXN2 Y D VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=3e-07
MXPD net33 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0 net29 C net33 VNW p12 l=1.3e-07 w=8.7e-07
MXP1 net25 B net29 VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y A net25 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BX2MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=4.9e-07
MXN5 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=6e-07
MXPA_2 Y A net25__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 net25__2 B net29__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP1_2 net29__2 C net33__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP2_2 net33__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 net33 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP1 net29 C net33 VNW p12 l=1.3e-07 w=8.7e-07
MXP0 net25 B net29 VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A net25 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BX4MTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=5e-07
mXI0_MXNA1_2 A AN VSS VPW n12 l=1.3e-07 w=5e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y C VSS VPW n12 l=1.3e-07 w=6e-07
MXN6 Y D VSS VPW n12 l=1.3e-07 w=6e-07
MXN6_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI0_MXPA1_2 A AN VDD VNW p12 l=1.3e-07 w=6.1e-07
MXPA_2 Y A net25__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 net25__2 B net29__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP4_2 net29__2 C net33__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 net33__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5_3 net33__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4_3 net29__3 C net33__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_3 net25__3 B net29__3 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_3 Y A net25__3 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_4 Y A net25__4 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_4 net25__4 B net29__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP4_4 net29__4 C net33__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_4 net33__4 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP5 net33 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net29 C net33 VNW p12 l=1.3e-07 w=8.7e-07
MXP3 net25 B net29 VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A net25 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4BXLMTR Y VDD VNW VPW VSS AN B C D
mXI0_MXNA1 A AN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 Y D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN7 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 A AN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net33 D VDD VNW p12 l=1.3e-07 w=4.7e-07
MXP10 net29 C net33 VNW p12 l=1.3e-07 w=4.7e-07
MXP9 net25 B net29 VNW p12 l=1.3e-07 w=4.7e-07
MXP8 Y A net25 VNW p12 l=1.3e-07 w=4.7e-07
.ends


.SUBCKT NOR4X12MTR Y VDD VNW VPW VSS A B C D
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNC Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNC_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB_2 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_3 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNB_3 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNC_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_3 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_4 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNC_4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB_4 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_4 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_5 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNB_5 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNC_5 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_5 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_6 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNC_6 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB_6 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_6 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_3 Y A net37__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_3 net37__3 B net40__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP7_3 net40__3 C net43__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net43__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net43__4 D VDD VNW p12 l=1.3e-07 w=7.8e-07
MXP7_4 net40__4 C net43__4 VNW p12 l=1.3e-07 w=7.8e-07
MXP5_4 net37__4 B net40__4 VNW p12 l=1.3e-07 w=7.8e-07
MXPA_4 Y A net37__4 VNW p12 l=1.3e-07 w=7.8e-07
MXPA_5 Y A net37__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_5 net37__5 B net40__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_5 net40__5 C net43__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_5 net43__5 D VDD VNW p12 l=1.3e-07 w=7.8e-07
MXP8_6 net43__6 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7_6 net40__6 C net43__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_6 net37__6 B net40__6 VNW p12 l=1.3e-07 w=8.1e-07
MXPA_6 Y A net37__6 VNW p12 l=1.3e-07 w=8.1e-07
MXPA_7 Y A net37__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_7 net37__7 B net40__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_7 net40__7 C net43__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_7 net43__7 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP8_8 net43__8 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7_8 net40__8 C net43__8 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_8 net37__8 B net40__8 VNW p12 l=1.3e-07 w=8.1e-07
MXPA_8 Y A net37__8 VNW p12 l=1.3e-07 w=8.1e-07
MXPA_9 Y A net37__9 VNW p12 l=1.3e-07 w=8.1e-07
MXP5_9 net37__9 B net40__9 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_9 net40__9 C net43__9 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_9 net43__9 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP8_10 net43__10 D VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7_10 net40__10 C net43__10 VNW p12 l=1.3e-07 w=7.8e-07
MXP5_10 net37__10 B net40__10 VNW p12 l=1.3e-07 w=7.8e-07
MXPA_10 Y A net37__10 VNW p12 l=1.3e-07 w=7.8e-07
MXPA_11 Y A net37__11 VNW p12 l=1.3e-07 w=7.8e-07
MXP5_11 net37__11 B net40__11 VNW p12 l=1.3e-07 w=7.8e-07
MXP7_11 net40__11 C net43__11 VNW p12 l=1.3e-07 w=7.8e-07
MXP8_11 net43__11 D VDD VNW p12 l=1.3e-07 w=7.8e-07
MXP8_12 net43__12 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7_12 net40__12 C net43__12 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_12 net37__12 B net40__12 VNW p12 l=1.3e-07 w=8.7e-07
MXPA_12 Y A net37__12 VNW p12 l=1.3e-07 w=8.7e-07
MXPA Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP7 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4X1MTR Y VDD VNW VPW VSS A B C D
MXN7 Y D VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y C VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN5 Y B VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4X2MTR Y VDD VNW VPW VSS A B C D
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP13_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4X4MTR Y VDD VNW VPW VSS A B C D
MXN14 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13 Y B VSS VPW n12 l=1.3e-07 w=6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=6e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_3 Y A net37__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_3 net37__3 B net40__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP12_3 net40__3 C net43__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net43__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net43__4 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_4 net40__4 C net43__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP17_4 net37__4 B net40__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP18_4 Y A net37__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP18 Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
MXP17 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4X6MTR Y VDD VNW VPW VSS A B C D
MXNA Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_3 Y B VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_3 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_3 Y A net37__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_3 net37__3 B net40__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP12_3 net40__3 C net43__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net43__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net43__4 D VDD VNW p12 l=1.3e-07 w=7.8e-07
MXP12_4 net40__4 C net43__4 VNW p12 l=1.3e-07 w=7.8e-07
MXP17_4 net37__4 B net40__4 VNW p12 l=1.3e-07 w=7.8e-07
MXP18_4 Y A net37__4 VNW p12 l=1.3e-07 w=7.8e-07
MXP18_5 Y A net37__5 VNW p12 l=1.3e-07 w=8.2e-07
MXP17_5 net37__5 B net40__5 VNW p12 l=1.3e-07 w=8.2e-07
MXP12_5 net40__5 C net43__5 VNW p12 l=1.3e-07 w=8.2e-07
MXP8_5 net43__5 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_6 net43__6 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_6 net40__6 C net43__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP17_6 net37__6 B net40__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP18_6 Y A net37__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP18 Y A net37 VNW p12 l=1.3e-07 w=8.1e-07
MXP17 net37 B net40 VNW p12 l=1.3e-07 w=8.1e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=8.1e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.1e-07
.ends


.SUBCKT NOR4X8MTR Y VDD VNW VPW VSS A B C D
MXN14 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B VSS VPW n12 l=1.3e-07 w=6e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=6e-07
MXNA_2 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXN9_2 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_3 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_3 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_3 Y B VSS VPW n12 l=1.3e-07 w=6.3e-07
MXNA_3 Y A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNA_4 Y A VSS VPW n12 l=1.3e-07 w=6e-07
MXN11_4 Y B VSS VPW n12 l=1.3e-07 w=6e-07
MXN9_4 Y C VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_4 Y D VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP8_2 net43__2 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 net40__2 C net43__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_2 net37__2 B net40__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 Y A net37__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_3 Y A net37__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_3 net37__3 B net40__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP12_3 net40__3 C net43__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net43__3 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net43__4 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_4 net40__4 C net43__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP19_4 net37__4 B net40__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP20_4 Y A net37__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP20_5 Y A net37__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP19_5 net37__5 B net40__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP12_5 net40__5 C net43__5 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_5 net43__5 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_6 net43__6 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_6 net40__6 C net43__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP19_6 net37__6 B net40__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP20_6 Y A net37__6 VNW p12 l=1.3e-07 w=8.1e-07
MXP20_7 Y A net37__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP19_7 net37__7 B net40__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP12_7 net40__7 C net43__7 VNW p12 l=1.3e-07 w=8.1e-07
MXP8_7 net43__7 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_8 net43__8 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_8 net40__8 C net43__8 VNW p12 l=1.3e-07 w=8.7e-07
MXP19_8 net37__8 B net40__8 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_8 Y A net37__8 VNW p12 l=1.3e-07 w=8.7e-07
MXP20 Y A net37 VNW p12 l=1.3e-07 w=8.7e-07
MXP19 net37 B net40 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT NOR4XLMTR Y VDD VNW VPW VSS A B C D
MXN10 Y D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 Y C VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 Y B VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNA Y A VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP8 net43 D VDD VNW p12 l=1.3e-07 w=4.7e-07
MXP12 net40 C net43 VNW p12 l=1.3e-07 w=4.7e-07
MXP13 net37 B net40 VNW p12 l=1.3e-07 w=4.7e-07
MXP14 Y A net37 VNW p12 l=1.3e-07 w=4.7e-07
.ends


.SUBCKT OA21X1MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OA21X2MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA21X4MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA21X8MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPB2_2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPB1_2 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 ny B0 VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA21XLMTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 ny B0 XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPB1 ny A0 XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 ny B0 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OA22X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 ny A1 net48 VPW n12 l=1.3e-07 w=2.3e-07
MXN3 ny A0 net48 VPW n12 l=1.3e-07 w=2.3e-07
MXN4 net48 B0 VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN5 net48 B1 VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP6 net67 A1 VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP5 ny A0 net67 VNW p12 l=1.3e-07 w=3.1e-07
MXP4 ny B0 net73 VNW p12 l=1.3e-07 w=3.1e-07
MXP8 net73 B1 VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OA22X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 ny A1 net45 VPW n12 l=1.3e-07 w=3.6e-07
MXN7 ny A0 net45 VPW n12 l=1.3e-07 w=3.6e-07
MXN8 net45 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN9 net45 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP7 net60 A1 VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP9 ny A0 net60 VNW p12 l=1.3e-07 w=5.1e-07
MXP10 ny B0 net66 VNW p12 l=1.3e-07 w=5.1e-07
MXP8 net66 B1 VDD VNW p12 l=1.3e-07 w=5.1e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA22X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 ny A1 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN10 ny A0 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 net45 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net45 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP11 net60 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12 ny A0 net60 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 ny B0 net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net66 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA22X8MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN13 ny A0 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 ny A1 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 ny A1 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 ny A0 net45 VPW n12 l=1.3e-07 w=7.1e-07
MXN14 net45 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15 net45 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 net45 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 net45 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP15_2 ny A0 net60__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14_2 net60__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP14 net60 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 ny A0 net60 VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 ny B0 net66__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net66__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net66 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16 ny B0 net66 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OA22XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 ny A1 net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 ny A0 net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net45 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net45 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP7 net60 A1 VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 ny A0 net60 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 ny B0 net66 VNW p12 l=1.3e-07 w=2.3e-07
MXP8 net66 B1 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI211X1MTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI211X2MTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI211X4MTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n2__2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPC1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPB1_2 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI211X8MTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC1_3 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2_3 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC2_4 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNC1_4 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n2__2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 XI0_n2__3 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 XI0_n2__3 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_4 XI0_n2__4 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y B0 XI0_n2__4 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPC1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2_3 XI0_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC1_3 Y A0 XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC1_4 Y A0 XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2_4 XI0_p1__4 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPB1_2 Y C0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPB1_3 Y C0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_3 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPA1_4 Y B0 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI0_MXPB1_4 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI211XLMTR Y VDD VNW VPW VSS A0 A1 B0 C0
mXI0_MXNC1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNC2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 XI0_n2 C0 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 XI0_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPC1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPC2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI21BX1MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT OAI21BX2MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=3.7e-07
.ends


.SUBCKT OAI21BX4MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXPB2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=7.4e-07
.ends


.SUBCKT OAI21BX8MTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_3 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_3 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_4 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_4 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXPB2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_3 Y A0 XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_3 XI1_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_4 XI1_p1__4 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_4 Y A0 XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y b0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21BXLMTR Y VDD VNW VPW VSS A0 A1 B0N
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y b0 XI1_n1 VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA1 b0 B0N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y b0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 b0 B0N VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT OAI21X1MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI21X2MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21X3MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1_2 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXPB2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT OAI21X4MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21X6MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_3 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_3 Y A0 XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_3 XI0_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21X8MTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_2 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_3 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_3 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB1_4 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNB2_4 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPB2_2 XI0_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_2 Y A0 XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_3 Y A0 XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_3 XI0_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2_4 XI0_p1__4 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1_4 Y A0 XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI21XLMTR Y VDD VNW VPW VSS A0 A1 B0
mXI0_MXNB2 XI0_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNB1 XI0_n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 Y B0 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPB2 XI0_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPB1 Y A0 XI0_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI221X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN2 net33 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net33 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 net25 A1 net33 VPW n12 l=1.3e-07 w=3.6e-07
MXN1 net25 A0 net33 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y C0 net25 VPW n12 l=1.3e-07 w=3.6e-07
MXP0 Y B0 net46 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 net46 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP2 net58 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP1 Y A0 net58 VNW p12 l=1.3e-07 w=6.2e-07
MXP3 Y C0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI221X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN7 net33 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 net33 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 net25 A1 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN8 net25 A0 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 net25 VPW n12 l=1.3e-07 w=7.1e-07
MXP5 Y B0 net073 VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net073 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP6 net059 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP7 Y A0 net059 VNW p12 l=1.3e-07 w=8.7e-07
MXP3 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI221X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN11 net33 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 net33 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10_2 net33 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 net33 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net25 A0 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net25 A1 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 net25 A1 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN12_2 net25 A0 net33 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 net25 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y C0 net25 VPW n12 l=1.3e-07 w=7.1e-07
MXP9_2 Y B0 net077__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net077__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net077 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y B0 net077 VNW p12 l=1.3e-07 w=8.7e-07
MXP11_2 Y A0 net069__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP10_2 net069__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net069 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP11 Y A0 net069 VNW p12 l=1.3e-07 w=8.7e-07
MXP3 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI221XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0
MXN10 net33 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net33 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net25 A1 net33 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net25 A0 net33 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 Y C0 net25 VPW n12 l=1.3e-07 w=1.8e-07
MXP5 Y B0 net069 VNW p12 l=1.3e-07 w=3.6e-07
MXP4 net069 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP7 net077 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP6 Y A0 net077 VNW p12 l=1.3e-07 w=3.6e-07
MXP3 Y C0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI222X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN2 net28 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 net28 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN0 net24 A1 net28 VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net24 A0 net28 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 Y C0 net24 VPW n12 l=1.3e-07 w=3.6e-07
MXN4 Y C1 net24 VPW n12 l=1.3e-07 w=3.6e-07
MXP6 Y B0 net089 VNW p12 l=1.3e-07 w=6.2e-07
MXP5 net089 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP9 net083 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP10 Y A0 net083 VNW p12 l=1.3e-07 w=6.2e-07
MXP7 Y C0 net59 VNW p12 l=1.3e-07 w=6.2e-07
MXP8 net59 C1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI222X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN8 net28 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN10 net28 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net24 A1 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN7 net24 A0 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXN5 Y C1 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXP12 Y B0 net094 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 net094 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP14 net088 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15 Y A0 net088 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 Y C0 net59 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net59 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI222X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN13 net28 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15 net28 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 net28 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 net28 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 net24 A0 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN14 net24 A1 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 net24 A1 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN12_2 net24 A0 net28 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y C0 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y C1 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y C1 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y C0 net24 VPW n12 l=1.3e-07 w=7.1e-07
MXP19_2 Y B0 net082__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 net082__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP16 net082 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP19 Y B0 net082 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A0 net092__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net092__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17 net092 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP18 Y A0 net092 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 Y C0 net59__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net59__2 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net59 C1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP20 Y C0 net59 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI222XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1 C0 C1
MXN2 net28 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net28 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net24 A1 net28 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net24 A0 net28 VPW n12 l=1.3e-07 w=3e-07
MXN6 Y C0 net24 VPW n12 l=1.3e-07 w=3e-07
MXN4 Y C1 net24 VPW n12 l=1.3e-07 w=3e-07
MXP14 Y B0 net082 VNW p12 l=1.3e-07 w=3.6e-07
MXP11 net082 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP12 net086 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP13 Y A0 net086 VNW p12 l=1.3e-07 w=3.6e-07
MXP15 Y C0 net59 VNW p12 l=1.3e-07 w=3.6e-07
MXP8 net59 C1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI22X1MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=3.6e-07
MXN0 Y A0 net072 VPW n12 l=1.3e-07 w=3.6e-07
MXN1 net072 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN2 net072 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP0 net22 A1 VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP1 Y A0 net22 VNW p12 l=1.3e-07 w=5.9e-07
MXP2 Y B0 net32 VNW p12 l=1.3e-07 w=5.9e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=5.9e-07
.ends


.SUBCKT OAI22X2MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN3 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN4 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP3 net22 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 Y A0 net22 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y B0 net32 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI22X4MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN3 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN3_2 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN4 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5_2 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4_2 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4_2 Y A0 net22__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP3_2 net22__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP3 net22 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 Y A0 net22 VNW p12 l=1.3e-07 w=8.7e-07
MXP5_2 Y B0 net32__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net32__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y B0 net32 VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI22X8MTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN8 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_2 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_3 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_3 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_4 net072 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_4 net072 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_2 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN7_2 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN7_3 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_3 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN6_4 Y A1 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXN7_4 Y A0 net072 VPW n12 l=1.3e-07 w=7.1e-07
MXP9_2 Y B0 net32__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_2 net32__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8_3 net32__3 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9_3 Y B0 net32__3 VNW p12 l=1.3e-07 w=8.7e-07
MXP9_4 Y B0 net32__4 VNW p12 l=1.3e-07 w=8.7e-07
MXP8_4 net32__4 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y B0 net32 VNW p12 l=1.3e-07 w=8.7e-07
MXP7_2 Y A0 net22__2 VNW p12 l=1.3e-07 w=8.1e-07
MXP6_2 net22__2 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP6_3 net22__3 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7_3 Y A0 net22__3 VNW p12 l=1.3e-07 w=8.1e-07
MXP7_4 Y A0 net22__4 VNW p12 l=1.3e-07 w=8.1e-07
MXP6_4 net22__4 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP6 net22 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP7 Y A0 net22 VNW p12 l=1.3e-07 w=8.1e-07
.ends


.SUBCKT OAI22XLMTR Y VDD VNW VPW VSS A0 A1 B0 B1
MXN6 Y A1 net072 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 Y A0 net072 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 net072 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 net072 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXP3 net22 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP4 Y A0 net22 VNW p12 l=1.3e-07 w=3.6e-07
MXP5 Y B0 net32 VNW p12 l=1.3e-07 w=3.6e-07
MXP8 net32 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2B11X1MTR Y VDD VNW VPW VSS A0 A1N B0 C0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNC2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNC1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y B0 XI1_n2 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB1 XI1_n2 C0 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPC2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPC1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2B11X2MTR Y VDD VNW VPW VSS A0 A1N B0 C0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNC2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNC1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n2 C0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPC2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPC1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B11X4MTR Y VDD VNW VPW VSS A0 A1N B0 C0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNC2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNC1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNC1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNC2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n2__2 C0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y B0 XI1_n2__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n2 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n2 C0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPC2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPC1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPC1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPC2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y C0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B11XLMTR Y VDD VNW VPW VSS A0 A1N B0 C0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNC2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNC1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y B0 XI1_n2 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n2 C0 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPC2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPC1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y C0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2B1X1MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2B1X2MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B1X4MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPB2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B1X8MTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_3 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_3 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_4 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_4 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPB2_2 XI1_p1__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y A0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_3 Y A0 XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_3 XI1_p1__3 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_4 XI1_p1__4 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_4 Y A0 XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B1XLMTR Y VDD VNW VPW VSS A0 A1N B0
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNB2 XI1_n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y B0 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPB2 XI1_p1 A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y A0 XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2B2X1MTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2B2X2MTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B2X4MTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2_2 XI1_p1A__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y A0 XI1_p1A__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_2 XI1_p1B__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y B0 XI1_p1B__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B2X8MTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 A1 A1N VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_3 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_4 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_3 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_3 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_4 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_4 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 A1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA2_2 XI1_p1A__2 A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y A0 XI1_p1A__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y A0 XI1_p1A__3 VNW p12 l=1.3e-07 w=8.1e-07
mXI1_MXPA2_3 XI1_p1A__3 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI1_MXPA2_4 XI1_p1A__4 A1 VDD VNW p12 l=1.3e-07 w=8.1e-07
mXI1_MXPA1_4 Y A0 XI1_p1A__4 VNW p12 l=1.3e-07 w=8.1e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_2 XI1_p1B__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y B0 XI1_p1B__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_3 Y B0 XI1_p1B__3 VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPB2_3 XI1_p1B__3 B1 VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPB2_4 XI1_p1B__4 B1 VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPB1_4 Y B0 XI1_p1B__4 VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2B2XLMTR Y VDD VNW VPW VSS A0 A1N B0 B1
mXI0_MXNA1 A1 A1N VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA2 Y A1 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y A0 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXPA1 A1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 XI1_p1A A1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y A0 XI1_p1A VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y B0 XI1_p1B VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB2 XI1_p1B B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2BB1X1MTR Y VDD VNW VPW VSS A0N A1N B0
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNA2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2BB1X2MTR Y VDD VNW VPW VSS A0N A1N B0
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI1_MXPA2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB1X4MTR Y VDD VNW VPW VSS A0N A1N B0
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA2_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI1_MXPA2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA2_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB1XLMTR Y VDD VNW VPW VSS A0N A1N B0
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI2BB2X1MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=3.3e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=6.2e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI2BB2X2MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB2X4MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_2 XI1_p1__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y B0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB2X8MTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA1_2 nmin1 A1N XI0_n1__2 VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 XI0_n1__2 A0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_2 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_3 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_3 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB1_4 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNB2_4 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA2_2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI0_MXPA1_2 nmin1 A1N VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y nmin1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_2 XI1_p1__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_2 Y B0 XI1_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_3 Y B0 XI1_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_3 XI1_p1__3 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2_4 XI1_p1__4 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1_4 Y B0 XI1_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI2BB2XLMTR Y VDD VNW VPW VSS A0N A1N B0 B1
mXI0_MXNA2 XI0_n1 A0N VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 nmin1 A1N XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB2 XI1_n1 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNB1 XI1_n1 B0 VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y nmin1 XI1_n1 VPW n12 l=1.3e-07 w=3e-07
mXI0_MXPA2 nmin1 A0N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 nmin1 A1N VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPB2 XI1_p1 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPB1 Y B0 XI1_p1 VNW p12 l=1.3e-07 w=3.6e-07
mXI1_MXPA1 Y nmin1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI31X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0
MXN3 n1 A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN2 n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXPA2 net42 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP1 net039 A1 net42 VNW p12 l=1.3e-07 w=6.2e-07
MXP2 Y A0 net039 VNW p12 l=1.3e-07 w=6.2e-07
MXP3 Y B0 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI31X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0
MXN6 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN5 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN4 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXPA2 net42 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP4 net039 A1 net42 VNW p12 l=1.3e-07 w=8.7e-07
MXP5 Y A0 net039 VNW p12 l=1.3e-07 w=8.7e-07
MXP6 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI31X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0
MXN9 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN7_2 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8_2 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9_2 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXNB0_2 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXPA2_2 net42__2 A2 VDD VNW p12 l=1.3e-07 w=8.2e-07
MXP10_2 net039__2 A1 net42__2 VNW p12 l=1.3e-07 w=8.2e-07
MXP11_2 Y A0 net039__2 VNW p12 l=1.3e-07 w=8.2e-07
MXP11 Y A0 net039 VNW p12 l=1.3e-07 w=8.2e-07
MXP10 net039 A1 net42 VNW p12 l=1.3e-07 w=8.2e-07
MXPA2 net42 A2 VDD VNW p12 l=1.3e-07 w=8.2e-07
MXP9 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9_2 Y B0 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI31XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0
MXN6 n1 A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN5 n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXPA2 net42 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP4 net039 A1 net42 VNW p12 l=1.3e-07 w=3.6e-07
MXP5 Y A0 net039 VNW p12 l=1.3e-07 w=3.6e-07
MXP6 Y B0 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI32X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
MXN3 n1 A2 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN4 n1 A1 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN5 n1 A0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN1 Y B0 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXN2 Y B1 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXP1 net59 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP4 net67 A1 net59 VNW p12 l=1.3e-07 w=6.2e-07
MXP5 Y A0 net67 VNW p12 l=1.3e-07 w=6.2e-07
MXP3 Y B0 net55 VNW p12 l=1.3e-07 w=6.2e-07
MXP2 net55 B1 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI32X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
MXN7 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN8 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN6 Y B1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXPA2 net59 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net67 A1 net59 VNW p12 l=1.3e-07 w=8.7e-07
MXP9 Y A0 net67 VNW p12 l=1.3e-07 w=8.7e-07
MXP7 Y B0 net55 VNW p12 l=1.3e-07 w=8.7e-07
MXP6 net55 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI32X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
MXN12 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 n1 A0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 n1 A1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12_2 n1 A2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 Y B1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN10 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN10_2 Y B0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN11_2 Y B1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXP10_2 net59__2 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP13_2 net67__2 A1 net59__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14_2 Y A0 net67__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 Y A0 net67 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 net67 A1 net59 VNW p12 l=1.3e-07 w=8.7e-07
MXP10 net59 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP11_2 net55__2 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP12_2 Y B0 net55__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 Y B0 net55 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 net55 B1 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI32XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1
MXN16 n1 A2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN17 n1 A1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN18 n1 A0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXNB0 Y B0 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 Y B1 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXPA2 net59 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP17 net67 A1 net59 VNW p12 l=1.3e-07 w=3.6e-07
MXP18 Y A0 net67 VNW p12 l=1.3e-07 w=3.6e-07
MXP16 Y B0 net55 VNW p12 l=1.3e-07 w=3.6e-07
MXP15 net55 B1 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OAI33X1MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN4 VSS B2 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXN5 VSS B1 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXN6 VSS B0 n1 VPW n12 l=1.3e-07 w=3.6e-07
MXN2 n1 A0 Y VPW n12 l=1.3e-07 w=3.6e-07
MXN1 n1 A1 Y VPW n12 l=1.3e-07 w=3.6e-07
MXN3 n1 A2 Y VPW n12 l=1.3e-07 w=3.6e-07
MXP1 net77 B2 VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 net73 B1 net77 VNW p12 l=1.3e-07 w=6.2e-07
MXP4 Y B0 net73 VNW p12 l=1.3e-07 w=6.2e-07
MXP6 Y A0 net89 VNW p12 l=1.3e-07 w=6.2e-07
MXP5 net89 A1 net81 VNW p12 l=1.3e-07 w=6.2e-07
MXP2 net81 A2 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OAI33X2MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN10 n1 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN11 n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN12 n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN9 Y A0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN7 Y A1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN8 Y A2 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXP7 net77 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP9 net73 B1 net77 VNW p12 l=1.3e-07 w=8.7e-07
MXP10 Y B0 net73 VNW p12 l=1.3e-07 w=8.7e-07
MXP12 Y A0 net89 VNW p12 l=1.3e-07 w=8.7e-07
MXP11 net89 A1 net81 VNW p12 l=1.3e-07 w=8.7e-07
MXP8 net81 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI33X4MTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN16 n1 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN17 n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN18 n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN18_2 n1 B0 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN17_2 n1 B1 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN16_2 n1 B2 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN15 Y A2 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN13 Y A1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN14 Y A0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN14_2 Y A0 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN13_2 Y A1 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXN15_2 Y A2 n1 VPW n12 l=1.3e-07 w=7.1e-07
MXP14_2 net77__2 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP15_2 net73__2 B1 net77__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP16_2 Y B0 net73__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP16 Y B0 net73 VNW p12 l=1.3e-07 w=8.7e-07
MXP15 net73 B1 net77 VNW p12 l=1.3e-07 w=8.7e-07
MXP14 net77 B2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP13_2 net81__2 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP17_2 net89__2 A1 net81__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18_2 Y A0 net89__2 VNW p12 l=1.3e-07 w=8.7e-07
MXP18 Y A0 net89 VNW p12 l=1.3e-07 w=8.1e-07
MXP17 net89 A1 net81 VNW p12 l=1.3e-07 w=8.7e-07
MXP13 net81 A2 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OAI33XLMTR Y VDD VNW VPW VSS A0 A1 A2 B0 B1 B2
MXN9 n1 B2 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 n1 B1 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN11 n1 B0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN18 Y A0 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 Y A1 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 Y A2 n1 VPW n12 l=1.3e-07 w=1.8e-07
MXP7 net77 B2 VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP8 net73 B1 net77 VNW p12 l=1.3e-07 w=3.6e-07
MXP9 Y B0 net73 VNW p12 l=1.3e-07 w=3.6e-07
MXP11 Y A0 net89 VNW p12 l=1.3e-07 w=3.6e-07
MXP10 net89 A1 net81 VNW p12 l=1.3e-07 w=3.6e-07
MXPA2 net81 A2 VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT OR2X12MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A XI0_p1__3 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p1__3 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 XI0_p1__4 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 ny A XI0_p1__4 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR2X1MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=3.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OR2X2MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR2X4MTR Y VDD VNW VPW VSS A B
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR2X6MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR2X8MTR Y VDD VNW VPW VSS A B
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA2_2 XI0_p1__2 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p1__2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 ny A XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p1 B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X12MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_3 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2_3 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3_2 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3_3 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_5 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_6 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_4 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_5 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_4 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_5 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_5 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_6 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X1MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=4.8e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=4.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OR3X2MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=3e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X4MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_2 ny A XI0_p2__2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X6MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA3_2 XI0_p1__2 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2_2 XI0_p2__2 B XI0_p1__2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1_2 ny A XI0_p2__2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=7.8e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR3X8MTR Y VDD VNW VPW VSS A B C
mXI0_MXNA1 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1_2 ny A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA2_2 ny B VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA3_2 ny C VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI1_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXPA1 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 ny A XI0_p2 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_2 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA2_3 XI0_p2 B XI0_p1 VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_2 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA3_3 XI0_p1 C VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X12MTR Y VDD VNW VPW VSS A B C D
MXN14 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN14_2 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN14_3 net43 D VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN14_4 net43 D VSS VPW n12 l=1.3e-07 w=3e-07
MXN13 net43 C VSS VPW n12 l=1.3e-07 w=3e-07
MXN13_2 net43 C VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN13_3 net43 C VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN13_4 net43 C VSS VPW n12 l=1.3e-07 w=3e-07
MXN13_5 net43 C VSS VPW n12 l=1.3e-07 w=3e-07
MXN13_6 net43 C VSS VPW n12 l=1.3e-07 w=3.1e-07
MXN12 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN12_2 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN12_3 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA_2 net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA_3 net43 A VSS VPW n12 l=1.3e-07 w=3.1e-07
MXNA_4 net43 A VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI0_MXNA1_2 Y net43 VSS VPW n12 l=1.3e-07 w=3.5e-07
mXI0_MXNA1_3 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_5 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_6 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_7 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 net62 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_3 net62 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_4 net62 D VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_5 net62 D VDD VNW p12 l=1.3e-07 w=1.23e-06
MXP20 net66 C net62 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_2 net66 C net62 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_3 net66 C net62 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_4 net66 C net62 VNW p12 l=1.3e-07 w=8.7e-07
MXP20_5 net66 C net62 VNW p12 l=1.3e-07 w=1.23e-06
MXP21 net70 B net66 VNW p12 l=1.3e-07 w=1.23e-06
MXP21_2 net70 B net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP21_3 net70 B net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP21_4 net70 B net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP21_5 net70 B net66 VNW p12 l=1.3e-07 w=8.7e-07
MXP22 net43 A net70 VNW p12 l=1.3e-07 w=8.7e-07
MXP22_2 net43 A net70 VNW p12 l=1.3e-07 w=8.7e-07
MXP22_3 net43 A net70 VNW p12 l=1.3e-07 w=8.7e-07
MXP22_4 net43 A net70 VNW p12 l=1.3e-07 w=8.7e-07
MXP22_5 net43 A net70 VNW p12 l=1.3e-07 w=1.23e-06
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_5 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_6 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X1MTR Y VDD VNW VPW VSS A B C D
MXNA net43 A VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN0 net43 B VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN1 net43 C VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN2 net43 D VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP7 net43 A net70 VNW p12 l=1.3e-07 w=4.9e-07
MXP6 net70 B net66 VNW p12 l=1.3e-07 w=4.9e-07
MXP5 net66 C net62 VNW p12 l=1.3e-07 w=4.9e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT OR4X2MTR Y VDD VNW VPW VSS A B C D
MXNA net43 A VSS VPW n12 l=1.3e-07 w=3e-07
MXN3 net43 B VSS VPW n12 l=1.3e-07 w=3e-07
MXN4 net43 C VSS VPW n12 l=1.3e-07 w=3e-07
MXN5 net43 D VSS VPW n12 l=1.3e-07 w=3e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP10 net43 A net70 VNW p12 l=1.3e-07 w=7.9e-07
MXP9 net70 B net66 VNW p12 l=1.3e-07 w=7.9e-07
MXP8 net66 C net62 VNW p12 l=1.3e-07 w=7.9e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X4MTR Y VDD VNW VPW VSS A B C D
MXN8 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN7 net43 C VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN6 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_2 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP11 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP11_2 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP12 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP12_2 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP13 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP13_2 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X6MTR Y VDD VNW VPW VSS A B C D
MXNA net43 A VSS VPW n12 l=1.3e-07 w=4.6e-07
MXNA_2 net43 A VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN9 net43 B VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN9_2 net43 B VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN10 net43 C VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN10_2 net43 C VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN11 net43 D VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN11_2 net43 D VSS VPW n12 l=1.3e-07 w=4.6e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP16 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP16_2 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP16_3 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP15 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP15_2 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP15_3 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP14 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP14_2 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP14_3 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_2 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_3 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT OR4X8MTR Y VDD VNW VPW VSS A B C D
MXN14 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN14_2 net43 D VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN13 net43 C VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN13_2 net43 C VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN12 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN12_2 net43 B VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXNA_2 net43 A VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI0_MXNA1 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_2 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_3 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1_4 Y net43 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_2 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_3 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP0_4 net62 D VDD VNW p12 l=1.3e-07 w=8e-07
MXP17 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP17_2 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP17_3 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP17_4 net66 C net62 VNW p12 l=1.3e-07 w=8e-07
MXP18 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP18_2 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP18_3 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP18_4 net70 B net66 VNW p12 l=1.3e-07 w=8e-07
MXP19 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP19_2 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP19_3 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
MXP19_4 net43 A net70 VNW p12 l=1.3e-07 w=8e-07
mXI0_MXPA1 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_2 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_3 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1_4 Y net43 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX12MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=3.2e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=5e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=4.5e-07
MXN3_2 nmin OE net31 VPW n12 l=1.3e-07 w=4.5e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN0_3 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_5 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_6 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=3.9e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=6.5e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=3e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=8e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP0_3 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_5 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX16MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=4.1e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN3_2 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=6.9e-07
MXN0_3 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_5 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_6 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_7 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_8 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=8e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=5.2e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=8.6e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_3 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_5 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_7 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_8 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX1MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT TBUFX20MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=5.2e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=4.4e-07
MXN4_2 net31 nmen VSS VPW n12 l=1.3e-07 w=4.4e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=6.5e-07
MXN3_2 nmin OE net31 VPW n12 l=1.3e-07 w=6.5e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_3 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_4 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_5 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_6 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_7 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_8 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_9 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_10 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP4_2 nmin OE VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=8e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=8e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_3 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_4 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_5 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_7 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_8 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_9 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_10 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX24MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=6.3e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=5.2e-07
MXN4_2 net31 nmen VSS VPW n12 l=1.3e-07 w=5.2e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN3_2 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN3_3 nmin OE net31 VPW n12 l=1.3e-07 w=6.1e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_3 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_4 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN0_5 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_5 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_6 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_7 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_8 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_9 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_10 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_11 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2_12 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=7.7e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP5_3 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP5_4 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=6.6e-07
MXP4_2 nmin OE VDD VNW p12 l=1.3e-07 w=6.6e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_3 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_4 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP0_5 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_5 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_6 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_7 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_8 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_9 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_10 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_11 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2_12 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT TBUFX2MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=3e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.2e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=3.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=7e-07
.ends


.SUBCKT TBUFX3MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=2.3e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=5.3e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=3e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=6.6e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=6.6e-07
.ends


.SUBCKT TBUFX4MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=3e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=3.6e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
.ends


.SUBCKT TBUFX6MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=1.9e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=3e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=3.7e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=7.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.6e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=3e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=5.6e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=8.7e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=7.9e-07
.ends


.SUBCKT TBUFX8MTR Y VDD VNW VPW VSS A OE
mX_g0_MXNA1 nmen OE VSS VPW n12 l=1.3e-07 w=3e-07
MXN4 net31 nmen VSS VPW n12 l=1.3e-07 w=3.6e-07
MXN3 nmin OE net31 VPW n12 l=1.3e-07 w=6.4e-07
MXN0 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN0_2 net31 A VSS VPW n12 l=1.3e-07 w=6.1e-07
MXN2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_2 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_3 Y net31 VSS VPW n12 l=1.3e-07 w=6.5e-07
MXN2_4 Y net31 VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXPA1 nmen OE VDD VNW p12 l=1.3e-07 w=3e-07
MXP4 nmin OE VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP5 nmin nmen net31 VNW p12 l=1.3e-07 w=3e-07
MXP5_2 nmin nmen net31 VNW p12 l=1.3e-07 w=5e-07
MXP0 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP0_2 nmin A VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_2 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_3 Y nmin VDD VNW p12 l=1.3e-07 w=8e-07
MXP2_4 Y nmin VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends




.SUBCKT XNOR2X1MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=3e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=3e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=3.8e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=3.8e-07
.ends


.SUBCKT XNOR2X2MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=5.7e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=7.2e-07
.ends


.SUBCKT XNOR2X4MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_2 Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_2 Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN_2 Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=7.6e-07
mXI2_MXPOEN_2 Y A nb VNW p12 l=1.3e-07 w=7.6e-07
.ends


.SUBCKT XNOR2X8MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_3 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_4 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=5.3e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_2 Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_3 Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_4 Y A bb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_2 Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_3 Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_4 Y na nb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_3 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_4 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN_2 Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN_3 Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN_4 Y na bb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=7.6e-07
mXI2_MXPOEN_2 Y A nb VNW p12 l=1.3e-07 w=7.6e-07
mXI2_MXPOEN_3 Y A nb VNW p12 l=1.3e-07 w=7.6e-07
mXI2_MXPOEN_4 Y A nb VNW p12 l=1.3e-07 w=7.6e-07
.ends


.SUBCKT XNOR2XLMTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE Y A bb VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE Y na nb VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN Y na bb VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN Y A nb VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT XNOR3X1MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI52_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=3.7e-07
mXI53_MXNOE ny na bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI52_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=4.6e-07
mXI53_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT XNOR3X2MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=6e-07
mXI48_MXNOE ny na bnc VPW n12 l=1.3e-07 w=5.5e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI4_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI8_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=7.2e-07
mXI48_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=7.2e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XNOR3X4MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_2 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny na bnc VPW n12 l=1.3e-07 w=5.5e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.6e-07
mXI7_MXPA1_2 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI8_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=7.2e-07
mXI4_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=7.2e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XNOR3X8MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_2 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_3 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_4 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny na bnc VPW n12 l=1.3e-07 w=5.5e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.6e-07
mXI7_MXPA1_2 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.6e-07
mXI7_MXPA1_3 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI7_MXPA1_4 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI8_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=7.2e-07
mXI4_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=7.2e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XNOR3XLMTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=4.8e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=2e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=3e-07
mXI8_MXNOE ny C nbnc VPW n12 l=1.3e-07 w=3e-07
mXI4_MXNOE ny na bnc VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=5.8e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=5.8e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=4.8e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=1.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI8_MXPOEN ny na nbnc VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN ny C bnc VNW p12 l=1.3e-07 w=5.8e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT XOR2X1MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=3e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=3e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=3.8e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=3.8e-07
.ends


.SUBCKT XOR2X2MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=5.7e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=7.2e-07
.ends


.SUBCKT XOR2X3MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=4.5e-07
mXI2_MXNOE_2 Y A nb VPW n12 l=1.3e-07 w=4.5e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI4_MXNOE_2 Y na bb VPW n12 l=1.3e-07 w=4.5e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=4.7e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=5.7e-07
mXI2_MXPOEN_2 Y na nb VNW p12 l=1.3e-07 w=5.7e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=5.7e-07
mXI4_MXPOEN_2 Y A bb VNW p12 l=1.3e-07 w=5.7e-07
.ends


.SUBCKT XOR2X4MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_2 Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_2 Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN_2 Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=7.6e-07
mXI4_MXPOEN_2 Y A bb VNW p12 l=1.3e-07 w=7.6e-07
.ends


.SUBCKT XOR2X8MTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_2 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_3 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI1_MXNA1_4 nb B VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_2 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_3 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNA1_4 bb nb VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI0_MXNA1_2 na A VSS VPW n12 l=1.3e-07 w=5.2e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_2 Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_3 Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI2_MXNOE_4 Y A nb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_2 Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_3 Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE_4 Y na bb VPW n12 l=1.3e-07 w=6e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_2 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_3 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI1_MXPA1_4 nb B VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_2 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_3 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPA1_4 bb nb VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI0_MXPA1_2 na A VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN_2 Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN_3 Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI2_MXPOEN_4 Y na nb VNW p12 l=1.3e-07 w=6.1e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=7.6e-07
mXI4_MXPOEN_2 Y A bb VNW p12 l=1.3e-07 w=7.6e-07
mXI4_MXPOEN_3 Y A bb VNW p12 l=1.3e-07 w=7.6e-07
mXI4_MXPOEN_4 Y A bb VNW p12 l=1.3e-07 w=7.6e-07
.ends


.SUBCKT XOR2XLMTR Y VDD VNW VPW VSS A B
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 bb nb VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 na A VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXNOE Y A nb VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE Y na bb VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI3_MXPA1 bb nb VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI0_MXPA1 na A VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI2_MXPOEN Y na nb VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN Y A bb VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT XOR3X1MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=3.7e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=4.6e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT XOR3X2MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=7.4e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XOR3X4MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_2 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI7_MXPA1_2 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=7.4e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XOR3X8MTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=6e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=4.5e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=4e-07
mXI5_MXNA1_2 bc nc VSS VPW n12 l=1.3e-07 w=3.2e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_2 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_3 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI7_MXNA1_4 nbnc bnc VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=6e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=5.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=2.6e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_2 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_3 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI9_MXNA1_4 Y ny VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=7.6e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=7.2e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4e-07
mXI5_MXPA1_2 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI7_MXPA1_2 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI7_MXPA1_3 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.5e-07
mXI7_MXPA1_4 nbnc bnc VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=7.4e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3.2e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_2 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_3 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI9_MXPA1_4 Y ny VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT XOR3XLMTR Y VDD VNW VPW VSS A B C
mXI2_MXNA1 nc A VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI3_MXNOE bnc B nc VPW n12 l=1.3e-07 w=4.8e-07
mXI6_MXNOE bnc nb bc VPW n12 l=1.3e-07 w=3.7e-07
mXI5_MXNA1 bc nc VSS VPW n12 l=1.3e-07 w=3.7e-07
mXI1_MXNA1 nb B VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI7_MXNA1 nbnc bnc VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI8_MXNOE ny na nbnc VPW n12 l=1.3e-07 w=2.1e-07
mXI4_MXNOE ny C bnc VPW n12 l=1.3e-07 w=4.8e-07
mXI0_MXNA1 na C VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI9_MXNA1 Y ny VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI2_MXPA1 nc A VDD VNW p12 l=1.3e-07 w=5.8e-07
mXI3_MXPOEN bnc nb nc VNW p12 l=1.3e-07 w=5.8e-07
mXI6_MXPOEN bnc B bc VNW p12 l=1.3e-07 w=4.8e-07
mXI5_MXPA1 bc nc VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI1_MXPA1 nb B VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPA1 nbnc bnc VDD VNW p12 l=1.3e-07 w=2.5e-07
mXI8_MXPOEN ny C nbnc VNW p12 l=1.3e-07 w=2.5e-07
mXI4_MXPOEN ny na bnc VNW p12 l=1.3e-07 w=5.7e-07
mXI0_MXPA1 na C VDD VNW p12 l=1.3e-07 w=3e-07
mXI9_MXPA1 Y ny VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends

