* 
* No part of this file can be released without the consent of SMIC.
*
* Note: SMIC recommends that users set VNTOL=1E-9 at .option for more smooth convergence.
******************************************************************************************
* 0.11um Mixed Signal 1P8M with MIM Salicide 1.2V/3.3V RF SPICE Model (for HSPICE only)  *
******************************************************************************************
*
* Release version    : 1.14
*
* Release date       : 03/30/2016
*
* Simulation tool    : Synopsys Star-HSPICE version 2006.09
*
*  Resistor   :
*        *------------------------------------------------------------------* 
*        |                 |                Resistor subckt                 |
*        *==================================================================*
*        | N+ poly SAB     |    rnposab_ckt_rf     |    rnposab_ckt_rf_3t   |
*        *------------------------------------------------------------------*
*        | p+ poly SAB     |    rpposab_ckt_rf     |    rpposab_ckt_rf_3t   |
*        *------------------------------------------------------------------*
*        | HRP poly        |    rhrpo_ckt_rf      |     rhrpo_ckt_rf_3t     |
*        *------------------------------------------------------------------*

******************************                                   
*Non-silicide N+ Poly resistor               
******************************                      
.subckt rnposab_ckt_rf port1 port2 l=l_rf w=w_rf devt='temper' mismod_res_rf=0
.param  
*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = '1/sqrt(weff*leff)'
+arsh = 1.0E-05

+rsh       = '275.50+DRSH_RNPOSAB_RF+rshmis'   rtc1     = -9.93E-04     rtc2  = 1.07E-06    
+dw        = '1.68E-08-2.7E-9+DDW_RNPOSAB_RF'  dl       = -1.33e-7
+jc1a      = 3.04E-05                jc1b     = -3.29E-09 
+jc2a      = -1.18E-08               jc2b     = -2.99E-13
+rvc1      = 'jc1a+jc1b/l'           rvc2     = '(jc2a+jc2b/l)/l' 
+weff      = 'w*0.9-2*dw'                leff     = 'l*0.9-2*dl'
+tcoef     = '1.0+(devt-25.0)*(rtc1+rtc2*(devt-25.0))' 
*RF component value
+Ls_rf      = 'max((0.007035*pwr(w*0.9*1e6+0.19294,1.0366)*(0.135+pwr((l*0.9)/(w*0.9)+0.2,-2.221*pwr(w*0.9*1e6,-0.1078)+4.864)))*1e-9,1e-12)'
+Cf_rf      = 'max((0.08566*pwr(w*0.9*1e6+0.2,-0.8872)*(0.006+pwr((l*0.9)/(w*0.9)+0.0202,0.2368*pwr(w*0.9*1e6,-1.7352)-3.026)))*1e-15,1e-18)'
+Rsub_rf    = 'max(165.3+2389.6*pwr(w*0.9*1e6,-0.9242)+174.3*pwr(w*0.9*1e6+2.0705,4)*pwr(l*0.9*1e6+0.02666,-0.4314*pwr(w*0.9*1e6,1.2708)-1.916),1e-5)'
+Csub_rf    = 'max((0.03194*pwr(w*0.9*1e6+0.2,1.5946)*(6.783+pwr(l*0.9*w*0.9*1e12+0.13226,-0.347*pwr(w*0.9*1e6,0.87)+1.4215)))*1e-15,1e-18)'
+Cox_rf     = 'max((0.01085*pwr(w*0.9*1e6+0.2,0.5126)*(10+pwr(l*0.9*w*0.9*1e12+0.4065,0.9025*pwr(w*0.9*1e6,-1.7592)+1.0813)))*1e-15,1e-18)'
+Rs2_rf     = 'max(0.39+0.44455*pwr(w*0.9*1e6+0.13192,-0.3454)*(0.155+exp(5+0.06201*(pwr(w*0.9*1e6,1.26)+3.094)*(l*0.9)/(w*0.9))),1e-5)'
* equivalent circuit
Ls 1 port2    l=Ls_rf
Cf port1 1    c=Cf_rf
Rs port1 1    r='rsh*leff/weff*tcoef*max(1.0+rvc1*abs(v(port1,1))+rvc2*v(port1,1)*v(port1,1),0.834)'
Rs2 1 port2   r=Rs2_rf
Rsub1 2 0     r=Rsub_rf
Csub1 2 0     c=Csub_rf
Cox1 port1 2  c=Cox_rf
Rsub2 3 0     r=Rsub_rf
Csub2 3 0     c=Csub_rf
Cox2 port2 3  c=Cox_rf
.ends rnposab_ckt_rf
***************************************************
*Non-silicide N+ Poly resistor (three terminal)              
***************************************************
.subckt rnposab_ckt_rf_3t port1 port2 pwell l=l_rf w=w_rf devt='temper' mismod_res_rf=0
.param  
*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = '1/sqrt(weff*leff)'
+arsh = 1.0E-05

+rsh       = '275.50+DRSH_RNPOSAB_RF+rshmis'   rtc1     = -9.93E-04     rtc2  = 1.07E-06    
+dw        = '1.68E-08-2.7E-9+DDW_RNPOSAB_RF'  dl       = -1.33e-7
+jc1a      = 3.04E-05                jc1b     = -3.29E-09 
+jc2a      = -1.18E-08               jc2b     = -2.99E-13
+rvc1      = 'jc1a+jc1b/l'           rvc2     = '(jc2a+jc2b/l)/l' 
+weff      = 'w*0.9-2*dw'                leff     = 'l*0.9-2*dl'
+tcoef     = '1.0+(devt-25.0)*(rtc1+rtc2*(devt-25.0))' 
*RF component value
+Ls_rf      = 'max((0.007035*pwr(w*0.9*1e6+0.19294,1.0366)*(0.135+pwr((l*0.9)/(w*0.9)+0.2,-2.221*pwr(w*0.9*1e6,-0.1078)+4.864)))*1e-9,1e-12)'
+Cf_rf      = 'max((0.08566*pwr(w*0.9*1e6+0.2,-0.8872)*(0.006+pwr((l*0.9)/(w*0.9)+0.0202,0.2368*pwr(w*0.9*1e6,-1.7352)-3.026)))*1e-15,1e-18)'
+Rsub_rf    = 'max(165.3+2389.6*pwr(w*0.9*1e6,-0.9242)+174.3*pwr(w*0.9*1e6+2.0705,4)*pwr(l*0.9*1e6+0.02666,-0.4314*pwr(w*0.9*1e6,1.2708)-1.916),1e-5)'
+Csub_rf    = 'max((0.03194*pwr(w*0.9*1e6+0.2,1.5946)*(6.783+pwr(l*0.9*w*0.9*1e12+0.13226,-0.347*pwr(w*0.9*1e6,0.87)+1.4215)))*1e-15,1e-18)'
+Cox_rf     = 'max((0.01085*pwr(w*0.9*1e6+0.2,0.5126)*(10+pwr(l*0.9*w*0.9*1e12+0.4065,0.9025*pwr(w*0.9*1e6,-1.7592)+1.0813)))*1e-15,1e-18)'
+Rs2_rf     = 'max(0.39+0.44455*pwr(w*0.9*1e6+0.13192,-0.3454)*(0.155+exp(5+0.06201*(pwr(w*0.9*1e6,1.26)+3.094)*(l*0.9)/(w*0.9))),1e-5)'
* equivalent circuit
Ls 1 port2    l=Ls_rf
Cf port1 1    c=Cf_rf
Rs port1 1    r='rsh*leff/weff*tcoef*max(1.0+rvc1*abs(v(port1,1))+rvc2*v(port1,1)*v(port1,1),0.834)'
Rs2 1 port2   r=Rs2_rf
Rsub1 2 pwell     r=Rsub_rf
Csub1 2 pwell     c=Csub_rf
Cox1 port1 2  c=Cox_rf
Rsub2 3 pwell     r=Rsub_rf
Csub2 3 pwell     c=Csub_rf
Cox2 port2 3  c=Cox_rf
.ends rnposab_ckt_rf_3T
******************************                                   
*Non-silicide P+ Poly resistor               
******************************                      
.subckt rpposab_ckt_rf port1 port2 l=l_rf w=w_rf devt='temper' mismod_res_rf=0
.param
*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = '1/sqrt(weff*leff)'
+arsh = 3.4E-06

+rsh       = '321.5+DRSH_RPPOSAB_RF+rshmis'    rtc1     = -5.75E-05     rtc2  = 6.10E-07    
+dw        = '1.28E-08-2.7E-9+DDW_RPPOSAB_RF'  dl       = -2.68e-7
*+vc1      = -5.07E-05               vc2      = -7.96E-05 
+jc1a      = 2.16E-05                jc1b     = -1.77E-9 
+jc2a      = -7.61E-10               jc2b     = -1.79E-14
+rvc1      = 'jc1a+jc1b/l'           rvc2     = '(jc2a+jc2b/l)/l' 
+weff      = 'w*0.9-2*dw'                leff     = 'l*0.9-2*dl'
+tcoef     = '1.0+(devt-25.0)*(rtc1+rtc2*(devt-25.0))'  
*RF component value
+Ls_rf      = 'max(((0.0129*w*1e6+0.0006)*pwr(l/w,2.3758*pwr(w*1e6,0.1048)))*1e-9,1e-12)'
+Cf_rf      = 'max((0.8913*pwr(l/w,-1.1526))*1e-15,1e-18)'
+Rsub_rf    = 'max(71.885*l/w + 70.958,1e-3)'
+Csub_rf    = 'max((1.5*pwr(l/w,0.4337))*1e-15,1e-18)'
+Cox_rf     = 'max((0.046*w*l*1e12+1.5358)*1e-15,1e-18)'
+Rs2_rf     = 'max(2000*l/w,1e-5)'
* equivalent circuit
Ls 1 port2    l=Ls_rf
Cf port1 1    c=Cf_rf
Rs port1 1    r='rsh*leff/weff*tcoef*max(1.0+rvc1*abs(v(port1,1))+rvc2*v(port1,1)*v(port1,1),0.890)'
Rs2 1 port2   r=Rs2_rf
Cf2   port1 4 c='Cf_rf*0.1'
Rs3   4 port2 r='Rs2_rf*10'
Rsub1 2 0     r=Rsub_rf
Csub1 2 0     c=Csub_rf
Cox1 port1 2  c=Cox_rf
Rsub2 3 0     r=Rsub_rf
Csub2 3 0     c=Csub_rf
Cox2 port2 3  c=Cox_rf
.ends rpposab_ckt_rf
************************************************ 
*Non-silicide P+ Poly resistor (three terminal)
************************************************ 
.subckt rpposab_ckt_rf_3t port1 port2 pwell l=l_rf w=w_rf devt='temper' mismod_res_rf=0
.param
*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = '1/sqrt(weff*leff)'
+arsh = 3.4E-06

+rsh       = '321.5+DRSH_RPPOSAB_RF+rshmis'    rtc1     = -5.75E-05     rtc2  = 6.10E-07    
+dw        = '1.28E-08-2.7E-9+DDW_RPPOSAB_RF'  dl       = -2.68e-7
*+vc1      = -5.07E-05               vc2      = -7.96E-05 
+jc1a      = 2.16E-05                jc1b     = -1.77E-9 
+jc2a      = -7.61E-10               jc2b     = -1.79E-14
+rvc1      = 'jc1a+jc1b/l'           rvc2     = '(jc2a+jc2b/l)/l' 
+weff      = 'w*0.9-2*dw'                leff     = 'l*0.9-2*dl'
+tcoef     = '1.0+(devt-25.0)*(rtc1+rtc2*(devt-25.0))'  
*RF component value
+Ls_rf      = 'max(((0.0129*w*1e6+0.0006)*pwr(l/w,2.3758*pwr(w*1e6,0.1048)))*1e-9,1e-12)'
+Cf_rf      = 'max((0.8913*pwr(l/w,-1.1526))*1e-15,1e-18)'
+Rsub_rf    = 'max(71.885*l/w + 70.958,1e-3)'
+Csub_rf    = 'max((1.5*pwr(l/w,0.4337))*1e-15,1e-18)'
+Cox_rf     = 'max((0.046*w*l*1e12+1.5358)*1e-15,1e-18)'
+Rs2_rf     = 'max(2000*l/w,1e-5)'
* equivalent circuit
Ls 1 port2    l=Ls_rf
Cf port1 1    c=Cf_rf
Rs port1 1    r='rsh*leff/weff*tcoef*max(1.0+rvc1*abs(v(port1,1))+rvc2*v(port1,1)*v(port1,1),0.890)'
Rs2 1 port2   r=Rs2_rf
Cf2   port1 4 c='Cf_rf*0.1'
Rs3   4 port2 r='Rs2_rf*10'
Rsub1 2 pwell     r=Rsub_rf
Csub1 2 pwell     c=Csub_rf
Cox1 port1 2  c=Cox_rf
Rsub2 3 pwell     r=Rsub_rf
Csub2 3 pwell     c=Csub_rf
Cox2 port2 3  c=Cox_rf
.ends rpposab_ckt_rf_3t

*********************************                                   
* Non-Silicide HR Poly resistor *               
*********************************                      
.subckt rhrpo_ckt_rf port1 port2 l=l_rf w=w_rf mismod_res_rf=0
.param
*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = '1/sqrt(weff*l*0.9)'
+arsh = 1.55E-05
*****base model parameter*****  
+rsh      = '963+drsh_rhrpo_rf+rshmis'
+rtc1     = -6.77E-04                    rtc2   = 2.08E-06
+dw       = '2.27E-08-2.7E-9+ddw_rhrpo_rf'
+rint0 = 2.08E-4                    rint1 = 0
+rinttc1 = -6.46E-04                rinttc2 = -1.12E-06
+jc1a = 8.89E-05                    jc1b = -4.49E-09
+jc2a = -2.53E-09                   jc2b = -6.64E-14
+rintjc1a = 0.365                   rintjc1b = 1.45E+3
+rintjc2a = -13.1689                rintjc2b = -1.52E+7
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+rvc1 = 'jc1a + jc1b / (l*0.9)'           rvc2 = '(jc2a + jc2b / (l*0.9)) / (l*0.9)'
+weff = 'w*0.9-2*dw'
+rintvc1 = 'rintjc1a + rintjc1b * weff'  rintvc2 = 'rintjc2a + rintjc2b * weff'
+rinttcoef(temper) = '1.0+(temper-25.0)*(rinttc1+rinttc2*(temper-25.0))'
+Ls_rf	  = 'max((4.246819E-02*pwr(w*1e6,-9.933603E-01)+0.00426)*pwr(l*1e6,(4.312050E-01*pwr(w*1e6,-5.234278E-01)+2.61))*0.9*1e-9, 1e-13)'
+Cf_rf	  = 'max(((8.2020E-04*pwr(w*1e6,1.9584)+0.022)*l*1e6+0.16284)*(9.0016*pwr(l*1e6,-0.5239))*1e-15,1e-18)'
+Rs2_rf	  = 'max(1445.2*pwr(l/w,2.5309),1e-3)'
+Rsub_rf  = 'max((210.2*(l/w)-127.15)*(1.01-0.0059*exp(0.0659*l/w)), 1e-3)'
+Csub_rf  = 'max((0.01*w*l*1e12+1.21)*(0.6274*exp(0.0077*l*1e6))*1e-15,1e-18)'
+Cox_rf   = 'max((0.0512*w*l*1e12-0.5)*1.629*pwr(w*1e6,-0.2921)*1e-15, 1e-18)'
Ls_rf 1 port2    Ls_rf 
Cf_rf port1 1    Cf_rf
*Rinta_rf port1 na '(rint0/weff+rint1/(weff*weff))*rinttcoef(temper)*max(1.0+rintvc1*abs(v(port1,na))+rintvc2*v(port1,na)*v(port1,na), 0.82)'
Rinta_rf port1 na '(rint0/weff+rint1/(weff*weff))*rinttcoef(temper)*max(min(1.0+rintvc1*abs(v(port1,na))+rintvc2*v(port1,na)*v(port1,na),1.5),0.5)'
*Rs_rf na nb    'rsh*l/weff*tcoef(temper)*max(1.0+rvc1*abs(v(na,nb))+rvc2*v(na,nb)*v(na,nb),0.89)'
Rs_rf na nb 'rsh*(l*0.9)/weff*tcoef(temper)*max(min(1.0+rvc1*abs(v(na,nb))+rvc2*v(na,nb)*v(na,nb),1.5),0.5)'
*Rintb_rf nb 1 '(rint0/weff+rint1/(weff*weff))*rinttcoef(temper)*max(1.0+rintvc1*abs(v(nb,1))+rintvc2*v(nb,1)*v(nb,1), 0.82)'
Rintb_rf nb 1 '(rint0/weff+rint1/(weff*weff))*rinttcoef(temper)*max(min(1.0+rintvc1*abs(v(nb,1))+rintvc2*v(nb,1)*v(nb,1),1.5),0.5)'
Rs2_rf 1 port2   Rs2_rf
Cf2_rf port1 4   '0.1*Cf_rf'
Rs3_rf 4 port2   '10*Rs2_rf'
Rsub1_rf 2 0     Rsub_rf
Csub1_rf 2 0     Csub_rf
Cox1_rf port1 2  Cox_rf
Rsub2_rf 3 0     Rsub_rf
Csub2_rf 3 0     Csub_rf
Cox2_rf port2 3  Cox_rf 
.ends rhrpo_ckt_rf
**********************************************                                   
* Non-Silicide HR Poly resistor (3-terminal) *               
**********************************************                      
.subckt rhrpo_ckt_rf_3t port1 port2 B l=l_rf w=w_rf mismod_res_rf=0
.param
*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = '1/sqrt(weff*l*0.9)'
+arsh = 1.55E-05
*****base model parameter*****  
+rsh      = '963+drsh_rhrpo_rf_3t+rshmis'
+rtc1     = -6.77E-04                    rtc2   = 2.08E-06
+dw       = '2.27E-08-2.7E-9+ddw_rhrpo_rf_3t'
+rint0 = 2.08E-4                    rint1 = 0
+rinttc1 = -6.46E-04                rinttc2 = -1.12E-06
+jc1a = 8.89E-05                    jc1b = -4.49E-09
+jc2a = -2.53E-09                   jc2b = -6.64E-14
+rintjc1a = 0.365                   rintjc1b = 1.45E+3
+rintjc2a = -13.1689                rintjc2b = -1.52E+7
+tcoef(temper)     = '1.0+(temper-25.0)*(rtc1+rtc2*(temper-25.0))' 
+rvc1 = 'jc1a + jc1b / (l*0.9)'           rvc2 = '(jc2a + jc2b / (l*0.9)) / (l*0.9)'
+weff = 'w*0.9-2*dw'
+rintvc1 = 'rintjc1a + rintjc1b * weff'  rintvc2 = 'rintjc2a + rintjc2b * weff'
+rinttcoef(temper) = '1.0+(temper-25.0)*(rinttc1+rinttc2*(temper-25.0))'
+Ls_rf	  = 'max((4.246819E-02*pwr(w*1e6,-9.933603E-01)+0.00426)*pwr(l*1e6,(4.312050E-01*pwr(w*1e6,-5.234278E-01)+2.61))*0.9*1e-9, 1e-13)'
+Cf_rf	  = 'max(((8.2020E-04*pwr(w*1e6,1.9584)+0.022)*l*1e6+0.16284)*(9.0016*pwr(l*1e6,-0.5239))*1e-15,1e-18)'
+Rs2_rf	  = 'max(1445.2*pwr(l/w,2.5309),1e-3)'
+Rsub_rf  = 'max((210.2*(l/w)-127.15)*(1.01-0.0059*exp(0.0659*l/w)), 1e-3)'
+Csub_rf  = 'max((0.01*w*l*1e12+1.21)*(0.6274*exp(0.0077*l*1e6))*1e-15,1e-18)'
+Cox_rf   = 'max((0.0512*w*l*1e12-0.5)*1.629*pwr(w*1e6,-0.2921)*1e-15, 1e-18)'
Ls_rf 1 port2    Ls_rf 
Cf_rf port1 1    Cf_rf
Rinta_rf port1 na '(rint0/weff+rint1/(weff*weff))*rinttcoef(temper)*max(min(1.0+rintvc1*abs(v(port1,na))+rintvc2*v(port1,na)*v(port1,na),1.5),0.5)'
Rs_rf na nb 'rsh*(l*0.9)/weff*tcoef(temper)*max(min(1.0+rvc1*abs(v(na,nb))+rvc2*v(na,nb)*v(na,nb),1.5),0.5)'
Rintb_rf nb 1 '(rint0/weff+rint1/(weff*weff))*rinttcoef(temper)*max(min(1.0+rintvc1*abs(v(nb,1))+rintvc2*v(nb,1)*v(nb,1),1.5),0.5)'
Rs2_rf 1 port2   Rs2_rf
Cf2_rf port1 4   '0.1*Cf_rf'
Rs3_rf 4 port2   '10*Rs2_rf'
Rsub1_rf 2 B     Rsub_rf
Csub1_rf 2 B     Csub_rf
Cox1_rf port1 2  Cox_rf
Rsub2_rf 3 B     Rsub_rf
Csub2_rf 3 B     Csub_rf
Cox2_rf port2 3  Cox_rf 
.ends rhrpo_ckt_rf_3t


