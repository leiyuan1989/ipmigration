.model mn15 nmos4 l=1 w=1 n=1
.model mp15 pmos4 l=1 w=1 n=1