****Sub-Circuit for CLKLAHAQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHAQHSV1 CK E ECK BC VDD VSS
MM51 s c VSS VPW N12LL W=200.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=200.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=260.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=200.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM0 ten BC VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=220.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=320.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=260.00n L=60.00n
MM45 s c nt21 VNW P12LL W=540.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=540.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=500.00n L=60.00n
MM1 ten BC VDD VNW P12LL W=300.00n L=60.00n
MM54 nt21 pm VDD VNW P12LL W=540.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=330.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=460.00n L=60.00n
MM39 pm cn nt11 VNW P12LL W=500.00n L=60.00n
.ENDS CLKLAHAQHSV1
****Sub-Circuit for CLKLAHAQHSV2, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHAQHSV2 CK E ECK BC VDD VSS
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM39 pm cn nt11 VNW P12LL W=440.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=250.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=540.00n L=60.00n
MM45 s c nt21 VNW P12LL W=440.00n L=60.00n
MM54 nt21 pm VDD VNW P12LL W=540.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=540.00n L=60.00n
MM1 ten BC VDD VNW P12LL W=340.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=440.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=350.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=350.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=350.00n L=60.00n
MM51 s c VSS VPW N12LL W=350.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=430.00n L=60.00n
MM0 ten BC VSS VPW N12LL W=270.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=350.00n L=60.00n
.ENDS CLKLAHAQHSV2
****Sub-Circuit for CLKLAHAQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHAQHSV4 CK E ECK BC VDD VSS
MM51 s c VSS VPW N12LL W=300.00n L=60.00n
MM49 m pm VSS VPW N12LL W=300.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=300.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=260.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=300.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM0 ten BC VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=220.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=860.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=260.00n L=60.00n
MM45 s c nt21 VNW P12LL W=600.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=600.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=600.00n L=60.00n
MM1 ten BC VDD VNW P12LL W=300.00n L=60.00n
MM54 nt21 pm VDD VNW P12LL W=590.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=330.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.2u L=60.00n
MM39 pm cn nt11 VNW P12LL W=600.00n L=60.00n
.ENDS CLKLAHAQHSV4
****Sub-Circuit for CLKLAHAQHSV8, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHAQHSV8 CK E ECK BC VDD VSS
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM39 pm cn nt11 VNW P12LL W=540.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=250.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=1.3u L=60.00n
MM45 s c nt21 VNW P12LL W=1.08u L=60.00n
MM54 nt21 pm VDD VNW P12LL W=1.3u L=60.00n
MM21 ECK s VDD VNW P12LL W=2.16u L=60.00n
MM1 ten BC VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=540.00n L=60.00n
MM51 s c VSS VPW N12LL W=860.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=430.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=860.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=860.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=1.72u L=60.00n
MM0 ten BC VSS VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=430.00n L=60.00n
.ENDS CLKLAHAQHSV8
****Sub-Circuit for CLKLAHQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHQHSV1 CK E ECK FC VDD VSS
MM51 hnet12 FC VSS VPW N12LL W=300.00n L=60.00n
MM49 m pm VSS VPW N12LL W=300.00n L=60.00n
MM43 s pm VSS VPW N12LL W=230.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=300.00n L=60.00n
MM44 s c VSS VPW N12LL W=230.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=270n L=60.00n
MM27 cn CK VSS VPW N12LL W=220n L=60.00n
MM22 ECK s VSS VPW N12LL W=340.00n L=60.00n
MM36 pm c hnet12 VPW N12LL W=300.00n L=60.00n
MM45 s c hnet31 VNW P12LL W=550.00n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=550.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=590.0n L=60.00n
MM54 hnet13 FC VDD VNW P12LL W=590.0n L=60.00n
MM14 hnet21 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400n L=60.00n
MM28 cn CK VDD VNW P12LL W=330n L=60.00n
MM21 ECK s VDD VNW P12LL W=440.00n L=60.00n
MM39 pm cn hnet11 VNW P12LL W=590.0n L=60.00n
.ENDS CLKLAHQHSV1
****Sub-Circuit for CLKLAHQHSV2, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHQHSV2 CK E ECK FC VDD VSS
MM22 ECK s VSS VPW N12LL W=430.00n L=60.00n
MM44 s c VSS VPW N12LL W=270.00n L=60.00n
MM43 s pm VSS VPW N12LL W=270.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM51 hnet12 FC VSS VPW N12LL W=350.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=350.00n L=60.00n
MM36 pm c hnet12 VPW N12LL W=350.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270n L=60.00n
MM30 c cn VSS VPW N12LL W=350n L=60.00n
MM21 ECK s VDD VNW P12LL W=540.00n L=60.00n
MM45 s c hnet31 VNW P12LL W=500.00n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=500.00n L=60.00n
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM14 hnet21 c pm VNW P12LL W=250.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=250.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=440.0n L=60.00n
MM39 pm cn hnet11 VNW P12LL W=440.0n L=60.00n
MM54 hnet13 FC VDD VNW P12LL W=440.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=340n L=60.00n
MM29 c cn VDD VNW P12LL W=440n L=60.00n
.ENDS CLKLAHQHSV2
****Sub-Circuit for CLKLAHQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHQHSV4 CK E ECK FC VDD VSS
MM51 hnet12 FC VSS VPW N12LL W=340.00n L=60.00n
MM49 m pm VSS VPW N12LL W=400.00n L=60.00n
MM43 s pm VSS VPW N12LL W=280.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=340.00n L=60.00n
MM44 s c VSS VPW N12LL W=280.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=270n L=60.00n
MM27 cn CK VSS VPW N12LL W=220n L=60.00n
MM22 ECK s VSS VPW N12LL W=860n L=60.00n
MM36 pm c hnet12 VPW N12LL W=340.00n L=60.00n
MM45 s c hnet31 VNW P12LL W=640.00n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=640.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=650.0n L=60.00n
MM54 hnet13 FC VDD VNW P12LL W=650.0n L=60.00n
MM14 hnet21 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400n L=60.00n
MM28 cn CK VDD VNW P12LL W=330n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.2u L=60.00n
MM39 pm cn hnet11 VNW P12LL W=650.0n L=60.00n
.ENDS CLKLAHQHSV4
****Sub-Circuit for CLKLAHQHSV8, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHQHSV8 CK E ECK FC VDD VSS
MM22 ECK s VSS VPW N12LL W=1.72u L=60.00n
MM44 s c VSS VPW N12LL W=580.00n L=60.00n
MM43 s pm VSS VPW N12LL W=580.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM51 hnet12 FC VSS VPW N12LL W=430.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=430.00n L=60.00n
MM36 pm c hnet12 VPW N12LL W=430.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270n L=60.00n
MM30 c cn VSS VPW N12LL W=430n L=60.00n
MM21 ECK s VDD VNW P12LL W=2.16u L=60.00n
MM45 s c hnet31 VNW P12LL W=1080n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=1080n L=60.00n
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM14 hnet21 c pm VNW P12LL W=250.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=250.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=540.00n L=60.00n
MM39 pm cn hnet11 VNW P12LL W=540.00n L=60.00n
MM54 hnet13 FC VDD VNW P12LL W=540.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340n L=60.00n
MM29 c cn VDD VNW P12LL W=540n L=60.00n
.ENDS CLKLAHQHSV8
****Sub-Circuit for CLKLANAQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANAQHSV1 CK E ECK BC VDD VSS
MM51 nt22 BC VSS VPW N12LL W=300.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c nt22 VPW N12LL W=300.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=260.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=300.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=290.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=260.00n L=60.00n
MM45 s m nt21 VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=400.00n L=60.00n
MM54 nt21 BC VDD VNW P12LL W=300.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=360.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=460.00n L=60.00n
MM39 pm c nt11 VNW P12LL W=400.00n L=60.00n
.ENDS CLKLANAQHSV1
****Sub-Circuit for CLKLANAQHSV2, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT CLKLANAQHSV2 CK E ECK BC VDD VSS
MM39 pm c nt11 VNW P12LL W=440.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=440.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=250.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM50 m pm VDD VNW P12LL W=350.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM29 c cn VDD VNW P12LL W=430.00n L=60.00n
MM54 nt21 BC VDD VNW P12LL W=350.00n L=60.00n
MM45 s m nt21 VNW P12LL W=350.00n L=60.00n
MM46 s c VDD VNW P12LL W=350.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=540.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=350.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=350.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM49 m pm VSS VPW N12LL W=280.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=350.00n L=60.00n
MM51 nt22 BC VSS VPW N12LL W=350.00n L=60.00n
MM43 s c nt22 VPW N12LL W=350.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=430.00n L=60.00n
.ENDS CLKLANAQHSV2
****Sub-Circuit for CLKLANAQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANAQHSV4 CK E ECK BC VDD VSS
MM51 nt22 BC VSS VPW N12LL W=430.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c nt22 VPW N12LL W=430.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=320.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=270.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=800.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=320.00n L=60.00n
MM45 s m nt21 VNW P12LL W=430.00n L=60.00n
MM46 s c VDD VNW P12LL W=430.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=450.00n L=60.00n
MM54 nt21 BC VDD VNW P12LL W=430.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=360.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.3u L=60.00n
MM39 pm c nt11 VNW P12LL W=450.00n L=60.00n
.ENDS CLKLANAQHSV4
****Sub-Circuit for CLKLANAQHSV8, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT CLKLANAQHSV8 CK E ECK BC VDD VSS
MM21 ECK s VDD VNW P12LL W=2.16u L=60.00n
MM46 s c VDD VNW P12LL W=860.00n L=60.00n
MM45 s m nt21 VNW P12LL W=860.00n L=60.00n
MM54 nt21 BC VDD VNW P12LL W=860.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM50 m pm VDD VNW P12LL W=540.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=250.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=540.00n L=60.00n
MM39 pm c nt11 VNW P12LL W=540.00n L=60.00n
MM43 s c nt22 VPW N12LL W=860.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=1.72u L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM51 nt22 BC VSS VPW N12LL W=860.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=860.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM49 m pm VSS VPW N12LL W=430.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=430.00n L=60.00n
.ENDS CLKLANAQHSV8
****Sub-Circuit for CLKLANQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV1 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK s VSS VPW N12LL W=290.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK s VDD VNW P12LL W=460.00n L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV1
****Sub-Circuit for CLKLANQHSV12, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV12 CK E ECK FC VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=860.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK pq VSS VPW N12LL W=2.46u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.2u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK pq VDD VNW P12LL W=3.9u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV12
****Sub-Circuit for CLKLANQHSV16, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV16 CK E ECK FC VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=860.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK pq VSS VPW N12LL W=3.42u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.2u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK pq VDD VNW P12LL W=5.2u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV16
****Sub-Circuit for CLKLANQHSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV2 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK s VSS VPW N12LL W=420.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK s VDD VNW P12LL W=650.00n L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV2
****Sub-Circuit for CLKLANQHSV20, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV20 CK E ECK FC VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=1.29u L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK pq VSS VPW N12LL W=4.2u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.74u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK pq VDD VNW P12LL W=6.5u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV20
****Sub-Circuit for CLKLANQHSV24, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV24 CK E ECK FC VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=1.29u L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK pq VSS VPW N12LL W=5.16u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.74u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK pq VDD VNW P12LL W=7.8u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV24
****Sub-Circuit for CLKLANQHSV3, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV3 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=360.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=360.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK s VSS VPW N12LL W=620.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=400.00n L=60.00n
MM46 s c VDD VNW P12LL W=400.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK s VDD VNW P12LL W=960.00n L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV3
****Sub-Circuit for CLKLANQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV4 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=430.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=260n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK s VSS VPW N12LL W=800.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=500.00n L=60.00n
MM46 s c VDD VNW P12LL W=500.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.3u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV4
****Sub-Circuit for CLKLANQHSV6, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV6 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=340.00n L=60.00n
MM49 m pm VSS VPW N12LL W=380.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=430.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=340.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=360n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM22 ECK s VSS VPW N12LL W=1.14u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=340.00n L=60.00n
MM45 s m VDD VNW P12LL W=440.00n L=60.00n
MM46 s c VDD VNW P12LL W=440.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=600.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=600.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540n L=60.00n
MM28 cn CK VDD VNW P12LL W=450n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.95u L=60.00n
MM39 pm c hnet24 VNW P12LL W=600.0n L=60.00n
.ENDS CLKLANQHSV6
****Sub-Circuit for CLKLANQHSV8, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV8 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=360.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=740.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=740.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=360n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM22 ECK s VSS VPW N12LL W=1.6u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=800.0n L=60.00n
MM46 s c VDD VNW P12LL W=800.0n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540n L=60.00n
MM28 cn CK VDD VNW P12LL W=450n L=60.00n
MM21 ECK s VDD VNW P12LL W=2.6u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV8

****Sub-Circuit for LAHHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHHSV1 D G Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 c pm VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=400.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHHSV1
****Sub-Circuit for LAHHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHHSV2 D G Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 c pm VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=570.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=570.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LAHHSV2
****Sub-Circuit for LAHHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHHSV4 D G Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 c pm VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=650.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LAHHSV4
****Sub-Circuit for LAHRNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRNHSV1 D G Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=340.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=340.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=600.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=560.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=560.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHRNHSV1
****Sub-Circuit for LAHRNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRNHSV2 D G Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=410.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=390.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=410.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=560.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=560.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHRNHSV2
****Sub-Circuit for LAHRNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRNHSV4 D G Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net117 cn pm VNW P12LL W=350.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=350.00n L=60.00n
MM10 pm c net128 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LAHRNHSV4
****Sub-Circuit for LAHRSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRSNHSV1 D G Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=330.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=330.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=330.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHRSNHSV1
****Sub-Circuit for LAHRSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRSNHSV2 D G Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LAHRSNHSV2
****Sub-Circuit for LAHRSNHSV4, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT LAHRSNHSV4 D G Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM51 pm s VSS VPW N12LL W=240.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=360.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=650.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=640.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=640.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=510.00n L=60.00n
.ENDS LAHRSNHSV4
****Sub-Circuit for LAHSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHSNHSV1 D G Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=290.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 c net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=430.00n L=60.00n
MM47 Q net0127 VDD VNW P12LL W=430.00n L=60.00n
MM14 net0285 cn net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 c net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHSNHSV1
****Sub-Circuit for LAHSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHSNHSV2 D G Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=430.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 c net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 cn net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q net0127 VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 cn net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 c net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=440.00n L=60.00n
.ENDS LAHSNHSV2
****Sub-Circuit for LAHSNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHSNHSV4 D G Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=860.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=405.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 c net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=320.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=650.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q net0127 VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 cn net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 c net0292 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=510.00n L=60.00n
.ENDS LAHSNHSV4
****Sub-Circuit for LALHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALHSV1 D GN Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=400.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALHSV1
****Sub-Circuit for LALHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALHSV2 D GN Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=570.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=570.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LALHSV2
****Sub-Circuit for LALHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALHSV4 D GN Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=650.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LALHSV4
****Sub-Circuit for LALRNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRNHSV1 D GN Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=230.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=230.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=230.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=200.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS LALRNHSV1
****Sub-Circuit for LALRNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRNHSV2 D GN Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=310.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=390.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=310.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net117 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net128 VNW P12LL W=560.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=560.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALRNHSV2
****Sub-Circuit for LALRNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRNHSV4 D GN Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=380.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net117 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net128 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LALRNHSV4
****Sub-Circuit for LALRSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRSNHSV1 D GN Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=330.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=330.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=330.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALRSNHSV1
****Sub-Circuit for LALRSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRSNHSV2 D GN Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM51 pm s VSS VPW N12LL W=200.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=550.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=250.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LALRSNHSV2
****Sub-Circuit for LALRSNHSV4, Mon May 30 19:34:53 CST 2011****
.SUBCKT LALRSNHSV4 D GN Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0145 VSS VPW N12LL W=860.00n L=60.00n
MM51 net0145 s VSS VPW N12LL W=200.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=360.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 cn net0145 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 net0145 c net69 VPW N12LL W=420.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=420.00n L=60.00n
MM0 net_0154 net0145 VSS VPW N12LL W=360.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM52 net0145 s net0252 VNW P12LL W=290.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=290.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=640.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q net0145 VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 c net0145 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0145 cn net0292 VNW P12LL W=605.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=550.00n L=60.00n
MM1 net_0154 net0145 VDD VNW P12LL W=510.00n L=60.00n
.ENDS LALRSNHSV4
****Sub-Circuit for LALSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALSNHSV1 D GN Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALSNHSV1
****Sub-Circuit for LALSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALSNHSV2 D GN Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=430.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 cn net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 c net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q net0127 VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 c net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 cn net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=440.00n L=60.00n
.ENDS LALSNHSV2
****Sub-Circuit for LALSNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALSNHSV4 D GN Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=860.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 cn net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 c net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=320.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=650.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q net0127 VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 c net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 cn net0292 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=510.00n L=60.00n
.ENDS LALSNHSV4