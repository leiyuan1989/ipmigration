* SPICE INPUT		Tue Jan 14 09:25:35 2020	buftld4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld4
.subckt buftld4 OE A GND Y VDD
M1 GND N_5 Y GND mn5  l=0.5u w=0.72u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_5 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M7 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M8 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 N_2 N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld4
* SPICE INPUT		Tue Jan 14 09:25:40 2020	buftld6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld6
.subckt buftld6 A OE VDD GND Y
M1 N_4 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M8 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M11 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_6 N_4 N_3 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld6
* SPICE INPUT		Tue Jan 14 09:25:45 2020	buftld8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld8
.subckt buftld8 OE A Y VDD GND
M1 GND N_5 Y GND mn5  l=0.5u w=0.72u m=1
M2 GND N_5 Y GND mn5  l=0.5u w=0.72u m=1
M3 GND N_5 Y GND mn5  l=0.5u w=0.72u m=1
M4 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M6 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_5 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_5 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M10 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M11 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M12 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_6 N_2 N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld8
* SPICE INPUT		Wed Jul 10 13:23:44 2019	ad01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d0
.subckt ad01d0 GND S CO VDD B CI A
M1 N_4 N_15 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_3 CI N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_10 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_14 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_15 CI GND GND mn5  l=0.5u w=0.5u m=1
M11 CO N_14 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_10 N_9 N_3 GND mn5  l=0.5u w=0.5u m=1
M13 S N_2 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_10 N_3 GND mn5  l=0.5u w=0.5u m=1
M15 N_3 N_15 N_2 VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 CI N_2 VDD mp5  l=0.42u w=0.52u m=1
M17 N_10 A VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_3 N_7 N_10 VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_7 N_10 N_3 VDD mp5  l=0.42u w=0.52u m=1
M21 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_4 N_14 VDD mp5  l=0.42u w=0.52u m=1
M23 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 CI VDD VDD mp5  l=0.42u w=0.52u m=1
M25 CO N_14 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_4 N_9 N_10 VDD mp5  l=0.42u w=0.52u m=1
M27 S N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
.ends ad01d0
* SPICE INPUT		Wed Jul 10 13:23:52 2019	ad01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d1
.subckt ad01d1 VDD S CO GND A B CI
M1 N_4 N_15 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_3 CI N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_9 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_14 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_15 CI GND GND mn5  l=0.5u w=0.5u m=1
M11 CO N_14 GND GND mn5  l=0.5u w=0.58u m=1
M12 N_9 N_8 N_3 GND mn5  l=0.5u w=0.5u m=1
M13 S N_2 GND GND mn5  l=0.5u w=0.58u m=1
M14 N_8 N_9 N_3 GND mn5  l=0.5u w=0.5u m=1
M15 N_3 N_15 N_2 VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 CI N_2 VDD mp5  l=0.42u w=0.52u m=1
M17 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_3 N_7 N_9 VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_7 N_9 N_3 VDD mp5  l=0.42u w=0.52u m=1
M21 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_4 N_14 VDD mp5  l=0.42u w=0.52u m=1
M23 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 CI VDD VDD mp5  l=0.42u w=0.52u m=1
M25 CO N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 N_4 N_8 N_9 VDD mp5  l=0.42u w=0.52u m=1
M27 S N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M28 N_4 N_9 N_8 VDD mp5  l=0.42u w=0.52u m=1
.ends ad01d1
* SPICE INPUT		Wed Jul 10 13:23:59 2019	ad01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d2
.subckt ad01d2 VDD S CO GND A B CI
M1 N_4 N_15 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_3 CI N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_9 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_14 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_15 CI GND GND mn5  l=0.5u w=0.5u m=1
M11 CO N_14 GND GND mn5  l=0.5u w=0.72u m=1
M12 N_9 N_8 N_3 GND mn5  l=0.5u w=0.5u m=1
M13 S N_2 GND GND mn5  l=0.5u w=0.72u m=1
M14 N_8 N_9 N_3 GND mn5  l=0.5u w=0.5u m=1
M15 N_3 N_15 N_2 VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 CI N_2 VDD mp5  l=0.42u w=0.52u m=1
M17 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_3 N_7 N_9 VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_7 N_9 N_3 VDD mp5  l=0.42u w=0.52u m=1
M21 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_4 N_14 VDD mp5  l=0.42u w=0.52u m=1
M23 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 CI VDD VDD mp5  l=0.42u w=0.52u m=1
M25 CO N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 N_4 N_8 N_9 VDD mp5  l=0.42u w=0.52u m=1
M27 S N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_4 N_9 N_8 VDD mp5  l=0.42u w=0.52u m=1
.ends ad01d2
* SPICE INPUT		Wed Jul 10 13:24:06 2019	ah01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d0
.subckt ah01d0 VDD CO S GND B A
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 S N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M3 GND A N_6 GND mn5  l=0.5u w=0.5u m=1
M4 CO N_8 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_21 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M7 S B N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_21 A N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 N_7 S VDD mp5  l=0.42u w=0.52u m=1
M11 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M12 CO N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M14 S B N_4 VDD mp5  l=0.42u w=0.52u m=1
M15 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_8 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ah01d0
* SPICE INPUT		Wed Jul 10 13:24:13 2019	ah01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d1
.subckt ah01d1 VDD CO S GND A B
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 S N_7 N_4 GND mn5  l=0.5u w=0.58u m=1
M3 GND A N_5 GND mn5  l=0.5u w=0.5u m=1
M4 S B N_5 GND mn5  l=0.5u w=0.58u m=1
M5 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_21 A N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_21 B GND GND mn5  l=0.5u w=0.5u m=1
M8 CO N_8 GND GND mn5  l=0.5u w=0.58u m=1
M9 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 S N_7 N_5 VDD mp5  l=0.42u w=0.76u m=1
M11 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M12 S B N_4 VDD mp5  l=0.42u w=0.76u m=1
M13 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_8 A VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M16 CO N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends ah01d1
* SPICE INPUT		Wed Jul 10 13:24:20 2019	ah01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d2
.subckt ah01d2 VDD CO S GND B A
M1 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M2 S N_4 N_5 GND mn5  l=0.5u w=0.72u m=1
M3 N_6 B S GND mn5  l=0.5u w=0.72u m=1
M4 N_6 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 A N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_12 B GND GND mn5  l=0.5u w=0.5u m=1
M7 CO N_8 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_5 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 S N_4 N_6 VDD mp5  l=0.42u w=0.96u m=1
M11 N_8 A VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M14 CO N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_5 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 S B N_5 VDD mp5  l=0.42u w=0.96u m=1
.ends ah01d2
* SPICE INPUT		Wed Jul 10 13:24:28 2019	an02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d0
.subckt an02d0 B A VDD Y GND
M1 N_8 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an02d0
* SPICE INPUT		Wed Jul 10 13:24:35 2019	an02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d1
.subckt an02d1 B A VDD Y GND
M1 N_8 A N_2 GND mn5  l=0.5u w=0.58u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.58u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an02d1
* SPICE INPUT		Wed Jul 10 13:24:42 2019	an02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d2
.subckt an02d2 B A VDD Y GND
M1 N_8 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends an02d2
* SPICE INPUT		Wed Jul 10 13:24:49 2019	an03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d0
.subckt an03d0 C B A GND Y VDD
M1 N_9 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 C VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an03d0
* SPICE INPUT		Wed Jul 10 13:24:56 2019	an03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d1
.subckt an03d1 C B A Y GND VDD
M1 N_9 A N_2 GND mn5  l=0.5u w=0.58u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.58u m=1
M3 N_10 C GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 C VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an03d1
* SPICE INPUT		Wed Jul 10 13:25:04 2019	an03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d2
.subckt an03d2 C B A Y GND VDD
M1 N_9 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 C VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends an03d2
* SPICE INPUT		Wed Jul 10 13:25:11 2019	an04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d0
.subckt an04d0 GND Y VDD D C B A
M1 N_6 A N_4 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.58u m=1
M3 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 D GND GND mn5  l=0.5u w=0.58u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 C VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 D VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an04d0
* SPICE INPUT		Wed Jul 10 13:25:18 2019	an04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d1
.subckt an04d1 GND Y VDD D C B A
M1 N_6 A N_4 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.58u m=1
M3 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 D GND GND mn5  l=0.5u w=0.58u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 C VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 D VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an04d1
* SPICE INPUT		Wed Jul 10 13:25:25 2019	an04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d2
.subckt an04d2 GND Y VDD A B C D
M1 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.58u m=1
M3 N_6 A N_4 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 D GND GND mn5  l=0.5u w=0.58u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 C VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 D VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends an04d2
* SPICE INPUT		Wed Jul 10 13:25:33 2019	an12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an12d0
.subckt an12d0 B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_14 N_4 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_14 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an12d0
* SPICE INPUT		Wed Jul 10 13:25:40 2019	an12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an12d1
.subckt an12d1 B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_14 N_4 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_14 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an12d1
* SPICE INPUT		Wed Jul 10 13:25:47 2019	an12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an12d2
.subckt an12d2 B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 N_4 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends an12d2
* SPICE INPUT		Wed Jul 10 13:25:54 2019	an13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an13d0
.subckt an13d0 C B AN GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an13d0
* SPICE INPUT		Wed Jul 10 13:26:01 2019	an13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an13d1
.subckt an13d1 C B AN VDD GND Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an13d1
* SPICE INPUT		Wed Jul 10 13:26:08 2019	an13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an13d2
.subckt an13d2 C B AN VDD GND Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an13d2
* SPICE INPUT		Wed Jul 10 13:26:15 2019	an23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an23d0
.subckt an23d0 C BN AN VDD Y GND
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_3 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_12 C GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_5 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an23d0
* SPICE INPUT		Wed Jul 10 13:26:23 2019	an23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an23d1
.subckt an23d1 C BN AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_5 N_2 GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_2 C VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends an23d1
* SPICE INPUT		Wed Jul 10 13:26:30 2019	an23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an23d2
.subckt an23d2 C BN AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_3 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_12 C GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_6 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an23d2
* SPICE INPUT		Wed Jul 10 13:26:37 2019	antenna
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=antenna
.subckt antenna GND VDD A
D1 A VDD dppnw_5  area=0.63p pj=3.2u
D2 GND A dnppw_5  area=0.49p pj=2.8u
.ends antenna
* SPICE INPUT		Wed Jul 10 13:26:44 2019	aoi211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d0
.subckt aoi211d0 A0 A1 B0 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 Y A1 N_15 GND mn5  l=0.5u w=0.5u m=1
M4 N_15 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M6 N_6 B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M7 N_6 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi211d0
* SPICE INPUT		Wed Jul 10 13:26:51 2019	aoi211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d1
.subckt aoi211d1 A0 A1 B0 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.58u m=1
M2 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M3 Y A1 N_10 GND mn5  l=0.5u w=0.58u m=1
M4 N_10 A0 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y C0 N_16 VDD mp5  l=0.42u w=0.76u m=1
M6 N_6 B0 N_16 VDD mp5  l=0.42u w=0.76u m=1
M7 N_6 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_6 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aoi211d1
* SPICE INPUT		Wed Jul 10 13:26:58 2019	aoi211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d2
.subckt aoi211d2 A0 A1 B0 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A1 N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_10 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y C0 N_16 VDD mp5  l=0.42u w=0.96u m=1
M6 N_6 B0 N_16 VDD mp5  l=0.42u w=0.96u m=1
M7 N_6 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_6 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi211d2
* SPICE INPUT		Wed Jul 10 13:27:05 2019	aoi21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d0
.subckt aoi21d0 A0 A1 B0 GND Y VDD
M1 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_12 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y B0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M5 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi21d0
* SPICE INPUT		Wed Jul 10 13:27:13 2019	aoi21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d1
.subckt aoi21d1 A0 A1 B0 GND Y VDD
M1 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 A1 Y GND mn5  l=0.5u w=0.58u m=1
M3 N_9 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y B0 N_7 VDD mp5  l=0.42u w=0.76u m=1
M5 N_7 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 N_7 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aoi21d1
* SPICE INPUT		Wed Jul 10 13:27:20 2019	aoi21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d2
.subckt aoi21d2 A0 A1 B0 GND Y VDD
M1 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 A1 Y GND mn5  l=0.5u w=0.72u m=1
M3 N_9 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 N_7 VDD mp5  l=0.42u w=0.96u m=1
M5 N_7 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_7 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi21d2
* SPICE INPUT		Wed Jul 10 13:27:27 2019	aoi221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d0
.subckt aoi221d0 C0 A0 A1 B1 B0 VDD GND Y
M1 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B1 N_12 GND mn5  l=0.5u w=0.5u m=1
M3 N_13 A1 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_13 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y C0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_11 A1 N_7 VDD mp5  l=0.42u w=0.52u m=1
M10 N_11 A0 N_7 VDD mp5  l=0.42u w=0.52u m=1
.ends aoi221d0
* SPICE INPUT		Wed Jul 10 13:27:34 2019	aoi221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d1
.subckt aoi221d1 B0 A0 A1 B1 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.58u m=1
M2 Y B1 N_12 GND mn5  l=0.5u w=0.58u m=1
M3 N_13 A1 Y GND mn5  l=0.5u w=0.58u m=1
M4 N_13 A0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.58u m=1
M6 Y C0 N_8 VDD mp5  l=0.42u w=0.76u m=1
M7 N_7 B1 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_7 A1 N_8 VDD mp5  l=0.42u w=0.76u m=1
M9 N_7 A0 N_8 VDD mp5  l=0.42u w=0.76u m=1
M10 N_7 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aoi221d1
* SPICE INPUT		Wed Jul 10 13:27:41 2019	aoi221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d2
.subckt aoi221d2 B0 A0 A1 B1 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y B1 N_12 GND mn5  l=0.5u w=0.72u m=1
M3 N_13 A1 Y GND mn5  l=0.5u w=0.72u m=1
M4 N_13 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y C0 N_8 VDD mp5  l=0.42u w=0.96u m=1
M7 N_7 B1 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_7 A1 N_8 VDD mp5  l=0.42u w=0.96u m=1
M9 N_7 A0 N_8 VDD mp5  l=0.42u w=0.96u m=1
M10 N_7 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi221d2
* SPICE INPUT		Wed Jul 10 13:27:49 2019	aoi22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d0
.subckt aoi22d0 B0 B1 A1 A0 GND VDD Y
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 Y B1 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_8 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_8 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 B0 Y VDD mp5  l=0.42u w=0.52u m=1
.ends aoi22d0
* SPICE INPUT		Wed Jul 10 13:27:56 2019	aoi22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d1
.subckt aoi22d1 B0 B1 A1 A0 Y VDD GND
M1 N_11 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 Y A1 N_11 GND mn5  l=0.5u w=0.58u m=1
M3 Y B1 N_10 GND mn5  l=0.5u w=0.58u m=1
M4 N_10 B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_6 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 N_6 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_6 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M8 N_6 B0 Y VDD mp5  l=0.42u w=0.76u m=1
.ends aoi22d1
* SPICE INPUT		Wed Jul 10 13:28:03 2019	aoi22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d2
.subckt aoi22d2 A0 A1 B0 B1 GND Y VDD
M1 Y B1 N_10 GND mn5  l=0.5u w=0.72u m=1
M2 N_10 B0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A1 N_11 GND mn5  l=0.5u w=0.72u m=1
M4 N_11 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_8 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M6 N_8 B0 Y VDD mp5  l=0.42u w=0.96u m=1
M7 N_8 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_8 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi22d2
* SPICE INPUT		Wed Jul 10 13:28:11 2019	aoi31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d0
.subckt aoi31d0 A0 A1 A2 B0 VDD Y GND
M1 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A2 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_11 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M6 N_7 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi31d0
* SPICE INPUT		Wed Jul 10 13:28:18 2019	aoi31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d1
.subckt aoi31d1 B0 A2 A1 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_11 A1 N_10 GND mn5  l=0.5u w=0.58u m=1
M3 N_11 A2 Y GND mn5  l=0.5u w=0.58u m=1
M4 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_9 A2 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y B0 N_9 VDD mp5  l=0.42u w=0.76u m=1
.ends aoi31d1
* SPICE INPUT		Wed Jul 10 13:28:25 2019	aoi31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d2
.subckt aoi31d2 B0 A2 A1 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_11 A1 N_10 GND mn5  l=0.5u w=0.72u m=1
M3 N_11 A2 Y GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_9 A2 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y B0 N_9 VDD mp5  l=0.42u w=0.96u m=1
.ends aoi31d2
* SPICE INPUT		Wed Jul 10 13:28:32 2019	aoi32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d0
.subckt aoi32d0 GND Y VDD A1 A0 A2 B1 B0
M1 N_5 B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B1 N_5 GND mn5  l=0.5u w=0.5u m=1
M3 Y A2 N_7 GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A1 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_6 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_12 B0 Y VDD mp5  l=0.42u w=0.52u m=1
M7 N_12 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_12 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi32d0
* SPICE INPUT		Wed Jul 10 13:28:40 2019	aoi32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d1
.subckt aoi32d1 GND Y VDD B0 B1 A2 A1 A0
M1 N_6 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_7 A1 N_6 GND mn5  l=0.5u w=0.58u m=1
M3 Y A2 N_7 GND mn5  l=0.5u w=0.58u m=1
M4 Y B1 N_5 GND mn5  l=0.5u w=0.58u m=1
M5 N_5 B0 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_9 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_9 A2 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_9 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M10 N_9 B0 Y VDD mp5  l=0.42u w=0.76u m=1
.ends aoi32d1
* SPICE INPUT		Wed Jul 10 13:28:47 2019	aoi32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d2
.subckt aoi32d2 GND Y VDD A0 A1 A2 B1 B0
M1 N_5 B0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_6 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B1 N_5 GND mn5  l=0.5u w=0.72u m=1
M4 Y A2 N_7 GND mn5  l=0.5u w=0.72u m=1
M5 N_7 A1 N_6 GND mn5  l=0.5u w=0.72u m=1
M6 N_12 B0 Y VDD mp5  l=0.42u w=0.96u m=1
M7 N_12 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_12 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M9 N_12 A2 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_12 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi32d2
* SPICE INPUT		Wed Jul 10 13:28:54 2019	aoi33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d0
.subckt aoi33d0 GND Y VDD B0 B1 B2 A2 A1 A0
M1 N_6 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A1 N_6 GND mn5  l=0.5u w=0.5u m=1
M3 Y A2 N_7 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 B2 Y GND mn5  l=0.5u w=0.5u m=1
M5 N_8 B1 N_5 GND mn5  l=0.5u w=0.5u m=1
M6 N_5 B0 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y B2 N_10 VDD mp5  l=0.42u w=0.52u m=1
M11 Y B1 N_10 VDD mp5  l=0.42u w=0.52u m=1
M12 Y B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends aoi33d0
* SPICE INPUT		Wed Jul 10 13:29:01 2019	aoi33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d1
.subckt aoi33d1 GND Y VDD B0 B1 B2 A2 A1 A0
M1 N_6 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_7 A1 N_6 GND mn5  l=0.5u w=0.58u m=1
M3 Y A2 N_7 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 B2 Y GND mn5  l=0.5u w=0.58u m=1
M5 N_8 B1 N_5 GND mn5  l=0.5u w=0.58u m=1
M6 N_5 B0 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_11 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_11 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_11 A2 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y B2 N_11 VDD mp5  l=0.42u w=0.76u m=1
M11 Y B1 N_11 VDD mp5  l=0.42u w=0.76u m=1
M12 Y B0 N_11 VDD mp5  l=0.42u w=0.76u m=1
.ends aoi33d1
* SPICE INPUT		Wed Jul 10 13:29:08 2019	aoi33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d2
.subckt aoi33d2 GND Y VDD A0 A1 B1 A2 B2 B0
M1 N_8 B1 N_5 GND mn5  l=0.5u w=0.72u m=1
M2 N_6 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_8 B2 Y GND mn5  l=0.5u w=0.72u m=1
M4 Y A2 N_7 GND mn5  l=0.5u w=0.72u m=1
M5 N_5 B0 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_7 A1 N_6 GND mn5  l=0.5u w=0.72u m=1
M7 Y B1 N_14 VDD mp5  l=0.42u w=0.96u m=1
M8 N_14 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y B2 N_14 VDD mp5  l=0.42u w=0.96u m=1
M10 N_14 A2 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 Y B0 N_14 VDD mp5  l=0.42u w=0.96u m=1
M12 N_14 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aoi33d2
* SPICE INPUT		Wed Jul 10 13:29:15 2019	aoim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d0
.subckt aoim21d0 A1N A0N B0 GND VDD Y
M1 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 A0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1N GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 N_13 VDD mp5  l=0.42u w=0.52u m=1
M6 N_13 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_14 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A1N N_14 VDD mp5  l=0.42u w=0.52u m=1
.ends aoim21d0
* SPICE INPUT		Wed Jul 10 13:29:22 2019	aoim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d1
.subckt aoim21d1 B0 A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_14 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_13 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y B0 N_13 VDD mp5  l=0.42u w=0.76u m=1
.ends aoim21d1
* SPICE INPUT		Wed Jul 10 13:29:30 2019	aoim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d2
.subckt aoim21d2 B0 A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_14 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_13 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y B0 N_13 VDD mp5  l=0.42u w=0.96u m=1
.ends aoim21d2
* SPICE INPUT		Wed Jul 10 13:29:37 2019	aoim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d0
.subckt aoim22d0 B1 B0 A1N A0N GND VDD Y
M1 N_2 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_16 B0 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_16 B1 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 A1N N_11 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_10 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends aoim22d0
* SPICE INPUT		Wed Jul 10 13:29:45 2019	aoim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d1
.subckt aoim22d1 B0 B1 A1N A0N VDD Y GND
M1 N_2 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B1 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_11 B0 Y GND mn5  l=0.5u w=0.58u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_18 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 A1N N_18 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B1 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_10 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y N_2 N_10 VDD mp5  l=0.42u w=0.76u m=1
.ends aoim22d1
* SPICE INPUT		Wed Jul 10 13:29:52 2019	aoim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d2
.subckt aoim22d2 B0 B1 A1N A0N GND Y VDD
M1 N_2 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B1 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_11 B0 Y GND mn5  l=0.5u w=0.72u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_18 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 A1N N_18 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B1 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_10 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y N_2 N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends aoim22d2
* SPICE INPUT		Wed Jul 10 13:29:59 2019	aoim31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim31d0
.subckt aoim31d0 B0 A2N A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_12 A1N N_11 VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 A2N N_12 VDD mp5  l=0.42u w=0.52u m=1
M9 N_10 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends aoim31d0
* SPICE INPUT		Wed Jul 10 13:30:07 2019	aoim31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim31d1
.subckt aoim31d1 B0 A2N A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y B0 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_15 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_16 A1N N_15 VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 A2N N_16 VDD mp5  l=0.42u w=0.52u m=1
M9 N_14 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y B0 N_14 VDD mp5  l=0.42u w=0.76u m=1
.ends aoim31d1
* SPICE INPUT		Wed Jul 10 13:30:14 2019	aoim31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim31d2
.subckt aoim31d2 B0 A2N A1N A0N GND VDD Y
M1 N_3 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_15 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_16 A1N N_15 VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 A2N N_16 VDD mp5  l=0.42u w=0.52u m=1
M9 N_14 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y B0 N_14 VDD mp5  l=0.42u w=0.96u m=1
.ends aoim31d2
* SPICE INPUT		Wed Jul 10 13:30:21 2019	aor211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d0
.subckt aor211d0 C0 B0 A0 A1 GND Y VDD
M1 N_11 A1 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 C0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 C0 N_18 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor211d0
* SPICE INPUT		Wed Jul 10 13:30:29 2019	aor211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d1
.subckt aor211d1 C0 B0 A0 A1 VDD Y GND
M1 N_11 A1 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 C0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 C0 N_18 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aor211d1
* SPICE INPUT		Wed Jul 10 13:30:36 2019	aor211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d2
.subckt aor211d2 A1 A0 B0 C0 GND Y VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_6 C0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 A1 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_6 C0 N_18 VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 B0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor211d2
* SPICE INPUT		Wed Jul 10 13:30:43 2019	aor21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d0
.subckt aor21d0 B0 A1 A0 VDD Y GND
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor21d0
* SPICE INPUT		Wed Jul 10 13:30:50 2019	aor21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d1
.subckt aor21d1 B0 A1 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_3 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_3 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
.ends aor21d1
* SPICE INPUT		Wed Jul 10 13:30:58 2019	aor21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d2
.subckt aor21d2 B0 A1 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_3 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_3 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
.ends aor21d2
* SPICE INPUT		Wed Jul 10 13:31:05 2019	aor221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d0
.subckt aor221d0 GND Y VDD C0 A0 A1 B1 B0
M1 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B1 N_4 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_14 A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A0 N_14 VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_14 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_14 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor221d0
* SPICE INPUT		Wed Jul 10 13:31:12 2019	aor221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d1
.subckt aor221d1 GND Y VDD C0 A0 A1 B1 B0
M1 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_8 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B1 N_4 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_14 A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A0 N_14 VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M11 N_14 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_14 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor221d1
* SPICE INPUT		Wed Jul 10 13:31:19 2019	aor221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d2
.subckt aor221d2 GND Y VDD C0 A0 A1 B1 B0
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_8 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B1 N_4 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_14 A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A0 N_14 VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 N_14 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_14 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor221d2
* SPICE INPUT		Wed Jul 10 13:31:26 2019	aor22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d0
.subckt aor22d0 B0 B1 A1 A0 Y GND VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_12 B1 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B1 N_9 VDD mp5  l=0.42u w=0.52u m=1
M10 N_9 B0 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends aor22d0
* SPICE INPUT		Wed Jul 10 13:31:34 2019	aor22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d1
.subckt aor22d1 A0 A1 B1 B0 GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 B1 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_8 B0 N_6 VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B1 N_8 VDD mp5  l=0.42u w=0.52u m=1
M9 N_8 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_8 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor22d1
* SPICE INPUT		Wed Jul 10 13:31:41 2019	aor22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d2
.subckt aor22d2 A0 A1 B1 B0 Y VDD GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 B1 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_7 B0 N_6 VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B1 N_7 VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor22d2
* SPICE INPUT		Wed Jul 10 13:31:48 2019	aor311d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor311d0
.subckt aor311d0 GND Y VDD A2 A0 A1 B0 C0
M1 N_7 A1 N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A0 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_15 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor311d0
* SPICE INPUT		Wed Jul 10 13:31:55 2019	aor311d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor311d1
.subckt aor311d1 GND Y VDD A2 A0 A1 B0 C0
M1 N_7 A1 N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A0 N_7 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_15 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aor311d1
* SPICE INPUT		Wed Jul 10 13:32:02 2019	aor311d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor311d2
.subckt aor311d2 GND Y VDD A2 A0 A1 B0 C0
M1 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A1 N_4 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A0 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_15 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aor311d2
* SPICE INPUT		Wed Jul 10 13:32:10 2019	aor31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d0
.subckt aor31d0 B0 A2 A1 A0 Y VDD GND
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A2 N_12 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_9 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor31d0
* SPICE INPUT		Wed Jul 10 13:32:17 2019	aor31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d1
.subckt aor31d1 B0 A2 A1 A0 GND Y VDD
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A2 N_12 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends aor31d1
* SPICE INPUT		Wed Jul 10 13:32:24 2019	aor31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d2
.subckt aor31d2 B0 A2 A1 A0 GND Y VDD
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A2 N_12 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aor31d2
* SPICE INPUT		Wed Jul 10 13:32:31 2019	buffd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd0
.subckt buffd0 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends buffd0
* SPICE INPUT		Wed Jul 10 13:32:39 2019	buffd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd1
.subckt buffd1 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends buffd1
* SPICE INPUT		Wed Jul 10 13:32:46 2019	buffd10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd10
.subckt buffd10 GND Y VDD A
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M7 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 N_4 A VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_4 A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buffd10
* SPICE INPUT		Wed Jul 10 13:32:53 2019	buffd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd2
.subckt buffd2 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.58u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends buffd2
* SPICE INPUT		Wed Jul 10 13:33:00 2019	buffd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd3
.subckt buffd3 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.74u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.34u m=1
M3 N_4 A GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.72u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.72u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends buffd3
* SPICE INPUT		Wed Jul 10 13:33:08 2019	buffd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd4
.subckt buffd4 GND Y VDD A
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buffd4
* SPICE INPUT		Wed Jul 10 13:33:15 2019	buffd5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd5
.subckt buffd5 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.613u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.613u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.574u m=1
M4 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y N_4 VDD VDD mp5  l=0.42u w=0.48u m=1
M8 VDD A N_4 VDD mp5  l=0.42u w=0.96u m=1
.ends buffd5
* SPICE INPUT		Wed Jul 10 13:33:22 2019	buffd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd6
.subckt buffd6 GND Y VDD A
M1 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buffd6
* SPICE INPUT		Wed Jul 10 13:33:30 2019	buffd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd8
.subckt buffd8 GND Y VDD A
M1 N_4 A GND GND mn5  l=0.5u w=0.54u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.54u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_4 A VDD VDD mp5  l=0.42u w=0.72u m=1
M8 N_4 A VDD VDD mp5  l=0.42u w=0.72u m=1
M9 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buffd8
* SPICE INPUT		Wed Jul 10 13:33:37 2019	buftd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd0
.subckt buftd0 OE A GND Y VDD
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_3 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 OE GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_3 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 OE N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftd0
* SPICE INPUT		Wed Jul 10 13:33:44 2019	buftd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd1
.subckt buftd1 OE A GND Y VDD
M1 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_3 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 OE GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_3 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 OE N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftd1
* SPICE INPUT		Wed Jul 10 13:33:51 2019	buftd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd2
.subckt buftd2 A OE Y GND VDD
M1 N_4 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_6 OE N_2 VDD mp5  l=0.42u w=0.52u m=1
.ends buftd2
* SPICE INPUT		Wed Jul 10 13:33:59 2019	buftld0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld0
.subckt buftld0 A OE GND VDD Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 N_2 N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld0
* SPICE INPUT		Wed Jul 10 13:34:06 2019	buftld1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld1
.subckt buftld1 A OE GND VDD Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 N_2 N_5 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld1
* SPICE INPUT		Wed Jul 10 13:34:13 2019	buftld2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld2
.subckt buftld2 A OE VDD Y GND
M1 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 OE N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_5 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_6 N_5 N_2 VDD mp5  l=0.42u w=0.52u m=1
.ends buftld2
* SPICE INPUT		Wed Jul 10 13:34:20 2019	dfbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb1
.subckt dfbfb1 VDD QN Q GND RN SN CKN D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_26 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_6 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CKN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_6 N_28 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M18 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_6 N_5 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_4 N_5 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_4 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_6 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M38 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfbfb1
* SPICE INPUT		Wed Jul 10 13:34:27 2019	dfbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb2
.subckt dfbfb2 VDD QN Q GND RN SN CKN D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_26 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_6 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CKN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_6 N_28 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M20 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_6 N_5 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_4 N_5 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_4 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_6 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M40 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfbfb2
* SPICE INPUT		Wed Jul 10 13:34:34 2019	dfbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb1
.subckt dfbrb1 VDD QN Q GND RN SN CK D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_6 N_26 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CK GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_6 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_8 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M13 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M14 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M17 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_6 N_5 VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_6 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M34 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M37 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfbrb1
* SPICE INPUT		Wed Jul 10 13:34:42 2019	dfbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb2
.subckt dfbrb2 VDD QN Q GND RN SN CK D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_6 N_26 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CK GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_6 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_8 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M20 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_6 N_5 VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_6 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M40 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfbrb2
* SPICE INPUT		Wed Jul 10 13:34:49 2019	dfbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq1
.subckt dfbrq1 VDD Q GND RN D SN CK
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 SN GND GND mn5  l=0.5u w=0.58u m=1
M3 N_26 N_3 Q GND mn5  l=0.5u w=0.58u m=1
M4 N_26 N_8 Q GND mn5  l=0.5u w=0.58u m=1
M5 N_25 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_3 N_25 GND mn5  l=0.5u w=0.5u m=1
M7 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_5 N_30 GND mn5  l=0.5u w=0.5u m=1
M10 N_31 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M13 N_21 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_21 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_29 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M17 N_6 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M18 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M21 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M23 Q N_3 N_18 VDD mp5  l=0.42u w=0.76u m=1
M24 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_18 N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.5u m=1
M27 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M31 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M34 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M36 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M37 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M38 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfbrq1
* SPICE INPUT		Wed Jul 10 13:34:56 2019	dfbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq2
.subckt dfbrq2 VDD Q GND SN D RN CK
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_24 SN GND GND mn5  l=0.5u w=0.72u m=1
M6 N_24 N_3 Q GND mn5  l=0.5u w=0.72u m=1
M7 Q N_8 N_24 GND mn5  l=0.5u w=0.72u m=1
M8 N_23 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_3 N_23 GND mn5  l=0.5u w=0.5u m=1
M10 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M11 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_8 N_5 N_30 GND mn5  l=0.5u w=0.5u m=1
M13 N_31 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M14 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_19 SN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_19 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_19 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M18 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_29 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M20 N_6 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M21 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M26 Q N_3 N_18 VDD mp5  l=0.42u w=0.96u m=1
M27 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_18 N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.5u m=1
M30 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M34 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M40 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
.ends dfbrq2
* SPICE INPUT		Wed Jul 10 13:35:03 2019	dfcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb1
.subckt dfcfb1 GND QN Q VDD RN D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_14 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_15 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_8 N_4 N_16 GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M18 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M19 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_22 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M23 N_21 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M24 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M29 N_25 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M33 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M36 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfcfb1
* SPICE INPUT		Wed Jul 10 13:35:11 2019	dfcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb2
.subckt dfcfb2 GND QN Q VDD RN D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_14 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_15 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_8 N_4 N_16 GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M18 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M19 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_22 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M23 N_21 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M24 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M29 N_25 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M33 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M36 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfcfb2
* SPICE INPUT		Wed Jul 10 13:35:18 2019	dfcfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfq1
.subckt dfcfq1 GND Q VDD CKN D RN
M1 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_16 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_16 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_15 GND mn5  l=0.5u w=0.5u m=1
M9 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_14 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_13 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_25 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_24 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 N_24 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_25 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_23 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_22 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_22 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_21 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_20 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_20 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcfq1
* SPICE INPUT		Wed Jul 10 13:35:25 2019	dfcfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfq2
.subckt dfcfq2 GND Q VDD CKN D RN
M1 N_16 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_16 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 N_4 N_15 GND mn5  l=0.5u w=0.5u m=1
M5 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M7 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_14 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_13 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_35 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_35 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_34 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M21 N_36 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M22 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M24 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M25 N_34 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_33 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_33 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_32 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_31 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M30 N_32 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M31 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_36 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfcfq2
* SPICE INPUT		Wed Jul 10 13:35:32 2019	dfcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb1
.subckt dfcrb1 VDD QN Q GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_26 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_26 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M10 N_25 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_24 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_24 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_23 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_23 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M27 N_17 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_14 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M33 N_15 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M34 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrb1
* SPICE INPUT		Wed Jul 10 13:35:39 2019	dfcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb2
.subckt dfcrb2 GND QN Q VDD CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_17 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_5 N_16 GND mn5  l=0.5u w=0.5u m=1
M10 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_25 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M27 N_24 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_21 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M33 N_22 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M34 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrb2
* SPICE INPUT		Wed Jul 10 13:35:47 2019	dfcrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrn1
.subckt dfcrn1 VDD QN GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_34 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_34 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_33 GND mn5  l=0.5u w=0.5u m=1
M8 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_17 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrn1
* SPICE INPUT		Wed Jul 10 13:35:54 2019	dfcrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrn2
.subckt dfcrn2 VDD QN GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_23 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_22 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_22 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_21 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_21 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_17 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrn2
* SPICE INPUT		Wed Jul 10 13:36:01 2019	dfcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq1
.subckt dfcrq1 VDD Q GND CK D RN
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 Q N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_9 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_18 N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.52u m=1
M21 N_18 N_3 Q VDD mp5  l=0.42u w=0.76u m=1
M22 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrq1
* SPICE INPUT		Wed Jul 10 13:36:08 2019	dfcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq2
.subckt dfcrq2 VDD Q GND RN D CK
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_18 N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_18 N_3 Q VDD mp5  l=0.42u w=0.96u m=1
M21 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrq2
* SPICE INPUT		Wed Jul 10 13:36:15 2019	dfnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb1
.subckt dfnfb1 VDD QN Q GND D CKN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_5 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnfb1
* SPICE INPUT		Wed Jul 10 13:36:22 2019	dfnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb2
.subckt dfnfb2 VDD QN Q GND CKN D
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_5 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M15 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M18 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfnfb2
* SPICE INPUT		Wed Jul 10 13:36:30 2019	dfnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb1
.subckt dfnrb1 VDD QN Q GND CK D
M1 QN N_10 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_10 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_32 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_31 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_30 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M11 N_6 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_10 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_10 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 VDD N_10 N_16 VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M20 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M21 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M25 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M26 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfnrb1
* SPICE INPUT		Wed Jul 10 13:36:37 2019	dfnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb2
.subckt dfnrb2 VDD QN Q GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M17 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfnrb2
* SPICE INPUT		Wed Jul 10 13:36:44 2019	dfnrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrn1
.subckt dfnrn1 VDD QN GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrn1
* SPICE INPUT		Wed Jul 10 13:36:51 2019	dfnrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrn2
.subckt dfnrn2 VDD QN GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrn2
* SPICE INPUT		Wed Jul 10 13:36:58 2019	dfnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq1
.subckt dfnrq1 VDD Q GND CK D
M1 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrq1
* SPICE INPUT		Wed Jul 10 13:37:05 2019	dfnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq2
.subckt dfnrq2 VDD Q GND CK D
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrq2
* SPICE INPUT		Wed Jul 10 13:37:13 2019	dfpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb1
.subckt dfpfb1 VDD Q QN GND CKN D SN
M1 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_36 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_36 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_33 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_33 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfpfb1
* SPICE INPUT		Wed Jul 10 13:37:20 2019	dfpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb2
.subckt dfpfb2 VDD Q QN GND CKN D SN
M1 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_36 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_36 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M10 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_33 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M32 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M33 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfpfb2
* SPICE INPUT		Wed Jul 10 13:37:27 2019	dfprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb1
.subckt dfprb1 VDD Q QN GND SN D CK
M1 N_4 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_33 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_33 N_12 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_34 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_34 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_10 GND GND mn5  l=0.5u w=0.58u m=1
M7 QN N_8 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_10 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_35 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_35 SN N_6 GND mn5  l=0.5u w=0.5u m=1
M11 N_38 N_7 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_36 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_4 N_36 GND mn5  l=0.5u w=0.5u m=1
M14 N_37 N_12 N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_37 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_38 SN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_12 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_4 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_15 N_12 N_5 VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 Q N_10 VDD VDD mp5  l=0.42u w=0.76u m=1
M24 QN N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M25 N_10 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_6 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_6 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_12 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_17 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M32 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_8 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_12 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprb1
* SPICE INPUT		Wed Jul 10 13:37:34 2019	dfprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb2
.subckt dfprb2 VDD Q QN GND SN D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_34 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_34 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M10 N_35 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_4 N_35 GND mn5  l=0.5u w=0.5u m=1
M12 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M13 N_36 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M14 N_36 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_37 SN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_37 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_4 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_7 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_7 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M30 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M32 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfprb2
* SPICE INPUT		Wed Jul 10 13:37:41 2019	dfprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq1
.subckt dfprq1 VDD Q GND CK D SN
M1 Q N_8 N_27 GND mn5  l=0.5u w=0.58u m=1
M2 N_27 SN GND GND mn5  l=0.5u w=0.58u m=1
M3 N_33 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 N_33 GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_32 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_31 GND mn5  l=0.5u w=0.5u m=1
M8 N_31 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_30 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_30 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M19 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_9 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_14 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_7 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_7 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_11 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprq1
* SPICE INPUT		Wed Jul 10 13:37:48 2019	dfprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq2
.subckt dfprq2 VDD Q GND CK D SN
M1 Q N_10 N_29 GND mn5  l=0.5u w=0.72u m=1
M2 N_29 SN GND GND mn5  l=0.5u w=0.72u m=1
M3 N_35 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_34 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 N_10 N_35 GND mn5  l=0.5u w=0.5u m=1
M6 N_34 N_5 N_10 GND mn5  l=0.5u w=0.5u m=1
M7 N_10 N_4 N_33 GND mn5  l=0.5u w=0.5u m=1
M8 N_33 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_32 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_32 N_7 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M13 N_30 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_30 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_11 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_16 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_11 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_15 N_5 N_10 VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_9 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_13 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_5 N_7 VDD mp5  l=0.42u w=0.5u m=1
M29 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_4 N_10 VDD mp5  l=0.42u w=0.5u m=1
M31 VDD N_5 N_4 VDD mp5  l=0.42u w=0.5u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprq2
* SPICE INPUT		Wed Jul 10 13:37:55 2019	dl01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d0
.subckt dl01d0 A GND VDD Y
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dl01d0
* SPICE INPUT		Wed Jul 10 13:38:03 2019	dl01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d1
.subckt dl01d1 A GND VDD Y
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dl01d1
* SPICE INPUT		Wed Jul 10 13:38:10 2019	dl01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d2
.subckt dl01d2 A GND VDD Y
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dl01d2
* SPICE INPUT		Wed Jul 10 13:38:17 2019	dl02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d0
.subckt dl02d0 A Y VDD GND
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=1u w=0.5u m=1
M3 N_4 N_3 GND GND mn5  l=1u w=0.5u m=1
M4 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_5 N_4 VDD VDD mp5  l=0.84u w=0.52u m=1
M7 N_4 N_3 VDD VDD mp5  l=0.84u w=0.52u m=1
M8 N_3 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dl02d0
* SPICE INPUT		Wed Jul 10 13:38:24 2019	dl02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d1
.subckt dl02d1 A VDD Y GND
M1 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_4 GND GND mn5  l=1u w=0.5u m=1
M3 N_4 N_3 GND GND mn5  l=1u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_3 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.84u w=0.52u m=1
M7 N_4 N_3 VDD VDD mp5  l=0.84u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dl02d1
* SPICE INPUT		Wed Jul 10 13:38:32 2019	dl02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d2
.subckt dl02d2 A VDD Y GND
M1 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_4 GND GND mn5  l=1u w=0.5u m=1
M3 N_4 N_3 GND GND mn5  l=1u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_3 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.84u w=0.52u m=1
M7 N_4 N_3 VDD VDD mp5  l=0.84u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dl02d2
* SPICE INPUT		Wed Jul 10 14:07:11 2019	fillercap16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap16
.subckt fillercap16 VDD GND
M1 GND VDD GND GND mn5  l=6.582u w=0.72u m=1
M2 VDD GND VDD VDD mp5  l=6.582u w=0.96u m=1
.ends fillercap16
* SPICE INPUT		Wed Jul 10 14:07:18 2019	fillercap32
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap32
.subckt fillercap32 VDD GND
M1 GND VDD GND GND mn5  l=14.198u w=0.72u m=1
M2 VDD GND VDD VDD mp5  l=14.198u w=0.96u m=1
.ends fillercap32
* SPICE INPUT		Wed Jul 10 14:06:57 2019	fillercap4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap4
.subckt fillercap4 VDD GND
M1 GND VDD GND GND mn5  l=0.874u w=0.72u m=1
M2 VDD GND VDD VDD mp5  l=0.874u w=0.96u m=1
.ends fillercap4
* SPICE INPUT		Wed Jul 10 14:07:25 2019	fillercap64
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap64
.subckt fillercap64 VDD GND
M1 GND VDD GND GND mn5  l=29.43u w=0.72u m=1
M2 VDD GND VDD VDD mp5  l=29.43u w=0.96u m=1
.ends fillercap64
* SPICE INPUT		Wed Jul 10 14:07:04 2019	fillercap8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap8
.subckt fillercap8 VDD GND
M1 GND VDD GND GND mn5  l=2.774u w=0.72u m=1
M2 VDD GND VDD VDD mp5  l=2.774u w=0.96u m=1
.ends fillercap8
* SPICE INPUT		Wed Jul 10 13:38:39 2019	inv0d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d0
.subckt inv0d0 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.5u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends inv0d0
* SPICE INPUT		Wed Jul 10 13:38:46 2019	inv0d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d1
.subckt inv0d1 VDD Y GND A
M1 Y A GND GND mn5  l=0.5u w=0.58u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends inv0d1
* SPICE INPUT		Wed Jul 10 13:38:53 2019	inv0d10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d10
.subckt inv0d10 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A GND GND mn5  l=0.5u w=0.72u m=1
M5 Y A GND GND mn5  l=0.5u w=0.72u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d10
* SPICE INPUT		Wed Jul 10 13:39:00 2019	inv0d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d2
.subckt inv0d2 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d2
* SPICE INPUT		Wed Jul 10 13:39:08 2019	inv0d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d3
.subckt inv0d3 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.54u m=1
M2 Y A GND GND mn5  l=0.5u w=0.54u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.72u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.72u m=1
.ends inv0d3
* SPICE INPUT		Wed Jul 10 13:39:15 2019	inv0d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d4
.subckt inv0d4 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d4
* SPICE INPUT		Wed Jul 10 13:39:22 2019	inv0d5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d5
.subckt inv0d5 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.6u m=1
M2 Y A GND GND mn5  l=0.5u w=0.6u m=1
M3 Y A GND GND mn5  l=0.5u w=0.6u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.8u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.8u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.8u m=1
.ends inv0d5
* SPICE INPUT		Wed Jul 10 13:39:29 2019	inv0d6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d6
.subckt inv0d6 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d6
* SPICE INPUT		Wed Jul 10 13:39:36 2019	inv0d8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d8
.subckt inv0d8 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A GND GND mn5  l=0.5u w=0.72u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d8
* SPICE INPUT		Wed Jul 10 13:39:43 2019	invtd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtd0
.subckt invtd0 GND Y VDD OE A
M1 N_4 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_6 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y OE N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends invtd0
* SPICE INPUT		Wed Jul 10 13:39:51 2019	invtd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtd1
.subckt invtd1 A OE VDD GND Y
M1 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A GND GND mn5  l=0.5u w=0.58u m=1
M3 Y N_2 N_9 GND mn5  l=0.5u w=0.58u m=1
M4 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_14 A VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y OE N_14 VDD mp5  l=0.42u w=0.76u m=1
.ends invtd1
* SPICE INPUT		Wed Jul 10 13:39:58 2019	invtd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtd2
.subckt invtd2 A OE VDD GND Y
M1 N_2 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y N_2 N_9 GND mn5  l=0.5u w=0.72u m=1
M4 N_2 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_14 A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y OE N_14 VDD mp5  l=0.42u w=0.96u m=1
.ends invtd2
* SPICE INPUT		Wed Jul 10 13:40:05 2019	invtld0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld0
.subckt invtld0 GND Y VDD OE A
M1 N_4 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 Y OE N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_6 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 Y N_4 N_13 VDD mp5  l=0.42u w=0.52u m=1
M6 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends invtld0
* SPICE INPUT		Wed Jul 10 13:40:12 2019	invtld1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld1
.subckt invtld1 OE A GND VDD Y
M1 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A GND GND mn5  l=0.5u w=0.58u m=1
M3 Y OE N_9 GND mn5  l=0.5u w=0.58u m=1
M4 N_5 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_14 A VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y N_5 N_14 VDD mp5  l=0.42u w=0.76u m=1
.ends invtld1
* SPICE INPUT		Wed Jul 10 13:40:19 2019	invtld2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld2
.subckt invtld2 OE A GND VDD Y
M1 N_5 OE GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y OE N_9 GND mn5  l=0.5u w=0.72u m=1
M4 N_5 OE VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_14 A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y N_5 N_14 VDD mp5  l=0.42u w=0.96u m=1
.ends invtld2
* SPICE INPUT		Wed Jul 10 13:40:26 2019	labhb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=labhb1
.subckt labhb1 VDD QN Q GND RN D SN G
M1 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M4 N_22 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_22 RN N_21 GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_5 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 N_24 RN N_23 GND mn5  l=0.5u w=0.5u m=1
M10 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M11 Q N_7 GND GND mn5  l=0.5u w=0.58u m=1
M12 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_23 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_6 N_14 VDD mp5  l=0.42u w=0.52u m=1
M15 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_4 N_13 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_7 N_6 N_16 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 Q N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends labhb1
* SPICE INPUT		Wed Jul 10 13:40:34 2019	labhb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=labhb2
.subckt labhb2 VDD QN Q GND RN D SN G
M1 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M4 N_22 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_22 RN N_21 GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_5 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 N_24 RN N_23 GND mn5  l=0.5u w=0.5u m=1
M10 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M11 Q N_7 GND GND mn5  l=0.5u w=0.72u m=1
M12 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_23 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_6 N_14 VDD mp5  l=0.42u w=0.52u m=1
M15 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_4 N_13 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_7 N_6 N_16 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 Q N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends labhb2
* SPICE INPUT		Wed Jul 10 13:40:41 2019	lablb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb1
.subckt lablb1 VDD QN Q GND RN D SN GN
M1 N_6 SN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_22 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_22 RN N_21 GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_4 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 N_24 RN N_23 GND mn5  l=0.5u w=0.5u m=1
M10 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M11 Q N_7 GND GND mn5  l=0.5u w=0.58u m=1
M12 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_6 N_14 VDD mp5  l=0.42u w=0.52u m=1
M15 N_6 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_5 N_13 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_7 N_6 N_16 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 Q N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lablb1
* SPICE INPUT		Wed Jul 10 13:40:48 2019	lablb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb2
.subckt lablb2 VDD QN Q GND RN D SN GN
M1 N_6 SN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_22 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_22 RN N_21 GND mn5  l=0.5u w=0.5u m=1
M6 N_24 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_4 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 N_24 RN N_23 GND mn5  l=0.5u w=0.5u m=1
M10 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M11 Q N_7 GND GND mn5  l=0.5u w=0.72u m=1
M12 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M14 N_15 N_6 N_14 VDD mp5  l=0.42u w=0.52u m=1
M15 N_6 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_5 N_13 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_7 N_6 N_16 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 Q N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lablb2
* SPICE INPUT		Wed Jul 10 13:40:55 2019	lachb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb1
.subckt lachb1 RN D G GND QN Q VDD
M1 N_5 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_3 GND mn5  l=0.5u w=0.5u m=1
M6 N_21 RN N_20 GND mn5  l=0.5u w=0.5u m=1
M7 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_3 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_20 N_7 N_3 GND mn5  l=0.5u w=0.5u m=1
M11 N_21 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_7 G VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_3 N_7 N_31 VDD mp5  l=0.42u w=0.52u m=1
M16 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_32 N_5 N_3 VDD mp5  l=0.42u w=0.52u m=1
M18 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M19 Q N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_32 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lachb1
* SPICE INPUT		Wed Jul 10 13:41:02 2019	lachb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb2
.subckt lachb2 RN D G GND QN Q VDD
M1 N_5 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_3 GND mn5  l=0.5u w=0.5u m=1
M6 N_21 RN N_20 GND mn5  l=0.5u w=0.5u m=1
M7 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_3 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_20 N_7 N_3 GND mn5  l=0.5u w=0.5u m=1
M11 N_21 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_7 G VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_3 N_7 N_31 VDD mp5  l=0.42u w=0.52u m=1
M16 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_32 N_5 N_3 VDD mp5  l=0.42u w=0.52u m=1
M18 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 Q N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_32 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lachb2
* SPICE INPUT		Wed Jul 10 13:41:10 2019	lachq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachq1
.subckt lachq1 RN D G VDD GND Q
M1 N_3 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_6 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_16 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_17 RN N_16 GND mn5  l=0.5u w=0.5u m=1
M5 N_2 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_4 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_17 N_3 N_4 GND mn5  l=0.5u w=0.5u m=1
M8 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M9 N_18 N_6 N_4 GND mn5  l=0.5u w=0.5u m=1
M10 N_19 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_3 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 G VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 D VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_4 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M15 N_4 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M16 Q N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_29 N_3 N_4 VDD mp5  l=0.42u w=0.52u m=1
M19 N_29 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lachq1
* SPICE INPUT		Wed Jul 10 13:41:17 2019	lachq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachq2
.subckt lachq2 RN D G VDD GND Q
M1 N_3 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_6 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_16 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_17 RN N_16 GND mn5  l=0.5u w=0.5u m=1
M5 N_2 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_4 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_17 N_3 N_4 GND mn5  l=0.5u w=0.5u m=1
M8 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M9 N_18 N_6 N_4 GND mn5  l=0.5u w=0.5u m=1
M10 N_19 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_3 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_6 G VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 D VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_4 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M15 N_4 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M16 Q N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M17 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_29 N_3 N_4 VDD mp5  l=0.42u w=0.52u m=1
M19 N_29 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lachq2
* SPICE INPUT		Wed Jul 10 13:41:24 2019	laclb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb1
.subckt laclb1 RN D GN GND QN Q VDD
M1 N_7 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_3 GND mn5  l=0.5u w=0.5u m=1
M6 N_21 RN N_20 GND mn5  l=0.5u w=0.5u m=1
M7 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_3 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_20 N_7 N_3 GND mn5  l=0.5u w=0.5u m=1
M11 N_21 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_5 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_3 N_7 N_31 VDD mp5  l=0.42u w=0.52u m=1
M16 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_32 N_5 N_3 VDD mp5  l=0.42u w=0.52u m=1
M18 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M19 Q N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_32 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends laclb1
* SPICE INPUT		Wed Jul 10 13:41:31 2019	laclb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb2
.subckt laclb2 RN D GN GND QN Q VDD
M1 N_7 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_3 GND mn5  l=0.5u w=0.5u m=1
M6 N_21 RN N_20 GND mn5  l=0.5u w=0.5u m=1
M7 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_3 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_20 N_7 N_3 GND mn5  l=0.5u w=0.5u m=1
M11 N_21 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_5 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_3 N_7 N_31 VDD mp5  l=0.42u w=0.52u m=1
M16 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_32 N_5 N_3 VDD mp5  l=0.42u w=0.52u m=1
M18 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 Q N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_32 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends laclb2
* SPICE INPUT		Wed Jul 10 13:41:39 2019	laclq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclq1
.subckt laclq1 GN D RN VDD Q GND
M1 N_6 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_16 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 RN N_16 GND mn5  l=0.5u w=0.5u m=1
M7 N_19 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_2 GN GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_2 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_8 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M13 N_6 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_28 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_29 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_2 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_3 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_8 N_3 N_28 VDD mp5  l=0.42u w=0.52u m=1
M19 N_29 N_2 N_8 VDD mp5  l=0.42u w=0.52u m=1
.ends laclq1
* SPICE INPUT		Wed Jul 10 13:41:46 2019	laclq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclq2
.subckt laclq2 GN D RN VDD Q GND
M1 N_6 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_16 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 RN N_16 GND mn5  l=0.5u w=0.5u m=1
M7 N_19 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_2 GN GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_2 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_8 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 N_6 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_28 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_29 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_2 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_3 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_8 N_3 N_28 VDD mp5  l=0.42u w=0.52u m=1
M19 N_29 N_2 N_8 VDD mp5  l=0.42u w=0.52u m=1
.ends laclq2
* SPICE INPUT		Wed Jul 10 13:41:53 2019	lanhb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb1
.subckt lanhb1 D G GND QN Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_5 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_16 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_25 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_5 N_4 N_25 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 Q N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M18 N_26 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhb1
* SPICE INPUT		Wed Jul 10 13:42:00 2019	lanhb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb2
.subckt lanhb2 D G GND QN Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_5 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_16 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_25 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_5 N_4 N_25 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 Q N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M18 N_26 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhb2
* SPICE INPUT		Wed Jul 10 13:42:07 2019	lanhn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhn1
.subckt lanhn1 D G GND QN VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhn1
* SPICE INPUT		Wed Jul 10 13:42:14 2019	lanhn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhn2
.subckt lanhn2 D G GND QN VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhn2
* SPICE INPUT		Wed Jul 10 13:42:21 2019	lanhq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhq1
.subckt lanhq1 D G GND Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhq1
* SPICE INPUT		Wed Jul 10 13:42:29 2019	lanhq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhq2
.subckt lanhq2 D G GND Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhq2
* SPICE INPUT		Wed Jul 10 13:42:36 2019	lanht1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanht1
.subckt lanht1 GND Q VDD OE D G
M1 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 N_6 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_12 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_11 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q OE N_8 GND mn5  l=0.5u w=0.58u m=1
M10 N_3 OE GND GND mn5  l=0.5u w=0.5u m=1
M11 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_25 D VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 N_4 N_25 VDD mp5  l=0.42u w=0.52u m=1
M15 N_8 N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_26 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Q N_3 N_8 VDD mp5  l=0.42u w=0.76u m=1
M20 N_3 OE VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanht1
* SPICE INPUT		Wed Jul 10 13:42:43 2019	lanht2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanht2
.subckt lanht2 GND Q VDD OE D G
M1 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 N_6 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_12 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_11 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q OE N_8 GND mn5  l=0.5u w=0.72u m=1
M10 N_3 OE GND GND mn5  l=0.5u w=0.5u m=1
M11 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_25 D VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 N_4 N_25 VDD mp5  l=0.42u w=0.52u m=1
M15 N_8 N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_26 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Q N_3 N_8 VDD mp5  l=0.42u w=0.96u m=1
M20 N_3 OE VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanht2
* SPICE INPUT		Wed Jul 10 13:42:50 2019	lanlb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb1
.subckt lanlb1 GND QN Q VDD D GN
M1 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_7 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_6 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_11 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_10 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_6 N_5 N_22 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 Q N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_23 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_23 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlb1
* SPICE INPUT		Wed Jul 10 13:42:57 2019	lanlb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb2
.subckt lanlb2 GND QN Q VDD D GN
M1 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_7 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_6 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_11 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_10 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_6 N_5 N_22 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 Q N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_23 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_23 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlb2
* SPICE INPUT		Wed Jul 10 13:43:04 2019	lanln1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanln1
.subckt lanln1 D GN GND QN VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanln1
* SPICE INPUT		Wed Jul 10 13:43:11 2019	lanln2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanln2
.subckt lanln2 D GN GND QN VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanln2
* SPICE INPUT		Wed Jul 10 13:43:19 2019	lanlq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlq1
.subckt lanlq1 D GN GND Q VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlq1
* SPICE INPUT		Wed Jul 10 13:43:26 2019	lanlq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlq2
.subckt lanlq2 D GN GND Q VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlq2
* SPICE INPUT		Wed Jul 10 13:43:33 2019	laphb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb1
.subckt laphb1 GND QN Q VDD D SN G
M1 N_7 N_5 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M9 Q N_7 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 D VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_7 N_4 N_27 VDD mp5  l=0.42u w=0.52u m=1
M19 N_27 N_6 N_26 VDD mp5  l=0.42u w=0.52u m=1
M20 N_29 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends laphb1
* SPICE INPUT		Wed Jul 10 13:43:40 2019	laphb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb2
.subckt laphb2 GND QN Q VDD D SN G
M1 N_7 N_5 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M9 Q N_7 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 D VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_7 N_4 N_27 VDD mp5  l=0.42u w=0.52u m=1
M19 N_27 N_6 N_26 VDD mp5  l=0.42u w=0.52u m=1
M20 N_29 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M22 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends laphb2
* SPICE INPUT		Wed Jul 10 13:43:47 2019	laplb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb1
.subckt laplb1 GND QN Q VDD D SN GN
M1 N_7 N_4 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M9 Q N_7 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 D VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_7 N_5 N_27 VDD mp5  l=0.42u w=0.52u m=1
M19 N_27 N_6 N_26 VDD mp5  l=0.42u w=0.52u m=1
M20 N_29 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends laplb1
* SPICE INPUT		Wed Jul 10 13:43:55 2019	laplb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb2
.subckt laplb2 GND QN Q VDD D SN GN
M1 N_7 N_4 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 SN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M9 Q N_7 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_9 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_6 N_28 VDD mp5  l=0.42u w=0.52u m=1
M13 N_28 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 D VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_7 N_5 N_27 VDD mp5  l=0.42u w=0.52u m=1
M19 N_27 N_6 N_26 VDD mp5  l=0.42u w=0.52u m=1
M20 N_29 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M22 N_9 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends laplb2
* SPICE INPUT		Wed Jul 10 13:44:02 2019	mi02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d0
.subckt mi02d0 VDD Y GND S0 B A
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 N_3 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_5 S0 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y S0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mi02d0
* SPICE INPUT		Wed Jul 10 13:44:09 2019	mi02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d1
.subckt mi02d1 GND Y VDD A B S0
M1 N_5 B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 N_4 GND mn5  l=0.5u w=0.58u m=1
M3 Y S0 N_5 GND mn5  l=0.5u w=0.58u m=1
M4 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_3 N_5 VDD mp5  l=0.42u w=0.76u m=1
M7 N_5 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y S0 N_4 VDD mp5  l=0.42u w=0.76u m=1
M9 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mi02d1
* SPICE INPUT		Wed Jul 10 13:44:16 2019	mi02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d2
.subckt mi02d2 GND Y VDD S0 B A
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 N_4 GND mn5  l=0.5u w=0.72u m=1
M3 Y S0 N_5 GND mn5  l=0.5u w=0.72u m=1
M4 N_5 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y S0 N_4 VDD mp5  l=0.42u w=0.96u m=1
M8 Y N_3 N_5 VDD mp5  l=0.42u w=0.96u m=1
M9 N_5 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mi02d2
* SPICE INPUT		Wed Jul 10 13:44:23 2019	mi04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi04d0
.subckt mi04d0 VDD Y GND D C S0 B A S1
M1 N_11 N_13 N_15 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_7 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_10 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_7 S0 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_15 S1 N_12 GND mn5  l=0.5u w=0.5u m=1
M10 N_13 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M12 N_6 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 N_7 N_5 GND mn5  l=0.5u w=0.5u m=1
M14 N_5 C GND GND mn5  l=0.5u w=0.5u m=1
M15 Y N_15 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_15 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M17 N_12 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_11 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 S0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 S0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M23 N_10 N_7 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 S1 N_11 VDD mp5  l=0.42u w=0.52u m=1
M25 N_13 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 D VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 N_7 N_4 VDD mp5  l=0.42u w=0.52u m=1
M29 N_5 C VDD VDD mp5  l=0.42u w=0.52u m=1
M30 Y N_15 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mi04d0
* SPICE INPUT		Wed Jul 10 13:44:30 2019	mi04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi04d1
.subckt mi04d1 VDD Y GND C D S0 B A S1
M1 N_11 N_15 N_14 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_7 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M7 N_10 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_7 S0 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_14 S1 N_12 GND mn5  l=0.5u w=0.5u m=1
M10 N_15 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M12 N_6 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 N_7 N_5 GND mn5  l=0.5u w=0.5u m=1
M14 N_5 C GND GND mn5  l=0.5u w=0.5u m=1
M15 Y N_14 GND GND mn5  l=0.5u w=0.58u m=1
M16 N_14 N_15 N_12 VDD mp5  l=0.42u w=0.52u m=1
M17 N_12 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_11 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 S0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 S0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M23 N_10 N_7 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 S1 N_11 VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 D VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 N_7 N_4 VDD mp5  l=0.42u w=0.52u m=1
M29 N_5 C VDD VDD mp5  l=0.42u w=0.52u m=1
M30 Y N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends mi04d1
* SPICE INPUT		Wed Jul 10 13:44:37 2019	mi04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi04d2
.subckt mi04d2 GND Y VDD C D S0 B A S1
M1 N_11 N_13 N_14 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A GND GND mn5  l=0.5u w=0.5u m=1
M5 N_10 N_7 N_9 GND mn5  l=0.5u w=0.5u m=1
M6 N_6 S0 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_9 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_7 S0 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_14 S1 N_12 GND mn5  l=0.5u w=0.5u m=1
M10 N_13 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_6 N_7 N_4 GND mn5  l=0.5u w=0.5u m=1
M14 N_4 C GND GND mn5  l=0.5u w=0.5u m=1
M15 Y N_14 GND GND mn5  l=0.5u w=0.72u m=1
M16 N_14 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M17 N_12 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_10 A VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_4 S0 N_6 VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 S0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M23 N_9 N_7 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_14 S1 N_11 VDD mp5  l=0.42u w=0.52u m=1
M25 N_13 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_8 B VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 D VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_5 N_7 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_4 C VDD VDD mp5  l=0.42u w=0.52u m=1
M30 Y N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends mi04d2
* SPICE INPUT		Wed Jul 10 13:44:45 2019	mx02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d0
.subckt mx02d0 VDD Y GND S0 B A
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 S0 N_5 VDD mp5  l=0.42u w=0.52u m=1
M11 N_7 N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mx02d0
* SPICE INPUT		Wed Jul 10 13:44:52 2019	mx02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d1
.subckt mx02d1 GND Y VDD S0 B A
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 S0 N_5 VDD mp5  l=0.42u w=0.52u m=1
M11 N_7 N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mx02d1
* SPICE INPUT		Wed Jul 10 13:44:59 2019	mx02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d2
.subckt mx02d2 GND Y VDD S0 B A
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_7 B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 S0 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_7 B VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 S0 N_5 VDD mp5  l=0.42u w=0.52u m=1
M11 N_7 N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mx02d2
* SPICE INPUT		Wed Jul 10 13:45:06 2019	mx04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d0
.subckt mx04d0 GND Y VDD S1 A B S0 D C
M1 N_3 N_14 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 S1 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_8 D GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 B GND GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_10 N_3 GND mn5  l=0.5u w=0.5u m=1
M9 N_13 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_14 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_4 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_10 S0 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_3 S0 N_11 GND mn5  l=0.5u w=0.5u m=1
M14 N_4 N_14 N_2 VDD mp5  l=0.42u w=0.5u m=1
M15 N_2 S1 N_3 VDD mp5  l=0.42u w=0.5u m=1
M16 N_7 C VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_8 N_10 N_4 VDD mp5  l=0.42u w=0.5u m=1
M18 N_8 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_11 B VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_3 N_10 N_11 VDD mp5  l=0.42u w=0.5u m=1
M22 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_4 S0 N_7 VDD mp5  l=0.42u w=0.5u m=1
M25 N_10 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_3 S0 N_13 VDD mp5  l=0.42u w=0.5u m=1
.ends mx04d0
* SPICE INPUT		Wed Jul 10 13:45:13 2019	mx04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d1
.subckt mx04d1 GND Y VDD S1 A B S0 D C
M1 N_3 N_14 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 S1 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_8 D GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 B GND GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_10 N_3 GND mn5  l=0.5u w=0.5u m=1
M9 N_13 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_14 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_4 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_10 S0 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_3 S0 N_11 GND mn5  l=0.5u w=0.5u m=1
M14 N_4 N_14 N_2 VDD mp5  l=0.42u w=0.5u m=1
M15 N_2 S1 N_3 VDD mp5  l=0.42u w=0.5u m=1
M16 N_7 C VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_8 N_10 N_4 VDD mp5  l=0.42u w=0.5u m=1
M18 N_8 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_11 B VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_3 N_10 N_11 VDD mp5  l=0.42u w=0.5u m=1
M22 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_4 S0 N_7 VDD mp5  l=0.42u w=0.5u m=1
M25 N_10 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_3 S0 N_13 VDD mp5  l=0.42u w=0.5u m=1
.ends mx04d1
* SPICE INPUT		Wed Jul 10 13:45:20 2019	mx04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d2
.subckt mx04d2 GND Y VDD S1 A B S0 D C
M1 N_3 N_14 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 S1 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_8 D GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 B GND GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_10 N_3 GND mn5  l=0.5u w=0.5u m=1
M9 N_13 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_14 S1 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_4 S0 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_10 S0 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_3 S0 N_11 GND mn5  l=0.5u w=0.5u m=1
M14 N_4 N_14 N_2 VDD mp5  l=0.42u w=0.5u m=1
M15 N_2 S1 N_3 VDD mp5  l=0.42u w=0.5u m=1
M16 N_7 C VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_8 N_10 N_4 VDD mp5  l=0.42u w=0.5u m=1
M18 N_8 D VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_11 B VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_3 N_10 N_11 VDD mp5  l=0.42u w=0.5u m=1
M22 N_13 A VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 S1 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_4 S0 N_7 VDD mp5  l=0.42u w=0.5u m=1
M25 N_10 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_3 S0 N_13 VDD mp5  l=0.42u w=0.5u m=1
.ends mx04d2
* SPICE INPUT		Wed Jul 10 13:45:27 2019	nd02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d0
.subckt nd02d0 VDD Y GND B A
M1 Y A N_8 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd02d0
* SPICE INPUT		Wed Jul 10 13:45:35 2019	nd02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d1
.subckt nd02d1 VDD Y GND B A
M1 Y A N_8 GND mn5  l=0.5u w=0.58u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.58u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.76u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd02d1
* SPICE INPUT		Wed Jul 10 13:45:42 2019	nd02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d2
.subckt nd02d2 GND Y VDD B A
M1 Y A N_5 GND mn5  l=0.5u w=0.72u m=1
M2 N_5 B GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd02d2
* SPICE INPUT		Wed Jul 10 13:45:49 2019	nd03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d0
.subckt nd03d0 C B A Y VDD GND
M1 Y A N_8 GND mn5  l=0.5u w=0.5u m=1
M2 N_9 B N_8 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 C GND GND mn5  l=0.5u w=0.5u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd03d0
* SPICE INPUT		Wed Jul 10 13:45:56 2019	nd03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d1
.subckt nd03d1 A B C VDD GND Y
M1 N_9 C GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 B N_8 GND mn5  l=0.5u w=0.58u m=1
M3 Y A N_8 GND mn5  l=0.5u w=0.58u m=1
M4 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M5 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd03d1
* SPICE INPUT		Wed Jul 10 13:46:03 2019	nd03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d2
.subckt nd03d2 C B A Y VDD GND
M1 Y A N_8 GND mn5  l=0.5u w=0.72u m=1
M2 N_9 B N_8 GND mn5  l=0.5u w=0.72u m=1
M3 N_9 C GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M5 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd03d2
* SPICE INPUT		Wed Jul 10 13:46:10 2019	nd04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d0
.subckt nd04d0 C B D A GND VDD Y
M1 Y A N_9 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B N_9 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 C N_10 GND mn5  l=0.5u w=0.5u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y D VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd04d0
* SPICE INPUT		Wed Jul 10 13:46:17 2019	nd04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d1
.subckt nd04d1 GND Y VDD A B C D
M1 N_6 D GND GND mn5  l=0.5u w=0.58u m=1
M2 N_7 C N_6 GND mn5  l=0.5u w=0.58u m=1
M3 N_7 B N_5 GND mn5  l=0.5u w=0.58u m=1
M4 Y A N_5 GND mn5  l=0.5u w=0.58u m=1
M5 Y D VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M7 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd04d1
* SPICE INPUT		Wed Jul 10 13:46:24 2019	nd04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d2
.subckt nd04d2 D C B A Y VDD GND
M1 Y A N_9 GND mn5  l=0.5u w=0.72u m=1
M2 N_11 B N_9 GND mn5  l=0.5u w=0.72u m=1
M3 N_11 C N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_10 D GND GND mn5  l=0.5u w=0.72u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y D VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd04d2
* SPICE INPUT		Wed Jul 10 13:46:32 2019	nd12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d0
.subckt nd12d0 B AN Y VDD GND
M1 Y N_4 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd12d0
* SPICE INPUT		Wed Jul 10 13:46:39 2019	nd12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d1
.subckt nd12d1 B AN Y VDD GND
M1 Y N_4 N_12 GND mn5  l=0.5u w=0.58u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 B GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd12d1
* SPICE INPUT		Wed Jul 10 13:46:46 2019	nd12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d2
.subckt nd12d2 B AN Y VDD GND
M1 Y N_4 N_8 GND mn5  l=0.5u w=0.72u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd12d2
* SPICE INPUT		Wed Jul 10 13:46:53 2019	nd13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d0
.subckt nd13d0 GND Y VDD B C AN
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 C GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd13d0
* SPICE INPUT		Wed Jul 10 13:47:00 2019	nd13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d1
.subckt nd13d1 C AN B Y VDD GND
M1 Y N_5 N_9 GND mn5  l=0.5u w=0.58u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.58u m=1
M3 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.58u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd13d1
* SPICE INPUT		Wed Jul 10 13:47:07 2019	nd13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d2
.subckt nd13d2 C AN B Y VDD GND
M1 Y N_5 N_9 GND mn5  l=0.5u w=0.72u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.72u m=1
M3 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd13d2
* SPICE INPUT		Wed Jul 10 13:47:15 2019	nd14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d0
.subckt nd14d0 GND Y VDD B C D AN
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 C N_7 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 B N_6 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y D VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd14d0
* SPICE INPUT		Wed Jul 10 13:47:22 2019	nd14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d1
.subckt nd14d1 GND Y VDD B C D AN
M1 N_8 B N_6 GND mn5  l=0.5u w=0.58u m=1
M2 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M3 N_7 D GND GND mn5  l=0.5u w=0.58u m=1
M4 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 N_6 GND mn5  l=0.5u w=0.58u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.76u m=1
M7 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y D VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nd14d1
* SPICE INPUT		Wed Jul 10 13:47:29 2019	nd14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d2
.subckt nd14d2 GND Y VDD B C D AN
M1 N_8 B N_6 GND mn5  l=0.5u w=0.72u m=1
M2 N_8 C N_7 GND mn5  l=0.5u w=0.72u m=1
M3 N_7 D GND GND mn5  l=0.5u w=0.72u m=1
M4 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 N_6 GND mn5  l=0.5u w=0.72u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y D VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd14d2
* SPICE INPUT		Wed Jul 10 13:47:36 2019	nd23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd23d0
.subckt nd23d0 AN C BN GND Y VDD
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd23d0
* SPICE INPUT		Wed Jul 10 13:47:44 2019	nd23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd23d1
.subckt nd23d1 AN C BN GND Y VDD
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 N_11 GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_4 N_10 GND mn5  l=0.5u w=0.58u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.58u m=1
M5 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M10 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd23d1
* SPICE INPUT		Wed Jul 10 13:47:51 2019	nd23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd23d2
.subckt nd23d2 AN C BN GND Y VDD
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 N_11 GND mn5  l=0.5u w=0.72u m=1
M3 N_11 N_4 N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.72u m=1
M5 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd23d2
* SPICE INPUT		Wed Jul 10 13:47:58 2019	nd24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d0
.subckt nd24d0 GND Y VDD D AN C BN
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 C N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
M11 Y D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd24d0
* SPICE INPUT		Wed Jul 10 13:48:05 2019	nd24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d1
.subckt nd24d1 GND Y VDD D AN C BN
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 N_9 GND mn5  l=0.5u w=0.58u m=1
M3 N_9 N_3 N_8 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M5 N_7 D GND GND mn5  l=0.5u w=0.58u m=1
M6 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y C VDD VDD mp5  l=0.42u w=0.76u m=1
M11 Y D VDD VDD mp5  l=0.42u w=0.76u m=1
M12 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd24d1
* SPICE INPUT		Wed Jul 10 13:48:12 2019	nd24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d2
.subckt nd24d2 GND Y VDD D AN C BN
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 N_9 GND mn5  l=0.5u w=0.72u m=1
M3 N_9 N_3 N_8 GND mn5  l=0.5u w=0.72u m=1
M4 N_8 C N_7 GND mn5  l=0.5u w=0.72u m=1
M5 N_7 D GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M11 Y D VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd24d2
* SPICE INPUT		Wed Jul 10 13:48:19 2019	nr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d0
.subckt nr02d0 GND Y VDD B A
M1 Y A GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A VDD VDD mp5  l=0.42u w=0.52u m=1
M4 Y B N_7 VDD mp5  l=0.42u w=0.52u m=1
.ends nr02d0
* SPICE INPUT		Wed Jul 10 13:48:26 2019	nr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d1
.subckt nr02d1 GND Y VDD B A
M1 Y A GND GND mn5  l=0.5u w=0.58u m=1
M2 Y B GND GND mn5  l=0.5u w=0.58u m=1
M3 N_7 A VDD VDD mp5  l=0.42u w=0.76u m=1
M4 Y B N_7 VDD mp5  l=0.42u w=0.76u m=1
.ends nr02d1
* SPICE INPUT		Wed Jul 10 13:48:34 2019	nr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d2
.subckt nr02d2 GND Y VDD B A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y B GND GND mn5  l=0.5u w=0.72u m=1
M3 N_7 A VDD VDD mp5  l=0.42u w=0.96u m=1
M4 Y B N_7 VDD mp5  l=0.42u w=0.96u m=1
.ends nr02d2
* SPICE INPUT		Wed Jul 10 13:48:41 2019	nr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d0
.subckt nr03d0 A B C Y VDD GND
M1 Y C GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y A GND GND mn5  l=0.5u w=0.5u m=1
M4 Y C N_8 VDD mp5  l=0.42u w=0.52u m=1
M5 N_9 B N_8 VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr03d0
* SPICE INPUT		Wed Jul 10 13:48:48 2019	nr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d1
.subckt nr03d1 A B C GND VDD Y
M1 Y C GND GND mn5  l=0.5u w=0.58u m=1
M2 Y B GND GND mn5  l=0.5u w=0.58u m=1
M3 Y A GND GND mn5  l=0.5u w=0.58u m=1
M4 Y C N_11 VDD mp5  l=0.42u w=0.76u m=1
M5 N_12 B N_11 VDD mp5  l=0.42u w=0.76u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nr03d1
* SPICE INPUT		Wed Jul 10 13:48:55 2019	nr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d2
.subckt nr03d2 A B C GND VDD Y
M1 Y C GND GND mn5  l=0.5u w=0.72u m=1
M2 Y B GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C N_11 VDD mp5  l=0.42u w=0.96u m=1
M5 N_12 B N_11 VDD mp5  l=0.42u w=0.96u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nr03d2
* SPICE INPUT		Wed Jul 10 13:49:02 2019	nr04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d0
.subckt nr04d0 A B C D Y VDD GND
M1 Y D GND GND mn5  l=0.5u w=0.5u m=1
M2 Y C GND GND mn5  l=0.5u w=0.5u m=1
M3 Y B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y D N_9 VDD mp5  l=0.42u w=0.52u m=1
M6 N_11 C N_9 VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 B N_10 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr04d0
* SPICE INPUT		Wed Jul 10 13:49:10 2019	nr04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d1
.subckt nr04d1 A B C D GND VDD Y
M1 Y D GND GND mn5  l=0.5u w=0.58u m=1
M2 Y C GND GND mn5  l=0.5u w=0.58u m=1
M3 Y B GND GND mn5  l=0.5u w=0.58u m=1
M4 Y A GND GND mn5  l=0.5u w=0.58u m=1
M5 Y D N_12 VDD mp5  l=0.42u w=0.76u m=1
M6 N_14 C N_12 VDD mp5  l=0.42u w=0.76u m=1
M7 N_14 B N_13 VDD mp5  l=0.42u w=0.76u m=1
M8 N_13 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nr04d1
* SPICE INPUT		Wed Jul 10 13:49:17 2019	nr04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d2
.subckt nr04d2 A B C D GND VDD Y
M1 Y D GND GND mn5  l=0.5u w=0.72u m=1
M2 Y C GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A GND GND mn5  l=0.5u w=0.72u m=1
M5 Y D N_12 VDD mp5  l=0.42u w=0.96u m=1
M6 N_14 C N_12 VDD mp5  l=0.42u w=0.96u m=1
M7 N_14 B N_13 VDD mp5  l=0.42u w=0.96u m=1
M8 N_13 A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nr04d2
* SPICE INPUT		Wed Jul 10 13:49:24 2019	nr12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d0
.subckt nr12d0 AN B Y VDD GND
M1 Y B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 Y B N_8 VDD mp5  l=0.42u w=0.52u m=1
M5 N_8 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr12d0
* SPICE INPUT		Wed Jul 10 13:49:31 2019	nr12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d1
.subckt nr12d1 B AN GND VDD Y
M1 N_2 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.58u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_2 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M5 Y B N_12 VDD mp5  l=0.42u w=0.76u m=1
M6 N_12 N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends nr12d1
* SPICE INPUT		Wed Jul 10 13:49:38 2019	nr12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d2
.subckt nr12d2 B AN GND VDD Y
M1 N_2 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.72u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_2 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M5 Y B N_12 VDD mp5  l=0.42u w=0.96u m=1
M6 N_12 N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nr12d2
* SPICE INPUT		Wed Jul 10 13:49:45 2019	nr13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d0
.subckt nr13d0 AN B C Y VDD GND
M1 Y C GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_3 AN GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C N_9 VDD mp5  l=0.42u w=0.52u m=1
M6 N_10 B N_9 VDD mp5  l=0.42u w=0.52u m=1
M7 N_10 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr13d0
* SPICE INPUT		Wed Jul 10 13:49:53 2019	nr13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d1
.subckt nr13d1 C B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M3 Y B GND GND mn5  l=0.5u w=0.58u m=1
M4 Y C GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_10 N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_10 B N_9 VDD mp5  l=0.42u w=0.76u m=1
M8 Y C N_9 VDD mp5  l=0.42u w=0.76u m=1
.ends nr13d1
* SPICE INPUT		Wed Jul 10 13:50:00 2019	nr13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d2
.subckt nr13d2 C B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_14 B N_13 VDD mp5  l=0.42u w=0.96u m=1
M8 Y C N_13 VDD mp5  l=0.42u w=0.96u m=1
.ends nr13d2
* SPICE INPUT		Wed Jul 10 13:50:07 2019	nr14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d0
.subckt nr14d0 D C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 Y B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y C GND GND mn5  l=0.5u w=0.5u m=1
M5 Y D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_16 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M10 Y D N_14 VDD mp5  l=0.42u w=0.52u m=1
.ends nr14d0
* SPICE INPUT		Wed Jul 10 13:50:14 2019	nr14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d1
.subckt nr14d1 D C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M3 Y B GND GND mn5  l=0.5u w=0.58u m=1
M4 Y C GND GND mn5  l=0.5u w=0.58u m=1
M5 Y D GND GND mn5  l=0.5u w=0.58u m=1
M6 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_12 B N_11 VDD mp5  l=0.42u w=0.76u m=1
M9 N_12 C N_10 VDD mp5  l=0.42u w=0.76u m=1
M10 Y D N_10 VDD mp5  l=0.42u w=0.76u m=1
.ends nr14d1
* SPICE INPUT		Wed Jul 10 13:50:21 2019	nr14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d2
.subckt nr14d2 D C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C GND GND mn5  l=0.5u w=0.72u m=1
M5 Y D GND GND mn5  l=0.5u w=0.72u m=1
M6 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_12 B N_11 VDD mp5  l=0.42u w=0.96u m=1
M9 N_12 C N_10 VDD mp5  l=0.42u w=0.96u m=1
M10 Y D N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends nr14d2
* SPICE INPUT		Wed Jul 10 13:50:29 2019	nr23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr23d0
.subckt nr23d0 C AN BN GND VDD Y
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C GND GND mn5  l=0.5u w=0.5u m=1
M6 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_11 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M10 Y C N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends nr23d0
* SPICE INPUT		Wed Jul 10 13:50:36 2019	nr23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr23d1
.subckt nr23d1 C AN BN GND VDD Y
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y C GND GND mn5  l=0.5u w=0.58u m=1
M6 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_11 N_3 N_10 VDD mp5  l=0.42u w=0.76u m=1
M10 Y C N_10 VDD mp5  l=0.42u w=0.76u m=1
.ends nr23d1
* SPICE INPUT		Wed Jul 10 13:50:43 2019	nr23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr23d2
.subckt nr23d2 C AN BN GND VDD Y
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y C GND GND mn5  l=0.5u w=0.72u m=1
M6 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_11 N_3 N_10 VDD mp5  l=0.42u w=0.96u m=1
M10 Y C N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends nr23d2
* SPICE INPUT		Wed Jul 10 13:50:50 2019	nr24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d0
.subckt nr24d0 D C AN BN Y VDD GND
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y D GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_13 N_4 N_12 VDD mp5  l=0.42u w=0.52u m=1
M11 N_13 C N_11 VDD mp5  l=0.42u w=0.52u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends nr24d0
* SPICE INPUT		Wed Jul 10 13:50:57 2019	nr24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d1
.subckt nr24d1 D C AN BN Y VDD GND
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y C GND GND mn5  l=0.5u w=0.58u m=1
M6 Y D GND GND mn5  l=0.5u w=0.58u m=1
M7 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 N_13 N_4 N_12 VDD mp5  l=0.42u w=0.76u m=1
M11 N_13 C N_11 VDD mp5  l=0.42u w=0.76u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=0.76u m=1
.ends nr24d1
* SPICE INPUT		Wed Jul 10 13:51:04 2019	nr24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d2
.subckt nr24d2 D C AN BN Y VDD GND
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y C GND GND mn5  l=0.5u w=0.72u m=1
M6 Y D GND GND mn5  l=0.5u w=0.72u m=1
M7 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_13 N_4 N_12 VDD mp5  l=0.42u w=0.96u m=1
M11 N_13 C N_11 VDD mp5  l=0.42u w=0.96u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=0.96u m=1
.ends nr24d2
* SPICE INPUT		Wed Jul 10 13:51:12 2019	oai211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d0
.subckt oai211d0 C0 B0 A1 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 B0 N_16 GND mn5  l=0.5u w=0.5u m=1
M4 Y C0 N_16 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y A1 N_10 VDD mp5  l=0.42u w=0.52u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai211d0
* SPICE INPUT		Wed Jul 10 13:51:19 2019	oai211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d1
.subckt oai211d1 C0 B0 A1 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 B0 N_16 GND mn5  l=0.5u w=0.58u m=1
M4 Y C0 N_16 GND mn5  l=0.5u w=0.58u m=1
M5 N_10 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 Y A1 N_10 VDD mp5  l=0.42u w=0.76u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oai211d1
* SPICE INPUT		Wed Jul 10 13:51:26 2019	oai211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d2
.subckt oai211d2 A0 C0 A1 B0 Y VDD GND
M1 N_9 B0 N_10 GND mn5  l=0.5u w=0.72u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y C0 N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_9 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y A1 N_16 VDD mp5  l=0.42u w=0.96u m=1
M7 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_16 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oai211d2
* SPICE INPUT		Wed Jul 10 13:51:33 2019	oai21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d0
.subckt oai21d0 A0 B0 A1 VDD Y GND
M1 N_5 A1 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B0 N_5 GND mn5  l=0.5u w=0.5u m=1
M3 N_5 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 A1 Y VDD mp5  l=0.42u w=0.52u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_12 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai21d0
* SPICE INPUT		Wed Jul 10 13:51:41 2019	oai21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d1
.subckt oai21d1 A0 A1 B0 Y VDD GND
M1 N_5 B0 Y GND mn5  l=0.5u w=0.58u m=1
M2 N_5 A1 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_5 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M5 N_9 A1 Y VDD mp5  l=0.42u w=0.76u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oai21d1
* SPICE INPUT		Wed Jul 10 13:51:48 2019	oai21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d2
.subckt oai21d2 A0 A1 B0 Y VDD GND
M1 N_5 B0 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_5 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_5 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M5 N_9 A1 Y VDD mp5  l=0.42u w=0.96u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oai21d2
* SPICE INPUT		Wed Jul 10 13:51:55 2019	oai221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d0
.subckt oai221d0 C0 B1 A1 A0 B0 Y VDD GND
M1 N_7 B0 N_8 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 B1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_7 GND mn5  l=0.5u w=0.5u m=1
M6 N_13 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_12 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M10 N_13 B1 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oai221d0
* SPICE INPUT		Wed Jul 10 13:52:02 2019	oai221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d1
.subckt oai221d1 C0 B1 A1 A0 B0 Y VDD GND
M1 N_7 B0 N_8 GND mn5  l=0.5u w=0.58u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_8 B1 N_7 GND mn5  l=0.5u w=0.58u m=1
M5 Y C0 N_7 GND mn5  l=0.5u w=0.58u m=1
M6 N_13 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_12 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y A1 N_12 VDD mp5  l=0.42u w=0.76u m=1
M10 N_13 B1 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai221d1
* SPICE INPUT		Wed Jul 10 13:52:10 2019	oai221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d2
.subckt oai221d2 C0 B1 B0 A1 A0 Y VDD GND
M1 N_7 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_7 B0 N_8 GND mn5  l=0.5u w=0.72u m=1
M4 N_7 B1 N_8 GND mn5  l=0.5u w=0.72u m=1
M5 Y C0 N_8 GND mn5  l=0.5u w=0.72u m=1
M6 N_12 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y A1 N_12 VDD mp5  l=0.42u w=0.96u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_13 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_13 B1 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai221d2
* SPICE INPUT		Wed Jul 10 13:52:17 2019	oai222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d0
.subckt oai222d0 B0 A0 A1 B1 C0 C1 Y VDD GND
M1 N_11 C1 Y GND mn5  l=0.5u w=0.5u m=1
M2 N_11 C0 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B1 N_8 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_8 B0 N_11 GND mn5  l=0.5u w=0.5u m=1
M7 N_20 C1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C0 N_20 VDD mp5  l=0.42u w=0.52u m=1
M9 Y B1 N_9 VDD mp5  l=0.42u w=0.52u m=1
M10 Y A1 N_21 VDD mp5  l=0.42u w=0.52u m=1
M11 N_21 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_9 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai222d0
* SPICE INPUT		Wed Jul 10 13:52:24 2019	oai222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d1
.subckt oai222d1 C1 C0 B1 A1 A0 B0 GND VDD Y
M1 N_13 B0 N_10 GND mn5  l=0.5u w=0.58u m=1
M2 N_13 A0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_13 A1 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_10 B1 N_13 GND mn5  l=0.5u w=0.58u m=1
M5 N_10 C0 Y GND mn5  l=0.5u w=0.58u m=1
M6 Y C1 N_10 GND mn5  l=0.5u w=0.58u m=1
M7 N_12 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_21 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y A1 N_21 VDD mp5  l=0.42u w=0.76u m=1
M10 Y B1 N_12 VDD mp5  l=0.42u w=0.76u m=1
M11 Y C0 N_20 VDD mp5  l=0.42u w=0.76u m=1
M12 N_20 C1 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oai222d1
* SPICE INPUT		Wed Jul 10 13:52:31 2019	oai222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d2
.subckt oai222d2 GND Y VDD B0 A0 C1 B1 C0 A1
M1 N_4 C0 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_6 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_6 B0 N_4 GND mn5  l=0.5u w=0.72u m=1
M4 N_6 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 B1 N_6 GND mn5  l=0.5u w=0.72u m=1
M6 N_4 C1 Y GND mn5  l=0.5u w=0.72u m=1
M7 Y A1 N_24 VDD mp5  l=0.42u w=0.96u m=1
M8 N_13 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_24 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y C0 N_25 VDD mp5  l=0.42u w=0.96u m=1
M11 Y B1 N_13 VDD mp5  l=0.42u w=0.96u m=1
M12 VDD C1 N_25 VDD mp5  l=0.42u w=0.96u m=1
.ends oai222d2
* SPICE INPUT		Wed Jul 10 13:52:39 2019	oai22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d0
.subckt oai22d0 A0 A1 B1 B0 GND VDD Y
M1 Y B0 N_7 GND mn5  l=0.5u w=0.5u m=1
M2 Y B1 N_7 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_11 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M7 Y A1 N_10 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai22d0
* SPICE INPUT		Wed Jul 10 13:52:46 2019	oai22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d1
.subckt oai22d1 A1 A0 B0 B1 VDD Y GND
M1 Y B1 N_7 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B0 Y GND mn5  l=0.5u w=0.58u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_7 A1 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_11 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M6 N_11 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_10 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y A1 N_10 VDD mp5  l=0.42u w=0.76u m=1
.ends oai22d1
* SPICE INPUT		Wed Jul 10 13:52:53 2019	oai22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d2
.subckt oai22d2 A1 A0 B0 B1 VDD Y GND
M1 Y B1 N_7 GND mn5  l=0.5u w=0.72u m=1
M2 N_7 B0 Y GND mn5  l=0.5u w=0.72u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_7 A1 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_11 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M6 N_11 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_10 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y A1 N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends oai22d2
* SPICE INPUT		Wed Jul 10 13:53:00 2019	oai311d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai311d0
.subckt oai311d0 VDD Y GND C0 B0 A0 A1 A2
M1 N_11 A2 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_20 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_20 GND mn5  l=0.5u w=0.5u m=1
M6 N_7 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M7 N_8 A1 N_7 VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 VDD C0 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oai311d0
* SPICE INPUT		Wed Jul 10 13:53:07 2019	oai311d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai311d1
.subckt oai311d1 C0 A2 A1 A0 B0 VDD Y GND
M1 N_9 B0 N_18 GND mn5  l=0.5u w=0.58u m=1
M2 N_9 A0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 A1 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_9 A2 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y C0 N_18 GND mn5  l=0.5u w=0.58u m=1
M6 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_12 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_12 A1 N_11 VDD mp5  l=0.42u w=0.76u m=1
M9 N_11 A2 Y VDD mp5  l=0.42u w=0.76u m=1
M10 VDD C0 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai311d1
* SPICE INPUT		Wed Jul 10 13:53:14 2019	oai311d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai311d2
.subckt oai311d2 A0 B0 C0 A1 A2 Y VDD GND
M1 N_10 A2 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_10 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y C0 N_11 GND mn5  l=0.5u w=0.72u m=1
M4 N_10 B0 N_11 GND mn5  l=0.5u w=0.72u m=1
M5 N_10 A0 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_17 A2 Y VDD mp5  l=0.42u w=0.96u m=1
M7 N_18 A1 N_17 VDD mp5  l=0.42u w=0.96u m=1
M8 VDD C0 Y VDD mp5  l=0.42u w=0.96u m=1
M9 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_18 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oai311d2
* SPICE INPUT		Wed Jul 10 13:53:21 2019	oai31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d0
.subckt oai31d0 A2 A0 A1 B0 Y VDD GND
M1 Y B0 N_7 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_11 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 A0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A2 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oai31d0
* SPICE INPUT		Wed Jul 10 13:53:29 2019	oai31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d1
.subckt oai31d1 A2 A0 A1 B0 Y VDD GND
M1 Y B0 N_7 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_7 A2 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M6 N_11 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_11 A0 N_10 VDD mp5  l=0.42u w=0.76u m=1
M8 N_10 A2 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai31d1
* SPICE INPUT		Wed Jul 10 13:53:36 2019	oai31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d2
.subckt oai31d2 A2 B0 A0 A1 GND VDD Y
M1 N_8 A1 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B0 N_8 GND mn5  l=0.5u w=0.72u m=1
M4 N_8 A2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_15 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_15 A0 N_14 VDD mp5  l=0.42u w=0.96u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_14 A2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai31d2
* SPICE INPUT		Wed Jul 10 13:53:43 2019	oai321d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai321d0
.subckt oai321d0 B1 B0 A0 A1 A2 C0 VDD Y GND
M1 Y C0 N_10 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A2 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_10 B1 N_11 GND mn5  l=0.5u w=0.5u m=1
M7 N_17 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_19 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_19 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M12 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai321d0
* SPICE INPUT		Wed Jul 10 13:53:50 2019	oai321d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai321d1
.subckt oai321d1 A2 A1 A0 B0 B1 C0 GND Y VDD
M1 Y C0 N_11 GND mn5  l=0.5u w=0.58u m=1
M2 N_11 B1 N_10 GND mn5  l=0.5u w=0.58u m=1
M3 N_10 B0 N_11 GND mn5  l=0.5u w=0.58u m=1
M4 N_10 A0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_10 A1 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_10 A2 GND GND mn5  l=0.5u w=0.58u m=1
M7 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_15 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M9 N_15 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 N_14 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M11 N_14 A1 N_13 VDD mp5  l=0.42u w=0.76u m=1
M12 N_13 A2 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai321d1
* SPICE INPUT		Wed Jul 10 13:53:57 2019	oai321d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai321d2
.subckt oai321d2 A2 B0 B1 A1 A0 C0 GND Y VDD
M1 Y C0 N_9 GND mn5  l=0.5u w=0.72u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_8 B1 N_9 GND mn5  l=0.5u w=0.72u m=1
M5 N_8 B0 N_9 GND mn5  l=0.5u w=0.72u m=1
M6 N_8 A2 GND GND mn5  l=0.5u w=0.72u m=1
M7 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_14 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_14 A1 N_13 VDD mp5  l=0.42u w=0.96u m=1
M10 N_15 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M11 N_15 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_13 A2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai321d2
* SPICE INPUT		Wed Jul 10 13:54:05 2019	oai322d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai322d0
.subckt oai322d0 VDD Y GND B0 A0 A1 A2 B1 C0 C1
M1 N_11 B0 N_13 GND mn5  l=0.5u w=0.5u m=1
M2 Y C1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 C0 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_13 B1 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_13 A2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_13 A1 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 A0 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_8 C1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y C0 N_8 VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M11 Y A2 N_9 VDD mp5  l=0.42u w=0.52u m=1
M12 N_10 A1 N_9 VDD mp5  l=0.42u w=0.52u m=1
M13 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_3 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai322d0
* SPICE INPUT		Wed Jul 10 13:54:13 2019	oai322d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai322d1
.subckt oai322d1 Y VDD GND B0 A0 A1 A2 B1 C0 C1
M1 N_14 B0 N_12 GND mn5  l=0.5u w=0.58u m=1
M2 Y C1 N_12 GND mn5  l=0.5u w=0.58u m=1
M3 N_12 C0 Y GND mn5  l=0.5u w=0.58u m=1
M4 N_14 B1 N_12 GND mn5  l=0.5u w=0.58u m=1
M5 N_14 A2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_14 A1 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_14 A0 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_9 C1 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_9 C0 Y VDD mp5  l=0.42u w=0.76u m=1
M10 N_3 B1 Y VDD mp5  l=0.42u w=0.76u m=1
M11 N_10 A2 Y VDD mp5  l=0.42u w=0.76u m=1
M12 N_11 A1 N_10 VDD mp5  l=0.42u w=0.76u m=1
M13 N_11 A0 VDD VDD mp5  l=0.42u w=0.76u m=1
M14 N_3 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oai322d1
* SPICE INPUT		Wed Jul 10 13:54:20 2019	oai322d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai322d2
.subckt oai322d2 GND Y VDD A1 C1 A0 A2 B0 B1 C0
M1 N_3 B0 N_2 GND mn5  l=0.5u w=0.72u m=1
M2 N_2 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y C1 N_3 GND mn5  l=0.5u w=0.72u m=1
M4 N_2 B1 N_3 GND mn5  l=0.5u w=0.72u m=1
M5 N_2 A2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_3 C0 Y GND mn5  l=0.5u w=0.72u m=1
M7 N_2 A1 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_26 C1 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_12 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M10 N_26 C0 Y VDD mp5  l=0.42u w=0.96u m=1
M11 N_12 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_28 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 N_27 A2 Y VDD mp5  l=0.42u w=0.96u m=1
M14 N_28 A1 N_27 VDD mp5  l=0.42u w=0.96u m=1
.ends oai322d2
* SPICE INPUT		Wed Jul 10 13:54:27 2019	oai32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d0
.subckt oai32d0 A0 B1 A1 A2 B0 Y VDD GND
M1 N_7 B0 Y GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A2 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 B1 Y GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_16 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_17 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y B1 N_15 VDD mp5  l=0.42u w=0.52u m=1
M10 N_17 A0 N_16 VDD mp5  l=0.42u w=0.52u m=1
.ends oai32d0
* SPICE INPUT		Wed Jul 10 13:54:34 2019	oai32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d1
.subckt oai32d1 A2 B1 B0 A0 A1 GND VDD Y
M1 N_9 A1 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 A0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 B0 Y GND mn5  l=0.5u w=0.58u m=1
M4 N_9 B1 Y GND mn5  l=0.5u w=0.58u m=1
M5 N_9 A2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_13 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_13 A0 N_12 VDD mp5  l=0.42u w=0.76u m=1
M8 N_11 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y B1 N_11 VDD mp5  l=0.42u w=0.76u m=1
M10 N_12 A2 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oai32d1
* SPICE INPUT		Wed Jul 10 13:54:41 2019	oai32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d2
.subckt oai32d2 A2 B1 B0 A0 A1 GND VDD Y
M1 N_9 A1 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 B0 Y GND mn5  l=0.5u w=0.72u m=1
M4 N_9 B1 Y GND mn5  l=0.5u w=0.72u m=1
M5 N_9 A2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_13 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_13 A0 N_12 VDD mp5  l=0.42u w=0.96u m=1
M8 N_11 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y B1 N_11 VDD mp5  l=0.42u w=0.96u m=1
M10 N_12 A2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai32d2
* SPICE INPUT		Wed Jul 10 13:54:49 2019	oai33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d0
.subckt oai33d0 VDD Y GND B2 B1 B0 A1 A0 A2
M1 Y B0 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B2 N_12 GND mn5  l=0.5u w=0.5u m=1
M6 Y B1 N_12 GND mn5  l=0.5u w=0.5u m=1
M7 N_9 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_8 A0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M10 N_7 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M11 Y B2 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_9 B1 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends oai33d0
* SPICE INPUT		Wed Jul 10 13:54:56 2019	oai33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d1
.subckt oai33d1 VDD Y GND B2 B1 B0 A1 A0 A2
M1 Y B0 N_12 GND mn5  l=0.5u w=0.58u m=1
M2 N_12 A1 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_12 A0 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_12 A2 GND GND mn5  l=0.5u w=0.58u m=1
M5 Y B2 N_12 GND mn5  l=0.5u w=0.58u m=1
M6 Y B1 N_12 GND mn5  l=0.5u w=0.58u m=1
M7 N_9 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_8 A1 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_8 A0 N_7 VDD mp5  l=0.42u w=0.76u m=1
M10 N_7 A2 Y VDD mp5  l=0.42u w=0.76u m=1
M11 Y B2 N_6 VDD mp5  l=0.42u w=0.76u m=1
M12 N_9 B1 N_6 VDD mp5  l=0.42u w=0.76u m=1
.ends oai33d1
* SPICE INPUT		Wed Jul 10 13:55:03 2019	oai33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d2
.subckt oai33d2 VDD Y GND B2 B1 B0 A1 A0 A2
M1 N_14 A2 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_14 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B1 N_14 GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 N_14 GND mn5  l=0.5u w=0.72u m=1
M5 N_14 A1 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y B2 N_14 GND mn5  l=0.5u w=0.72u m=1
M7 N_7 A2 Y VDD mp5  l=0.42u w=0.96u m=1
M8 N_8 A0 N_7 VDD mp5  l=0.42u w=0.96u m=1
M9 N_9 B1 N_6 VDD mp5  l=0.42u w=0.96u m=1
M10 N_9 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 N_8 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 Y B2 N_6 VDD mp5  l=0.42u w=0.96u m=1
.ends oai33d2
* SPICE INPUT		Wed Jul 10 13:55:10 2019	oaim211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim211d0
.subckt oaim211d0 B0 C0 A0N A1N GND VDD Y
M1 N_11 A1N N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y C0 N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim211d0
* SPICE INPUT		Wed Jul 10 13:55:17 2019	oaim211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim211d1
.subckt oaim211d1 GND Y VDD C0 B0 A0N A1N
M1 N_7 A1N N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A0N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 N_4 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_8 B0 N_6 GND mn5  l=0.5u w=0.58u m=1
M5 Y C0 N_6 GND mn5  l=0.5u w=0.58u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oaim211d1
* SPICE INPUT		Wed Jul 10 13:55:25 2019	oaim211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim211d2
.subckt oaim211d2 GND Y VDD B0 C0 A0N A1N
M1 N_7 A1N N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A0N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C0 N_6 GND mn5  l=0.5u w=0.72u m=1
M5 N_8 B0 N_6 GND mn5  l=0.5u w=0.72u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oaim211d2
* SPICE INPUT		Wed Jul 10 13:55:32 2019	oaim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d0
.subckt oaim21d0 B0 A1N A0N VDD GND Y
M1 N_10 A0N N_3 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 N_9 GND mn5  l=0.5u w=0.5u m=1
M4 N_9 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim21d0
* SPICE INPUT		Wed Jul 10 13:55:39 2019	oaim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d1
.subckt oaim21d1 B0 A1N A0N VDD GND Y
M1 N_10 A0N N_3 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 N_9 GND mn5  l=0.5u w=0.58u m=1
M4 N_9 B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_3 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oaim21d1
* SPICE INPUT		Wed Jul 10 13:55:46 2019	oaim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d2
.subckt oaim21d2 B0 A1N A0N VDD GND Y
M1 N_10 A0N N_3 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 N_9 GND mn5  l=0.5u w=0.72u m=1
M4 N_9 B0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_3 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oaim21d2
* SPICE INPUT		Wed Jul 10 13:55:53 2019	oaim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d0
.subckt oaim22d0 B1 B0 A0N A1N Y VDD GND
M1 N_11 A1N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A0N N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 N_4 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_7 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_7 B1 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_18 B1 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oaim22d0
* SPICE INPUT		Wed Jul 10 13:56:00 2019	oaim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d1
.subckt oaim22d1 B1 B0 A0N A1N Y VDD GND
M1 N_11 A1N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A0N N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 N_4 Y GND mn5  l=0.5u w=0.58u m=1
M4 N_7 B0 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_7 B1 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M9 N_18 B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M10 N_18 B1 Y VDD mp5  l=0.42u w=0.76u m=1
.ends oaim22d1
* SPICE INPUT		Wed Jul 10 13:56:08 2019	oaim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d2
.subckt oaim22d2 B1 B0 A0N A1N Y VDD GND
M1 N_11 A1N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A0N N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 N_4 Y GND mn5  l=0.5u w=0.72u m=1
M4 N_7 B0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_7 B1 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_18 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_18 B1 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oaim22d2
* SPICE INPUT		Wed Jul 10 13:56:15 2019	oaim2m11d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim2m11d0
.subckt oaim2m11d0 C0 A0N B0N A1N VDD GND Y
M1 N_11 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_12 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A0N N_12 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_11 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_7 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B0N N_7 VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim2m11d0
* SPICE INPUT		Wed Jul 10 13:56:22 2019	oaim2m11d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim2m11d1
.subckt oaim2m11d1 C0 A0N B0N A1N VDD GND Y
M1 N_11 N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_12 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A0N N_12 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_11 GND mn5  l=0.5u w=0.58u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_7 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B0N N_7 VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends oaim2m11d1
* SPICE INPUT		Wed Jul 10 13:56:30 2019	oaim2m11d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim2m11d2
.subckt oaim2m11d2 C0 B0N A1N A0N VDD Y GND
M1 N_3 A0N N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 B0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y C0 N_11 GND mn5  l=0.5u w=0.72u m=1
M6 N_9 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 B0N N_9 VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oaim2m11d2
* SPICE INPUT		Wed Jul 10 13:56:37 2019	oaim31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim31d0
.subckt oaim31d0 GND Y VDD A1N A2N B0 A0N
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1N N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0N N_4 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A2N VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim31d0
* SPICE INPUT		Wed Jul 10 13:56:44 2019	oaim31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim31d1
.subckt oaim31d1 GND Y VDD A1N A2N A0N B0
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.58u m=1
M2 N_6 B0 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_8 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1N N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0N N_4 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_4 A2N VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim31d1
* SPICE INPUT		Wed Jul 10 13:56:51 2019	oaim31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim31d2
.subckt oaim31d2 GND Y VDD A1N A2N B0 A0N
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.72u m=1
M2 N_6 B0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_8 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1N N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0N N_4 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_4 A2N VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim31d2
* SPICE INPUT		Wed Jul 10 13:56:58 2019	or02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d0
.subckt or02d0 A B VDD GND Y
M1 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 B N_3 VDD mp5  l=0.42u w=0.52u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or02d0
* SPICE INPUT		Wed Jul 10 13:57:05 2019	or02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d1
.subckt or02d1 A B VDD GND Y
M1 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_12 B N_2 VDD mp5  l=0.42u w=0.52u m=1
M5 N_12 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends or02d1
* SPICE INPUT		Wed Jul 10 13:57:12 2019	or02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d2
.subckt or02d2 A B GND VDD Y
M1 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 B N_3 VDD mp5  l=0.42u w=0.52u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or02d2
* SPICE INPUT		Wed Jul 10 13:57:20 2019	or03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d0
.subckt or03d0 B A C GND VDD Y
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_13 C N_3 VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_14 B N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends or03d0
* SPICE INPUT		Wed Jul 10 13:57:27 2019	or03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d1
.subckt or03d1 B A C GND VDD Y
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_13 C N_3 VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_14 B N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends or03d1
* SPICE INPUT		Wed Jul 10 13:57:34 2019	or03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d2
.subckt or03d2 B A C GND VDD Y
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_13 C N_3 VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_14 B N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends or03d2
* SPICE INPUT		Wed Jul 10 13:57:41 2019	or04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d0
.subckt or04d0 A B D C VDD Y GND
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_14 D N_3 VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_16 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or04d0
* SPICE INPUT		Wed Jul 10 13:57:48 2019	or04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d1
.subckt or04d1 D A C B VDD Y GND
M1 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 D GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_14 D N_2 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends or04d1
* SPICE INPUT		Wed Jul 10 13:57:55 2019	or04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d2
.subckt or04d2 D A B C VDD Y GND
M1 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 D GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_15 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_14 D N_2 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends or04d2
* SPICE INPUT		Wed Jul 10 13:58:03 2019	or12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or12d0
.subckt or12d0 B AN VDD GND Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_14 B N_2 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or12d0
* SPICE INPUT		Wed Jul 10 13:58:10 2019	or12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or12d1
.subckt or12d1 AN B Y VDD GND
M1 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_2 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_14 B N_4 VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_2 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_14 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or12d1
* SPICE INPUT		Wed Jul 10 13:58:17 2019	or12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or12d2
.subckt or12d2 AN B Y VDD GND
M1 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_14 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 B N_2 VDD mp5  l=0.42u w=0.52u m=1
M7 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends or12d2
* SPICE INPUT		Wed Jul 10 13:58:24 2019	or13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or13d0
.subckt or13d0 C B AN Y VDD GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_15 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C N_16 VDD mp5  l=0.42u w=0.52u m=1
.ends or13d0
* SPICE INPUT		Wed Jul 10 13:58:32 2019	or13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or13d1
.subckt or13d1 AN C B GND VDD Y
M1 N_5 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_5 B GND GND mn5  l=0.5u w=0.5u m=1
M4 N_5 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 C N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or13d1
* SPICE INPUT		Wed Jul 10 13:58:39 2019	or13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or13d2
.subckt or13d2 C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 C N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends or13d2
* SPICE INPUT		Wed Jul 10 13:58:46 2019	or23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or23d0
.subckt or23d0 AN C BN Y VDD GND
M1 N_6 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 BN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_3 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_18 N_7 N_17 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C N_18 VDD mp5  l=0.42u w=0.52u m=1
M11 N_17 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_3 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or23d0
* SPICE INPUT		Wed Jul 10 13:58:53 2019	or23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or23d1
.subckt or23d1 AN C BN Y VDD GND
M1 N_5 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_5 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_2 C N_18 VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 N_5 N_17 VDD mp5  l=0.42u w=0.52u m=1
M10 N_17 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends or23d1
* SPICE INPUT		Wed Jul 10 13:59:00 2019	or23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or23d2
.subckt or23d2 BN C AN Y VDD GND
M1 N_6 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 BN GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_6 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_17 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 N_5 N_17 VDD mp5  l=0.42u w=0.52u m=1
M10 N_2 C N_18 VDD mp5  l=0.42u w=0.52u m=1
M11 N_5 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends or23d2
* SPICE INPUT		Wed Jul 10 13:59:08 2019	ora211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d0
.subckt ora211d0 C0 B0 A1 A0 GND Y VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_6 C0 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_17 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora211d0
* SPICE INPUT		Wed Jul 10 13:59:15 2019	ora211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d1
.subckt ora211d1 A1 B0 C0 A0 GND VDD Y
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_5 C0 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A1 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_5 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
.ends ora211d1
* SPICE INPUT		Wed Jul 10 13:59:22 2019	ora211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d2
.subckt ora211d2 A1 B0 C0 A0 VDD Y GND
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_5 C0 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A1 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_5 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
.ends ora211d2
* SPICE INPUT		Wed Jul 10 13:59:30 2019	ora21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d0
.subckt ora21d0 B0 A1 A0 Y VDD GND
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_6 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B0 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_5 A1 N_14 VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora21d0
* SPICE INPUT		Wed Jul 10 13:59:37 2019	ora21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d1
.subckt ora21d1 B0 A1 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 N_9 GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_14 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 A1 N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends ora21d1
* SPICE INPUT		Wed Jul 10 13:59:44 2019	ora21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d2
.subckt ora21d2 A1 B0 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_4 B0 N_9 GND mn5  l=0.5u w=0.5u m=1
M4 N_9 A1 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_14 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_4 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A1 N_14 VDD mp5  l=0.42u w=0.52u m=1
.ends ora21d2
* SPICE INPUT		Wed Jul 10 13:59:51 2019	ora311d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora311d1
.subckt ora311d1 C0 B0 A2 A1 A0 Y VDD GND
M1 Y N_7 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 B0 N_12 GND mn5  l=0.5u w=0.5u m=1
M6 N_12 C0 N_7 GND mn5  l=0.5u w=0.5u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_19 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_19 A1 N_18 VDD mp5  l=0.42u w=0.52u m=1
M10 N_18 A2 N_7 VDD mp5  l=0.42u w=0.52u m=1
M11 N_7 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_7 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora311d1
* SPICE INPUT		Wed Jul 10 13:59:58 2019	ora311d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora311d2
.subckt ora311d2 A0 A1 A2 B0 C0 Y VDD GND
M1 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_12 C0 N_7 GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B0 N_12 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_7 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_18 A2 N_7 VDD mp5  l=0.42u w=0.52u m=1
M11 N_19 A1 N_18 VDD mp5  l=0.42u w=0.52u m=1
M12 N_19 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora311d2
* SPICE INPUT		Wed Jul 10 14:00:06 2019	ora31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d0
.subckt ora31d0 B0 A2 A0 A1 Y VDD GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 B0 N_7 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 A0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A2 N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora31d0
* SPICE INPUT		Wed Jul 10 14:00:13 2019	ora31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d1
.subckt ora31d1 A0 A2 B0 A1 GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_10 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_15 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A2 N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_16 A0 N_15 VDD mp5  l=0.42u w=0.52u m=1
.ends ora31d1
* SPICE INPUT		Wed Jul 10 14:00:20 2019	ora31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d2
.subckt ora31d2 A0 A2 B0 A1 GND VDD Y
M1 N_10 A1 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_5 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_5 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 A2 N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_16 A0 N_15 VDD mp5  l=0.42u w=0.52u m=1
.ends ora31d2
* SPICE INPUT		Wed Jul 10 14:00:28 2019	sdbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb1
.subckt sdbfb1 VDD Q QN GND RN SN SI SE D CKN
M1 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M9 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M10 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M11 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_9 N_5 N_29 GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_4 N_55 GND mn5  l=0.5u w=0.5u m=1
M14 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M16 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M17 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_4 N_56 GND mn5  l=0.5u w=0.5u m=1
M20 N_57 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M21 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M23 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M24 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M25 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M26 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M28 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_4 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M34 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M44 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M45 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M46 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M47 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M48 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdbfb1
* SPICE INPUT		Wed Jul 10 14:00:35 2019	sdbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb2
.subckt sdbfb2 VDD Q QN GND RN SN SI SE D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_5 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_4 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_4 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M20 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M21 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M22 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M23 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M24 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M25 N_4 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.52u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M42 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M44 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M45 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M46 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M47 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M48 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdbfb2
* SPICE INPUT		Wed Jul 10 14:00:42 2019	sdbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb1
.subckt sdbrb1 VDD Q QN GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M18 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M19 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M20 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M21 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M22 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M23 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M24 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M42 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M44 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M45 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M46 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M47 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M48 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdbrb1
* SPICE INPUT		Wed Jul 10 14:00:50 2019	sdbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb2
.subckt sdbrb2 VDD Q QN GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M18 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M20 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M21 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M22 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M23 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M24 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M43 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M44 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M45 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M46 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M47 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M48 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
.ends sdbrb2
* SPICE INPUT		Wed Jul 10 14:00:57 2019	sdbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq1
.subckt sdbrq1 VDD Q GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_35 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_35 N_6 N_30 GND mn5  l=0.5u w=0.5u m=1
M6 N_36 SI N_30 GND mn5  l=0.5u w=0.5u m=1
M7 N_36 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_30 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_37 GND mn5  l=0.5u w=0.5u m=1
M10 N_37 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_28 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_28 N_3 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_38 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_38 GND mn5  l=0.5u w=0.5u m=1
M16 Q N_11 N_24 GND mn5  l=0.5u w=0.58u m=1
M17 N_24 N_3 Q GND mn5  l=0.5u w=0.58u m=1
M18 N_24 SN GND GND mn5  l=0.5u w=0.58u m=1
M19 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M20 N_39 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M21 N_39 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_12 N_3 N_26 GND mn5  l=0.5u w=0.5u m=1
M23 N_26 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M24 N_26 SN GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_22 N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M42 Q N_3 N_22 VDD mp5  l=0.42u w=0.76u m=1
M43 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M44 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M45 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M46 N_21 N_3 N_12 VDD mp5  l=0.42u w=0.5u m=1
M47 N_21 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M48 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdbrq1
* SPICE INPUT		Wed Jul 10 14:01:05 2019	sdbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq2
.subckt sdbrq2 VDD Q GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_35 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_35 N_6 N_30 GND mn5  l=0.5u w=0.5u m=1
M6 N_36 SI N_30 GND mn5  l=0.5u w=0.5u m=1
M7 N_36 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_30 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_37 GND mn5  l=0.5u w=0.5u m=1
M10 N_37 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_28 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_28 N_3 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_38 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_12 N_3 N_26 GND mn5  l=0.5u w=0.5u m=1
M16 N_26 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M17 N_26 SN GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 N_24 GND mn5  l=0.5u w=0.72u m=1
M19 N_24 N_3 Q GND mn5  l=0.5u w=0.72u m=1
M20 N_24 SN GND GND mn5  l=0.5u w=0.72u m=1
M21 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M22 N_11 N_5 N_38 GND mn5  l=0.5u w=0.5u m=1
M23 N_39 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M24 N_39 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_21 N_3 N_12 VDD mp5  l=0.42u w=0.5u m=1
M41 N_21 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M42 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M43 N_22 N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M44 Q N_3 N_22 VDD mp5  l=0.42u w=0.96u m=1
M45 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M46 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M47 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M48 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdbrq2
* SPICE INPUT		Wed Jul 10 14:01:12 2019	sdcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb1
.subckt sdcfb1 VDD Q QN GND RN SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_26 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M6 N_47 SI N_26 GND mn5  l=0.5u w=0.5u m=1
M7 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M9 N_48 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_11 N_5 N_49 GND mn5  l=0.5u w=0.5u m=1
M15 N_50 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M16 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M20 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M28 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M32 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M35 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M37 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M38 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M41 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M42 N_14 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M43 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M44 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends sdcfb1
* SPICE INPUT		Wed Jul 10 14:01:19 2019	sdcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb2
.subckt sdcfb2 VDD Q QN GND CKN D SE SI RN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M5 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M10 N_11 N_5 N_49 GND mn5  l=0.5u w=0.5u m=1
M11 N_50 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M12 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_28 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M14 N_47 SI N_28 GND mn5  l=0.5u w=0.5u m=1
M15 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M17 N_48 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 N_14 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M31 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M33 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M35 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M39 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M44 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdcfb2
* SPICE INPUT		Wed Jul 10 14:01:27 2019	sdcfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfq1
.subckt sdcfq1 VDD Q GND CKN D SE SI RN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_5 N_47 GND mn5  l=0.5u w=0.5u m=1
M4 N_48 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M6 N_48 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_44 D GND GND mn5  l=0.5u w=0.5u m=1
M10 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M11 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M13 N_27 N_6 N_44 GND mn5  l=0.5u w=0.5u m=1
M14 N_45 SI N_27 GND mn5  l=0.5u w=0.5u m=1
M15 N_45 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_4 N_27 GND mn5  l=0.5u w=0.5u m=1
M17 N_46 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_47 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M25 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_21 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_12 N_13 N_22 VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M33 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M38 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_10 N_13 N_19 VDD mp5  l=0.42u w=0.52u m=1
M41 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcfq1
* SPICE INPUT		Wed Jul 10 14:01:34 2019	sdcfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfq2
.subckt sdcfq2 VDD Q GND RN SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_48 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_48 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_44 D GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M12 N_25 N_6 N_44 GND mn5  l=0.5u w=0.5u m=1
M13 N_45 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M14 N_45 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M16 N_46 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_47 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_11 N_5 N_47 GND mn5  l=0.5u w=0.5u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_21 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_12 N_13 N_22 VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M30 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M37 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M38 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_10 N_13 N_19 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
.ends sdcfq2
* SPICE INPUT		Wed Jul 10 14:01:41 2019	sdcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb1
.subckt sdcrb1 VDD Q QN GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M5 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_50 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M13 N_11 N_4 N_49 GND mn5  l=0.5u w=0.5u m=1
M14 N_26 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M15 N_47 SI N_26 GND mn5  l=0.5u w=0.5u m=1
M16 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_5 N_26 GND mn5  l=0.5u w=0.5u m=1
M18 N_48 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M19 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M31 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M35 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M40 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M41 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M44 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrb1
* SPICE INPUT		Wed Jul 10 14:01:49 2019	sdcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb2
.subckt sdcrb2 VDD Q QN GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M5 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_50 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M13 N_11 N_4 N_49 GND mn5  l=0.5u w=0.5u m=1
M14 N_26 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M15 N_47 SI N_26 GND mn5  l=0.5u w=0.5u m=1
M16 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_5 N_26 GND mn5  l=0.5u w=0.5u m=1
M18 N_48 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M19 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M31 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M35 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M40 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M41 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M44 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrb2
* SPICE INPUT		Wed Jul 10 14:01:56 2019	sdcrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrn1
.subckt sdcrn1 VDD QN GND RN SI SE D CK
M1 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_42 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M9 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_24 N_6 N_42 GND mn5  l=0.5u w=0.5u m=1
M13 N_43 SI N_24 GND mn5  l=0.5u w=0.5u m=1
M14 N_43 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_5 N_24 GND mn5  l=0.5u w=0.5u m=1
M16 N_44 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_44 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M21 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M28 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_21 VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_10 N_13 N_18 VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrn1
* SPICE INPUT		Wed Jul 10 14:02:03 2019	sdcrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrn2
.subckt sdcrn2 VDD QN GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_42 D GND GND mn5  l=0.5u w=0.5u m=1
M5 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_24 N_6 N_42 GND mn5  l=0.5u w=0.5u m=1
M9 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M12 N_43 SI N_24 GND mn5  l=0.5u w=0.5u m=1
M13 N_43 SE GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_5 N_24 GND mn5  l=0.5u w=0.5u m=1
M15 N_44 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M16 N_44 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M26 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_12 N_13 N_21 VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_21 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M36 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 N_13 N_18 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
.ends sdcrn2
* SPICE INPUT		Wed Jul 10 14:02:11 2019	sdcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq1
.subckt sdcrq1 VDD Q GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_12 GND GND mn5  l=0.5u w=0.58u m=1
M4 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_13 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 RN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_47 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_43 D GND GND mn5  l=0.5u w=0.5u m=1
M10 N_47 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M11 N_11 N_4 N_46 GND mn5  l=0.5u w=0.5u m=1
M12 N_25 N_6 N_43 GND mn5  l=0.5u w=0.5u m=1
M13 N_44 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M14 N_44 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M16 N_45 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M24 Q N_12 N_15 VDD mp5  l=0.42u w=0.76u m=1
M25 N_15 N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_12 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_21 N_13 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M32 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M33 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M38 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_10 N_12 N_19 VDD mp5  l=0.42u w=0.52u m=1
M41 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_22 N_12 N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrq1
* SPICE INPUT		Wed Jul 10 14:02:18 2019	sdcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq2
.subckt sdcrq2 VDD Q GND RN SI SE D CK
M1 N_12 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M4 Q N_12 GND GND mn5  l=0.5u w=0.72u m=1
M5 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_13 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_47 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_43 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_47 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M12 N_11 N_4 N_46 GND mn5  l=0.5u w=0.5u m=1
M13 N_25 N_6 N_43 GND mn5  l=0.5u w=0.5u m=1
M14 N_44 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M15 N_44 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_45 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_12 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q N_12 N_15 VDD mp5  l=0.42u w=0.96u m=1
M26 N_15 N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_22 N_12 N_13 VDD mp5  l=0.42u w=0.52u m=1
M30 N_21 N_13 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M33 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M34 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M38 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M39 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 N_12 N_19 VDD mp5  l=0.42u w=0.52u m=1
M42 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrq2
* SPICE INPUT		Wed Jul 10 14:02:25 2019	sdnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb1
.subckt sdnfb1 GND QN Q VDD SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M6 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M7 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_17 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_11 N_5 N_18 GND mn5  l=0.5u w=0.5u m=1
M14 N_19 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M15 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M18 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M19 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M24 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M25 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_9 N_5 N_21 VDD mp5  l=0.42u w=0.52u m=1
M27 N_40 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M28 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_41 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M32 N_42 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M33 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M36 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends sdnfb1
* SPICE INPUT		Wed Jul 10 14:02:33 2019	sdnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb2
.subckt sdnfb2 GND QN Q VDD SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_19 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_5 N_18 GND mn5  l=0.5u w=0.5u m=1
M10 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M14 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_17 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M22 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M24 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_42 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_41 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M29 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M32 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M33 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_9 N_5 N_21 VDD mp5  l=0.42u w=0.52u m=1
M35 N_40 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M36 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdnfb2
* SPICE INPUT		Wed Jul 10 14:02:40 2019	sdnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb1
.subckt sdnrb1 GND QN Q VDD SI SE D CK
M1 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M3 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 N_4 N_18 GND mn5  l=0.5u w=0.5u m=1
M8 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M10 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M13 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M14 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M16 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M18 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M19 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_42 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M25 N_41 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M26 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M33 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M34 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_9 N_4 N_21 VDD mp5  l=0.42u w=0.52u m=1
M36 N_40 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
.ends sdnrb1
* SPICE INPUT		Wed Jul 10 14:02:47 2019	sdnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb2
.subckt sdnrb2 GND QN Q VDD SI SE D CK
M1 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_19 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 N_4 N_18 GND mn5  l=0.5u w=0.5u m=1
M6 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M8 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M14 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M19 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_42 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M23 N_41 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M24 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M31 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M32 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_9 N_4 N_21 VDD mp5  l=0.42u w=0.52u m=1
M34 N_40 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdnrb2
* SPICE INPUT		Wed Jul 10 14:02:54 2019	sdnrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrn1
.subckt sdnrn1 GND QN VDD SI SE D CK
M1 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M7 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M9 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M12 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M13 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M14 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M15 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M16 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M18 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M23 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M24 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_20 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_37 N_6 N_20 VDD mp5  l=0.42u w=0.52u m=1
M32 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_9 N_4 N_20 VDD mp5  l=0.42u w=0.52u m=1
M34 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
.ends sdnrn1
* SPICE INPUT		Wed Jul 10 14:03:02 2019	sdnrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrn2
.subckt sdnrn2 GND QN VDD CK D SE SI
M1 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M14 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M21 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M22 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M27 N_9 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M28 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_37 N_6 N_22 VDD mp5  l=0.42u w=0.52u m=1
M30 N_22 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdnrn2
* SPICE INPUT		Wed Jul 10 14:03:09 2019	sdnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq1
.subckt sdnrq1 GND Q VDD CK D SE SI
M1 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M2 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M10 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M12 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M13 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M14 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M19 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M20 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M24 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_9 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M26 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M29 N_37 N_6 N_22 VDD mp5  l=0.42u w=0.52u m=1
M30 N_22 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdnrq1
* SPICE INPUT		Wed Jul 10 14:03:16 2019	sdnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq2
.subckt sdnrq2 GND Q VDD CK D SE SI
M1 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M5 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M14 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M21 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M23 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M27 N_9 N_4 N_19 VDD mp5  l=0.42u w=0.52u m=1
M28 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_37 N_6 N_19 VDD mp5  l=0.42u w=0.52u m=1
M30 N_19 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdnrq2
* SPICE INPUT		Wed Jul 10 14:03:23 2019	sdpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb1
.subckt sdpfb1 VDD Q QN GND CKN D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.58u m=1
M2 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M5 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_46 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_5 N_45 GND mn5  l=0.5u w=0.5u m=1
M9 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M11 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_43 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M15 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M18 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.76u m=1
M23 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M25 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M29 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M30 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M38 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M39 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdpfb1
* SPICE INPUT		Wed Jul 10 14:03:31 2019	sdpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb2
.subckt sdpfb2 VDD Q QN GND CKN D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_46 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M5 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_5 N_45 GND mn5  l=0.5u w=0.5u m=1
M7 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M9 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M10 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_43 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M15 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M18 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.96u m=1
M23 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M28 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M32 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M38 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M39 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdpfb2
* SPICE INPUT		Wed Jul 10 14:03:38 2019	sdprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb1
.subckt sdprb1 VDD Q QN GND CK D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M5 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M10 N_43 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M12 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M13 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M15 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M18 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.76u m=1
M23 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M28 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M32 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M33 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M35 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M38 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M39 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprb1
* SPICE INPUT		Wed Jul 10 14:03:45 2019	sdprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb2
.subckt sdprb2 VDD Q QN GND CK D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M7 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M9 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_43 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M12 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M13 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M14 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M15 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M18 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.96u m=1
M23 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M28 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M32 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M33 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M35 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M36 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M38 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M39 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M41 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprb2
* SPICE INPUT		Wed Jul 10 14:03:53 2019	sdprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq1
.subckt sdprq1 VDD Q GND CK D SN SE SI
M1 N_43 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M2 N_43 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_42 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_44 SN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_41 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_4 N_42 GND mn5  l=0.5u w=0.5u m=1
M7 N_41 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_11 N_44 GND mn5  l=0.5u w=0.5u m=1
M9 Q N_11 N_37 GND mn5  l=0.5u w=0.58u m=1
M10 N_40 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_40 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M12 N_9 N_5 N_24 GND mn5  l=0.5u w=0.5u m=1
M13 N_37 SN GND GND mn5  l=0.5u w=0.58u m=1
M14 N_39 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_39 SI N_24 GND mn5  l=0.5u w=0.5u m=1
M16 N_24 N_6 N_38 GND mn5  l=0.5u w=0.5u m=1
M17 N_38 D GND GND mn5  l=0.5u w=0.5u m=1
M18 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M19 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M20 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_18 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_17 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M23 N_17 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_18 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M29 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_16 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_16 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M32 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M33 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M34 N_15 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_15 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_7 SE N_14 VDD mp5  l=0.42u w=0.5u m=1
M37 N_14 D VDD VDD mp5  l=0.42u w=0.5u m=1
M38 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprq1
* SPICE INPUT		Wed Jul 10 14:04:00 2019	sdprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq2
.subckt sdprq2 GND Q VDD CK D SE SI SN
M1 N_20 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_20 N_4 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 N_3 N_19 GND mn5  l=0.5u w=0.5u m=1
M4 N_19 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_18 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_18 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 Q N_10 N_14 GND mn5  l=0.5u w=0.72u m=1
M10 N_17 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M12 N_14 SN GND GND mn5  l=0.5u w=0.72u m=1
M13 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M14 N_16 SI N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_6 N_5 N_15 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 SE GND GND mn5  l=0.5u w=0.5u m=1
M19 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M20 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_44 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_44 N_3 N_10 VDD mp5  l=0.42u w=0.5u m=1
M23 N_43 N_4 N_10 VDD mp5  l=0.42u w=0.52u m=1
M24 N_43 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_9 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_42 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 Q N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_11 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_42 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M31 N_8 N_3 N_25 VDD mp5  l=0.42u w=0.5u m=1
M32 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M33 N_41 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_41 N_5 N_25 VDD mp5  l=0.42u w=0.5u m=1
M35 N_11 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M36 N_25 SE N_40 VDD mp5  l=0.42u w=0.5u m=1
M37 N_40 D VDD VDD mp5  l=0.42u w=0.5u m=1
M38 N_5 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprq2
* SPICE INPUT		Wed Jul 10 14:04:07 2019	tiehi
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tiehi
.subckt tiehi VDD Y GND
M1 N_5 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends tiehi
* SPICE INPUT		Wed Jul 10 14:04:14 2019	tielo
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tielo
.subckt tielo GND Y VDD
M1 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_5 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends tielo
* SPICE INPUT		Wed Jul 10 14:04:22 2019	tlatncad1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad1
.subckt tlatncad1 VDD ECK GND CK E
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_21 E GND GND mn5  l=0.5u w=0.5u m=1
M3 N_21 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_22 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_22 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 ECK N_5 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_6 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_3 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_9 E VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_10 N_3 N_5 VDD mp5  l=0.42u w=0.5u m=1
M13 N_9 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M14 N_10 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M15 N_11 N_5 ECK VDD mp5  l=0.42u w=0.76u m=1
M16 N_6 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_11 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends tlatncad1
* SPICE INPUT		Wed Jul 10 14:04:29 2019	tlatncad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad2
.subckt tlatncad2 VDD ECK GND CK E
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_21 E GND GND mn5  l=0.5u w=0.5u m=1
M3 N_21 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_22 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_22 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 ECK N_5 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_6 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M8 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M9 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M10 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_9 E VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_10 N_3 N_5 VDD mp5  l=0.42u w=0.5u m=1
M13 N_9 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M14 N_10 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M15 N_11 N_5 ECK VDD mp5  l=0.42u w=0.96u m=1
M16 N_6 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_11 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends tlatncad2
* SPICE INPUT		Wed Jul 10 14:04:36 2019	tlatncad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad4
.subckt tlatncad4 GND ECK VDD E CK
M1 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 ECK N_5 GND GND mn5  l=0.5u w=0.72u m=1
M5 ECK N_5 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_10 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M10 N_10 E GND GND mn5  l=0.5u w=0.5u m=1
M11 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_6 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_28 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_27 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M18 N_28 N_3 N_5 VDD mp5  l=0.42u w=0.5u m=1
M19 N_27 E VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_15 N_5 ECK VDD mp5  l=0.42u w=0.96u m=1
M22 ECK N_5 N_15 VDD mp5  l=0.42u w=0.96u m=1
.ends tlatncad4
* SPICE INPUT		Wed Jul 10 14:04:43 2019	tlatntscad1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad1
.subckt tlatntscad1 VDD ECK GND CK SE E
M1 N_4 E GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 SE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_27 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M7 N_28 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_28 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_7 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_8 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 ECK N_3 GND GND mn5  l=0.5u w=0.58u m=1
M12 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M13 N_11 E N_4 VDD mp5  l=0.42u w=0.52u m=1
M14 N_11 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_6 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_12 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_13 N_3 N_7 VDD mp5  l=0.42u w=0.5u m=1
M19 N_12 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_7 ECK VDD mp5  l=0.42u w=0.76u m=1
M22 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M24 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends tlatntscad1
* SPICE INPUT		Wed Jul 10 14:04:51 2019	tlatntscad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad2
.subckt tlatntscad2 VDD ECK GND CK SE E
M1 N_4 E GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 SE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_28 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_29 N_6 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_8 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M11 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M12 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M13 N_12 E N_4 VDD mp5  l=0.42u w=0.52u m=1
M14 N_12 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 VDD N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M17 N_13 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_14 N_3 N_8 VDD mp5  l=0.42u w=0.5u m=1
M19 N_13 N_6 N_8 VDD mp5  l=0.42u w=0.52u m=1
M20 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_15 N_8 ECK VDD mp5  l=0.42u w=0.96u m=1
M22 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M24 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends tlatntscad2
* SPICE INPUT		Wed Jul 10 14:04:58 2019	tlatntscad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad4
.subckt tlatntscad4 GND ECK VDD CK SE E
M1 N_4 E GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 SE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_12 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_7 GND GND mn5  l=0.5u w=0.72u m=1
M10 ECK N_7 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_8 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M13 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M14 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M15 ECK N_7 N_15 VDD mp5  l=0.42u w=0.96u m=1
M16 ECK N_7 N_15 VDD mp5  l=0.42u w=0.96u m=1
M17 N_33 E N_4 VDD mp5  l=0.42u w=0.52u m=1
M18 N_33 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 VDD N_3 N_6 VDD mp5  l=0.42u w=0.52u m=1
M21 N_34 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_35 N_3 N_7 VDD mp5  l=0.42u w=0.5u m=1
M23 N_34 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M24 N_35 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_15 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends tlatntscad4
* SPICE INPUT		Wed Jul 10 14:05:05 2019	xn02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d0
.subckt xn02d0 VDD Y GND A B
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_8 A N_6 VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends xn02d0
* SPICE INPUT		Wed Jul 10 14:05:12 2019	xn02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d1
.subckt xn02d1 VDD Y GND A B
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A N_4 GND mn5  l=0.5u w=0.5u m=1
M5 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M8 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_8 A N_6 VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends xn02d1
* SPICE INPUT		Wed Jul 10 14:05:19 2019	xn02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d2
.subckt xn02d2 VDD Y GND A B
M1 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A N_4 GND mn5  l=0.5u w=0.5u m=1
M6 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_7 N_5 N_4 VDD mp5  l=0.42u w=0.52u m=1
M11 N_8 A N_7 VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends xn02d2
* SPICE INPUT		Wed Jul 10 14:05:26 2019	xn03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d0
.subckt xn03d0 VDD Y GND C B A
M1 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M8 Y N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_9 C N_12 GND mn5  l=0.5u w=0.5u m=1
M11 N_12 N_11 N_6 GND mn5  l=0.5u w=0.5u m=1
M12 N_11 C VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.52u m=1
M16 N_9 B N_4 VDD mp5  l=0.42u w=0.52u m=1
M17 N_6 B N_5 VDD mp5  l=0.42u w=0.52u m=1
M18 N_10 B VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 C N_12 VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 N_11 N_12 VDD mp5  l=0.42u w=0.52u m=1
.ends xn03d0
* SPICE INPUT		Wed Jul 10 14:05:34 2019	xn03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d1
.subckt xn03d1 VDD Y GND C A B
M1 N_12 N_11 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_9 C N_12 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M6 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M8 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M10 Y N_12 GND GND mn5  l=0.5u w=0.58u m=1
M11 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M12 N_11 C VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_9 B N_4 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 B N_5 VDD mp5  l=0.42u w=0.52u m=1
M15 N_10 B VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 C N_12 VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 N_11 N_12 VDD mp5  l=0.42u w=0.52u m=1
.ends xn03d1
* SPICE INPUT		Wed Jul 10 14:05:41 2019	xn03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d2
.subckt xn03d2 VDD Y GND C A B
M1 N_12 N_11 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_9 C N_12 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M6 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M8 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M10 Y N_12 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M12 N_11 C VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_9 B N_4 VDD mp5  l=0.42u w=0.52u m=1
M14 N_6 B N_5 VDD mp5  l=0.42u w=0.52u m=1
M15 N_10 B VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.52u m=1
M17 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Y N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 C N_12 VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 N_11 N_12 VDD mp5  l=0.42u w=0.52u m=1
.ends xn03d2
* SPICE INPUT		Wed Jul 10 14:05:48 2019	xr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d0
.subckt xr02d0 VDD Y GND B A
M1 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_6 N_5 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_4 A N_6 VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_8 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends xr02d0
* SPICE INPUT		Wed Jul 10 14:05:55 2019	xr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d1
.subckt xr02d1 VDD Y GND B A
M1 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_6 N_5 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_4 A N_6 VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M11 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_8 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends xr02d1
* SPICE INPUT		Wed Jul 10 14:06:02 2019	xr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d2
.subckt xr02d2 VDD Y GND B A
M1 N_5 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_8 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A N_7 GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_5 N_4 GND mn5  l=0.5u w=0.5u m=1
M7 N_7 A N_4 VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 N_8 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_8 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
.ends xr02d2
* SPICE INPUT		Wed Jul 10 14:06:10 2019	xr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d0
.subckt xr03d0 VDD Y GND C B A
M1 N_9 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 C N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M9 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M10 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M11 Y N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_4 A VDD VDD mp5  l=0.42u w=0.5u m=1
M13 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M14 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.5u m=1
M15 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.5u m=1
M16 N_9 B N_4 VDD mp5  l=0.42u w=0.5u m=1
M17 N_6 B N_5 VDD mp5  l=0.42u w=0.5u m=1
M18 N_10 B VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_11 C VDD VDD mp5  l=0.42u w=0.5u m=1
M20 Y N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 N_11 N_12 VDD mp5  l=0.42u w=0.5u m=1
M22 N_9 C N_12 VDD mp5  l=0.42u w=0.5u m=1
.ends xr03d0
* SPICE INPUT		Wed Jul 10 14:06:17 2019	xr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d1
.subckt xr03d1 VDD Y GND C A B
M1 N_9 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 C N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 Y N_12 GND GND mn5  l=0.5u w=0.58u m=1
M9 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M12 N_9 B N_4 VDD mp5  l=0.42u w=0.5u m=1
M13 N_6 B N_5 VDD mp5  l=0.42u w=0.5u m=1
M14 N_10 B VDD VDD mp5  l=0.42u w=0.5u m=1
M15 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.5u m=1
M16 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.5u m=1
M17 Y N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 N_4 A VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_11 C VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_6 N_11 N_12 VDD mp5  l=0.42u w=0.5u m=1
M22 N_9 C N_12 VDD mp5  l=0.42u w=0.5u m=1
.ends xr03d1
* SPICE INPUT		Wed Jul 10 14:06:24 2019	xr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d2
.subckt xr03d2 VDD Y GND A B C
M1 N_9 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 C N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_4 B N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 B GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 N_10 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_6 N_10 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 Y N_12 GND GND mn5  l=0.5u w=0.72u m=1
M9 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M10 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_11 C GND GND mn5  l=0.5u w=0.5u m=1
M12 N_9 B N_4 VDD mp5  l=0.42u w=0.5u m=1
M13 N_6 B N_5 VDD mp5  l=0.42u w=0.5u m=1
M14 N_10 B VDD VDD mp5  l=0.42u w=0.5u m=1
M15 N_9 N_10 N_5 VDD mp5  l=0.42u w=0.5u m=1
M16 N_4 N_10 N_6 VDD mp5  l=0.42u w=0.5u m=1
M17 Y N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 N_4 A VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_11 C VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_6 N_11 N_12 VDD mp5  l=0.42u w=0.5u m=1
M22 N_9 C N_12 VDD mp5  l=0.42u w=0.5u m=1
.ends xr03d2
