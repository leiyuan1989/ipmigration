//* 
//* No part of this file can be released without the consent of SMIC.
//*
//******************************************************************************************
//* 0.11um Mixed Signal 1P8M with MIM Salicide 1.2V/3.3V RF SPICE Model (for SPECTRE only) *
//******************************************************************************************
//*
//* Release version    : 1.14
//*
//* Release date       : 03/30/2016
//*
//* Simulation tool    : Cadence spectre V10.1
//*
//*
//*  Resistor   :
//*        *------------------------------------------------------------------* 
//*        |                 |                Resistor subckt                 |
//*        *==================================================================*
//*        | N+ poly SAB     |    rnposab_ckt_rf     |    rnposab_ckt_rf_3t   |
//*        *------------------------------------------------------------------*
//*        | p+ poly SAB     |    rpposab_ckt_rf     |    rpposab_ckt_rf_3t   |
//*        *------------------------------------------------------------------*
//*        | HRP poly        |    rhrpo_ckt_rf      |     rhrpo_ckt_rf_3t     |
//*        *------------------------------------------------------------------*
//*
//*
simulator lang=spectre  insensitive=yes
ahdl_include "res_rf.va"
//************************************             
//* Non-silicide N+ poly resistor             
//************************************             
//* l=length, w=width                          
subckt rnposab_ckt_rf (port1 port2)               
parameters l=0 w=0 devt=temp mismod_res_rf=0
//*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = 1/sqrt(weff*leff)
+arsh = 1.0E-05

+  rtc1 = -9.93E-04    rtc2 = 1.07E-06
+ dw = 1.68E-08-2.7E-9+ddw_rnposab_rf   dl = -1.33e-7
+tref = 25                    rsh = 275.50+drsh_rnposab_rf+rshmis
//+vc1 = -5.53E-05            vc2 = -5.75E-04
+ rjc1a = 3.04E-05            rjc1b = -3.29E-09
+ rjc2a = -1.18E-08           rjc2b = -2.99E-13
+weff     = w*0.9-2*dw       leff   = l*0.9-2*dl
//RF component value
+ls_rf      = max((0.007035*pwr(w*0.9*1e6+0.19294,1.0366)*(0.135+pwr((l*0.9)/(w*0.9)+0.2,-2.221*pwr(w*0.9*1e6,-0.1078)+4.864)))*1e-9,1e-12)
+cf_rf      = max((0.08566*pwr(w*0.9*1e6+0.2,-0.8872)*(0.006+pwr((l*0.9)/(w*0.9)+0.0202,0.2368*pwr(w*0.9*1e6,-1.7352)-3.026)))*1e-15,1e-18)
+rsub_rf    = max(165.3+2389.6*pwr(w*0.9*1e6,-0.9242)+174.3*pwr(w*0.9*1e6+2.0705,4)*pwr(l*0.9*1e6+0.02666,-0.4314*pwr(w*0.9*1e6,1.2708)-1.916),1e-5)
+csub_rf    = max((0.03194*pwr(w*0.9*1e6+0.2,1.5946)*(6.783+pwr(l*0.9*w*0.9*1e12+0.13226,-0.347*pwr(w*0.9*1e6,0.87)+1.4215)))*1e-15,1e-18)
+cox_rf     = max((0.01085*pwr(w*0.9*1e6+0.2,0.5126)*(10+pwr(l*0.9*w*0.9*1e12+0.4065,0.9025*pwr(w*0.9*1e6,-1.7592)+1.0813)))*1e-15,1e-18)
+rs2_rf     = max(0.39+0.44455*pwr(w*0.9*1e6+0.13192,-0.3454)*(0.155+exp(5+0.06201*(pwr(w*0.9*1e6,1.26)+3.094)*(l*0.9)/(w*0.9))),1e-5)
//*equivalent circuit
ls    (1 port2) inductor   l=ls_rf
cf    (port1 1) capacitor  c=cf_rf
rs    (port1 1 port1 1)    polyres_rf_hdl lr=l wr=w rtemp=devt etch=dw etchl=dl tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rminvcoef=0.834
rs2   (1 port2) resistor   r=rs2_rf
rsub1 (2 0)     resistor   r=rsub_rf
csub1 (2 0)     capacitor  c=csub_rf
cox1  (port1 2) capacitor  c=cox_rf
rsub2 (3 0)     resistor   r=rsub_rf
csub2 (3 0)     capacitor  c=csub_rf
cox2  (port2 3) capacitor  c=cox_rf
ends rnposab_ckt_rf 
//*   
//*************************************************
//* Non-silicide N+ poly resistor (three terminal)          
//*************************************************
//* l=length, w=width                          
subckt rnposab_ckt_rf_3t (port1 port2 pwell)               
parameters l=0 w=0 devt=temp mismod_res_rf=0  
//*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = 1/sqrt(weff*leff)
+arsh = 1.0E-05

+  rtc1 = -9.93E-04    rtc2 = 1.07E-06
+ dw = 1.68E-08-2.7E-9+ddw_rnposab_rf   dl = -1.33e-7
+tref = 25                    rsh = 275.50+drsh_rnposab_rf+rshmis
+weff     = w*0.9-2*dw       leff   = l*0.9-2*dl
//+vc1 = -5.53E-05            vc2 = -5.75E-04
+ rjc1a = 3.04E-05            rjc1b = -3.29E-09
+ rjc2a = -1.18E-08           rjc2b = -2.99E-13
//RF component value
+ls_rf      = max((0.007035*pwr(w*0.9*1e6+0.19294,1.0366)*(0.135+pwr((l*0.9)/(w*0.9)+0.2,-2.221*pwr(w*0.9*1e6,-0.1078)+4.864)))*1e-9,1e-12)
+cf_rf      = max((0.08566*pwr(w*0.9*1e6+0.2,-0.8872)*(0.006+pwr((l*0.9)/(w*0.9)+0.0202,0.2368*pwr(w*0.9*1e6,-1.7352)-3.026)))*1e-15,1e-18)
+rsub_rf    = max(165.3+2389.6*pwr(w*0.9*1e6,-0.9242)+174.3*pwr(w*0.9*1e6+2.0705,4)*pwr(l*0.9*1e6+0.02666,-0.4314*pwr(w*0.9*1e6,1.2708)-1.916),1e-5)
+csub_rf    = max((0.03194*pwr(w*0.9*1e6+0.2,1.5946)*(6.783+pwr(l*0.9*w*0.9*1e12+0.13226,-0.347*pwr(w*0.9*1e6,0.87)+1.4215)))*1e-15,1e-18)
+cox_rf     = max((0.01085*pwr(w*0.9*1e6+0.2,0.5126)*(10+pwr(l*0.9*w*0.9*1e12+0.4065,0.9025*pwr(w*0.9*1e6,-1.7592)+1.0813)))*1e-15,1e-18)
+rs2_rf     = max(0.39+0.44455*pwr(w*0.9*1e6+0.13192,-0.3454)*(0.155+exp(5+0.06201*(pwr(w*0.9*1e6,1.26)+3.094)*(l*0.9)/(w*0.9))),1e-5)
//*equivalent circuit
ls    (1 port2) inductor   l=ls_rf
cf    (port1 1) capacitor  c=cf_rf
rs    (port1 1 port1 1)    polyres_rf_hdl lr=l wr=w rtemp=devt etch=dw etchl=dl tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rminvcoef=0.834
rs2   (1 port2) resistor   r=rs2_rf
rsub1 (2 pwell)     resistor   r=rsub_rf
csub1 (2 pwell)     capacitor  c=csub_rf
cox1  (port1 2) capacitor  c=cox_rf
rsub2 (3 pwell)     resistor   r=rsub_rf
csub2 (3 pwell)     capacitor  c=csub_rf
cox2  (port2 3) capacitor  c=cox_rf
ends rnposab_ckt_rf_3t 
//* 
//************************************             
//* Non-silicide P+ poly resistor             
//************************************             
//* l=length, w=width                            
subckt rpposab_ckt_rf (port1 port2)               
parameters l=0 w=0 devt=temp mismod_res_rf=0  
//*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = 1/sqrt(weff*leff)
+arsh = 3.4E-06

+  rtc1 = -5.75E-05    rtc2 = 6.10E-07
+ dw = 1.28E-08-2.7E-9+ddw_rpposab_rf   dl = -2.68e-7
+tref = 25                    rsh = 321.5+drsh_rpposab_rf+rshmis
+weff     = w*0.9-2*dw       leff   = l*0.9-2*dl
//+vc1 = -5.07E-05            vc2 = -7.96E-05
+ rjc1a = 2.16E-05            rjc1b = -1.77E-9
+ rjc2a = -7.61E-10           rjc2b = -1.79E-14
//RF component value
+ls_rf      = max(((0.0129*w*1e6+0.0006)*pwr(l/w,2.3758*pwr(w*1e6,0.1048)))*1e-9,1e-12)
+cf_rf      = max((0.8913*pwr(l/w,-1.1526))*1e-15,1e-18)
+rsub_rf    = max(71.885*l/w + 70.958,1e-3)
+csub_rf    = max((1.5*pwr(l/w,0.4337))*1e-15,1e-18)
+cox_rf     = max((0.046*w*l*1e12+1.5358)*1e-15,1e-18)
+rs2_rf     = max(2000*l/w,1e-5)
//*equivalent circuit
ls    (1 port2) inductor   l=ls_rf
cf    (port1 1) capacitor  c=cf_rf
rs    (port1 1 port1 1)    polyres_rf_hdl lr=l wr=w rtemp=devt etch=dw etchl=dl tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rminvcoef=0.890
rs2   (1 port2) resistor   r=rs2_rf
Cf2   (port1 4) capacitor  c=(Cf_rf*0.1)
Rs3   (4 port2) resistor   r=(Rs2_rf*10)
rsub1 (2 0)     resistor   r=rsub_rf
csub1 (2 0)     capacitor  c=csub_rf
cox1  (port1 2) capacitor  c=cox_rf
rsub2 (3 0)     resistor   r=rsub_rf
csub2 (3 0)     capacitor  c=csub_rf
cox2  (port2 3) capacitor  c=cox_rf
ends rpposab_ckt_rf 
//*      
//*************************************************
//* Non-silicide P+ poly resistor (three terminal)
//*************************************************
//* l=length, w=width                            
subckt rpposab_ckt_rf_3t (port1 port2 pwell)               
parameters l=0 w=0 devt=temp mismod_res_rf=0  
//*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = 1/sqrt(weff*leff)
+arsh = 3.4E-06

+  rtc1 = -5.75E-05    rtc2 = 6.10E-07
+ dw = 1.28E-08-2.7E-9+ddw_rpposab_rf   dl = -2.68e-7
+tref = 25                    rsh = 321.5+drsh_rpposab_rf+rshmis
+weff     = w*0.9-2*dw       leff   = l*0.9-2*dl
//+vc1 = -5.07E-05            vc2 = -7.96E-05
+ rjc1a = 2.16E-05            rjc1b = -1.77E-9
+ rjc2a = -7.61E-10           rjc2b = -1.79E-14
//RF component value
+ls_rf      = max(((0.0129*w*1e6+0.0006)*pwr(l/w,2.3758*pwr(w*1e6,0.1048)))*1e-9,1e-12)
+cf_rf      = max((0.8913*pwr(l/w,-1.1526))*1e-15,1e-18)
+rsub_rf    = max(71.885*l/w + 70.958,1e-3)
+csub_rf    = max((1.5*pwr(l/w,0.4337))*1e-15,1e-18)
+cox_rf     = max((0.046*w*l*1e12+1.5358)*1e-15,1e-18)
+rs2_rf     = max(2000*l/w,1e-5)
//*equivalent circuit
ls    (1 port2) inductor   l=ls_rf
cf    (port1 1) capacitor  c=cf_rf
rs    (port1 1 port1 1)    polyres_rf_hdl lr=l wr=w rtemp=devt etch=dw etchl=dl tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rminvcoef=0.890
rs2   (1 port2) resistor   r=rs2_rf
Cf2   (port1 4) capacitor  c=(Cf_rf*0.1)
Rs3   (4 port2) resistor   r=(Rs2_rf*10)
rsub1 (2 pwell) resistor   r=rsub_rf
csub1 (2 pwell) capacitor  c=csub_rf
cox1  (port1 2) capacitor  c=cox_rf
rsub2 (3 pwell) resistor   r=rsub_rf
csub2 (3 pwell) capacitor  c=csub_rf
cox2  (port2 3) capacitor  c=cox_rf
ends rpposab_ckt_rf_3t 
//*
//*                                                     
//******************************************************************
//*                non-silicide HR poly resistance                 *
//******************************************************************
subckt rhrpo_ckt_rf (port1 port2)
parameters l=0 w=0 mismod_res_rf=0
+devt=temp
//*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = 1/sqrt(weff*l*0.9)
+arsh = 1.55E-05
//
+ rtc1 = -6.77E-04 rtc2 = 2.08E-06
+ dw = 2.27E-08-2.7E-9+ddw_rhrpo_rf tref =25.0          rsh = 963+drsh_rhrpo_rf+rshmis
+ rjc1a = 8.89E-05     rjc1b = -4.49E-09
+ rjc2a = -2.53E-09    rjc2b = -6.64E-14
+ rint0 = 2.08E-4      rint1 = 0
+ rinttc1 = -6.46E-04  rinttc2 = -1.12E-06
+ rintjc1a = 0.365     rintjc1b = 1.45E+3
+ rintjc2a = -13.1689  rintjc2b = -1.52E+7
+weff     = w*0.9-2*dw       leff   = l*0.9
+tcoef     = 1.0+(devt-25.0)*(rtc1+rtc2*(devt-25.0))
+rintvc1 = rintjc1a + rintjc1b * weff  rintvc2 = rintjc2a + rintjc2b * weff
+rinttcoef = 1.0+(devt-25.0)*(rinttc1+rinttc2*(devt-25.0))
+rvc1 = rjc1a + rjc1b / (l*0.9)           rvc2 = (rjc2a + rjc2b / (l*0.9)) / (l*0.9)
//
+Ls_rf	  = max((4.246819E-02*pwr(w*1e6,-9.933603E-01)+0.00426)*pwr(l*1e6,(4.312050E-01*pwr(w*1e6,-5.234278E-01)+2.61))*0.9*1e-9, 1e-13)
+Cf_rf	  = max(((8.2020E-04*pwr(w*1e6,1.9584)+0.022)*l*1e6+0.16284)*(9.0016*pwr(l*1e6,-0.5239))*1e-15,1e-18)
+Rs2_rf	  = max(1445.2*pwr(l/w,2.5309),1e-3)
+Rsub_rf  = max((210.2*(l/w)-127.15)*(1.01-0.0059*exp(0.0659*l/w)), 1e-3)
+Csub_rf  = max((0.01*w*l*1e12+1.21)*(0.6274*exp(0.0077*l*1e6))*1e-15,1e-18)
+Cox_rf   = max((0.0512*w*l*1e12-0.5)*1.629*pwr(w*1e6,-0.2921)*1e-15, 1e-18)
//
ls_rf (1 port2)    inductor    l=Ls_rf 
cf_rf (port1 1)    capacitor   c=Cf_rf
//Rinta_rf (port1 na port1 na) absrint_rf_hdl wr=w rtemp=devt etch=dw rsh0=rint0 tc1=rinttc1 tc2=rinttc2 jc1a=rintjc1a jc1b=rintjc1b jc2a=rintjc2a jc2b=rintjc2b tnom=tref rminvcoef=0.5 rmaxvcoef=1.5
//rs_rf (na nb na nb) polyres_rf_hdl lr=l wr=w rtemp=devt etch=dw tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rminvcoef=0.5 rmaxvcoef=1.5
//Rintb_rf (nb 1 nb 1) absrint_rf_hdl wr=w rtemp=devt etch=dw rsh0=rint0 tc1=rinttc1 tc2=rinttc2 jc1a=rintjc1a jc1b=rintjc1b jc2a=rintjc2a jc2b=rintjc2b tnom=tref rminvcoef=0.5 rmaxvcoef=1.5
Rinta_rf (port1 na) bsource     r=(rint0/weff+rint1/(weff*weff))*rinttcoef*max(min(1.0+rintvc1*abs(v(port1,na))+rintvc2*v(port1,na)*v(port1,na),1.5),0.5)
rs_rf    (na nb) bsource     r=rsh*(l*0.9)/weff*tcoef*max(min(1.0+rvc1*abs(v(na,nb))+rvc2*v(na,nb)*v(na,nb),1.5),0.5)
Rintb_rf (nb 1) bsource     r=(rint0/weff+rint1/(weff*weff))*rinttcoef*max(min(1.0+rintvc1*abs(v(nb,1))+rintvc2*v(nb,1)*v(nb,1),1.5),0.5)
rs2_rf (1 port2)   resistor    r=Rs2_rf
cf2_rf (port1 4)   capacitor   c=0.1*Cf_rf
rs3_rf (4 port2)   resistor    r=10*Rs2_rf
rsub1_rf (2 0)     resistor    r=Rsub_rf
csub1_rf (2 0)     capacitor   c=Csub_rf
cox1_rf (port1 2)  capacitor   c=Cox_rf
rsub2_rf (3 0)     resistor    r=Rsub_rf
csub2_rf (3 0)     capacitor   c=Csub_rf
cox2_rf (port2 3)  capacitor   c=Cox_rf 
ends rhrpo_ckt_rf
//******************************************************************
//*        non-silicide HR poly resistance (three terminal)        *
//******************************************************************
subckt rhrpo_ckt_rf_3t (port1 port2 B)
parameters l=0 w=0 mismod_res_rf=0
+devt=temp
//*****mismatch parameters*****
+rshmis = arsh*geo_fac*sigma_mis_r_rf*mismod_res_rf
+geo_fac = 1/sqrt(weff*leff)
+arsh = 1.55E-05
//
+ rtc1 = -6.77E-04 rtc2 = 2.08E-06
+ dw = 2.27E-08-2.7E-9+ddw_rhrpo_rf tref =25.0          rsh = 963+drsh_rhrpo_rf+rshmis
+ rjc1a = 8.89E-05     rjc1b = -4.49E-09
+ rjc2a = -2.53E-09    rjc2b = -6.64E-14
+ rint0 = 2.08E-4      rint1 = 0
+ rinttc1 = -6.46E-04  rinttc2 = -1.12E-06
+ rintjc1a = 0.365     rintjc1b = 1.45E+3
+ rintjc2a = -13.1689  rintjc2b = -1.52E+7
+weff     = w*0.9-2*dw       leff   = l*0.9
+tcoef     = 1.0+(devt-25.0)*(rtc1+rtc2*(devt-25.0))
+rintvc1 = rintjc1a + rintjc1b * weff  rintvc2 = rintjc2a + rintjc2b * weff
+rinttcoef = 1.0+(devt-25.0)*(rinttc1+rinttc2*(devt-25.0))
+rvc1 = rjc1a + rjc1b / (l*0.9)           rvc2 = (rjc2a + rjc2b / (l*0.9)) / (l*0.9)
//
+Ls_rf	  = max((4.246819E-02*pwr(w*1e6,-9.933603E-01)+0.00426)*pwr(l*1e6,(4.312050E-01*pwr(w*1e6,-5.234278E-01)+2.61))*0.9*1e-9, 1e-13)
+Cf_rf	  = max(((8.2020E-04*pwr(w*1e6,1.9584)+0.022)*l*1e6+0.16284)*(9.0016*pwr(l*1e6,-0.5239))*1e-15,1e-18)
+Rs2_rf	  = max(1445.2*pwr(l/w,2.5309),1e-3)
+Rsub_rf  = max((210.2*(l/w)-127.15)*(1.01-0.0059*exp(0.0659*l/w)), 1e-3)
+Csub_rf  = max((0.01*w*l*1e12+1.21)*(0.6274*exp(0.0077*l*1e6))*1e-15,1e-18)
+Cox_rf   = max((0.0512*w*l*1e12-0.5)*1.629*pwr(w*1e6,-0.2921)*1e-15, 1e-18)
//
ls_rf (1 port2)    inductor    l=Ls_rf 
cf_rf (port1 1)    capacitor   c=Cf_rf
//Rinta_rf (port1 na port1 na) absrint_rf_hdl wr=w rtemp=devt etch=dw rsh0=rint0 tc1=rinttc1 tc2=rinttc2 jc1a=rintjc1a jc1b=rintjc1b jc2a=rintjc2a jc2b=rintjc2b tnom=tref rminvcoef=0.5 rmaxvcoef=1.5
//rs_rf (na nb na nb) polyres_rf_hdl lr=l wr=w rtemp=devt etch=dw tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rminvcoef=0.5 rmaxvcoef=1.5
//Rintb_rf (nb 1 nb 1) absrint_rf_hdl wr=w rtemp=devt etch=dw rsh0=rint0 tc1=rinttc1 tc2=rinttc2 jc1a=rintjc1a jc1b=rintjc1b jc2a=rintjc2a jc2b=rintjc2b tnom=tref rminvcoef=0.5 rmaxvcoef=1.5
Rinta_rf (port1 na) bsource     r=(rint0/weff+rint1/(weff*weff))*rinttcoef*max(min(1.0+rintvc1*abs(v(port1,na))+rintvc2*v(port1,na)*v(port1,na),1.5),0.5)
rs_rf    (na nb) bsource     r=rsh*(l*0.9)/weff*tcoef*max(min(1.0+rvc1*abs(v(na,nb))+rvc2*v(na,nb)*v(na,nb),1.5),0.5)
Rintb_rf (nb 1) bsource     r=(rint0/weff+rint1/(weff*weff))*rinttcoef*max(min(1.0+rintvc1*abs(v(nb,1))+rintvc2*v(nb,1)*v(nb,1),1.5),0.5)
rs2_rf (1 port2)   resistor    r=Rs2_rf
cf2_rf (port1 4)   capacitor   c=0.1*Cf_rf
rs3_rf (4 port2)   resistor    r=10*Rs2_rf
rsub1_rf (2 B)     resistor    r=Rsub_rf
csub1_rf (2 B)     capacitor   c=Csub_rf
cox1_rf (port1 2)  capacitor   c=Cox_rf
rsub2_rf (3 B)     resistor    r=Rsub_rf
csub2_rf (3 B)     capacitor   c=Csub_rf
cox2_rf (port2 3)  capacitor   c=Cox_rf 
ends rhrpo_ckt_rf_3t
//
