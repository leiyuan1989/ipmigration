
****Sub-Circuit for SDGRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNHSV1 CK D Q QN RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM52 QN ps VSS VPW N12LL W=290.00n L=60.00n
MM3 m c ps VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=410.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=270.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=410.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM53 QN ps VDD VNW P12LL W=440.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=530.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=410.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=530.00n L=60.00n
MM1 m pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS SDGRNHSV1
****Sub-Circuit for SDGRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNHSV2 CK D Q QN RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM52 QN ps VSS VPW N12LL W=430.00n L=60.00n
MM3 m c ps VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=410.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=340.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=270.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=410.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM53 QN ps VDD VNW P12LL W=650.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=530.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=410.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=530.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRNHSV2
****Sub-Circuit for SDGRNHSV4, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT SDGRNHSV4 CK D Q QN RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM52 QN ps VSS VPW N12LL W=860.00n L=60.00n
MM3 m c ps VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=360.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=410.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=270.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=410.00n L=60.00n
MM0 m pm VSS VPW N12LL W=390.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM53 QN ps VDD VNW P12LL W=1.3u L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=540.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=530.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=410.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=530.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRNHSV4
****Sub-Circuit for SDGRNQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNQHSV1 CK D Q RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM3 m c ps VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=380.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=250.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=380.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=530.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=500.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=380.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS SDGRNQHSV1
****Sub-Circuit for SDGRNQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNQHSV2 CK D Q RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM3 m c ps VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=330.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=330.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=380.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=340.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=250.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=380.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=500.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=380.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRNQHSV2
****Sub-Circuit for SDGRNQHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SDGRNQHSV4 CK D Q RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM3 m c ps VPW N12LL W=370.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=360.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=380.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=250.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=380.00n L=60.00n
MM0 m pm VSS VPW N12LL W=390.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=540.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=500.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=360.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=580.00n L=60.00n
.ENDS SDGRNQHSV4
****Sub-Circuit for SDGRSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRSNHSV1 CK D Q QN RN SE SI SN VDD VSS
MM45 net0370 SE net201 VPW N12LL W=300.00n L=60.00n
MM46 net201 SI VSS VPW N12LL W=300.00n L=60.00n
MM47 net0172 RN VSS VPW N12LL W=390.00n L=60.00n
MM48 net0370 SEN net213 VPW N12LL W=340.00n L=60.00n
MM49 net213 D net205 VPW N12LL W=390.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN OS VSS VPW N12LL W=290.00n L=60.00n
MM62 OS c net181 VPW N12LL W=260.00n L=60.00n
MM63 net181 S VSS VPW N12LL W=260.00n L=60.00n
MM61 M cn net193 VPW N12LL W=300.00n L=60.00n
MM58 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM70 net205 SN net0172 VPW N12LL W=390.00n L=60.00n
MM60 net193 net0370 VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=230.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=230.00n L=60.00n
MM24 net172 cn OS VPW N12LL W=200.00n L=60.00n
MM23 VSS NET64 net172 VPW N12LL W=200.00n L=60.00n
MM69 net213 SNN net0172 VPW N12LL W=300.00n L=60.00n
MM19 Q NET64 VSS VPW N12LL W=290.00n L=60.00n
MM17 NET64 OS VSS VPW N12LL W=260.00n L=60.00n
MM12 net240 c M VPW N12LL W=200.00n L=60.00n
MM11 VSS S net240 VPW N12LL W=200.00n L=60.00n
MM0 S M VSS VPW N12LL W=300.00n L=60.00n
MM66 net0418 SNN net296 VNW P12LL W=590.00n L=60.00n
MM50 net288 SI VDD VNW P12LL W=420.00n L=60.00n
MM51 net0370 SEN net288 VNW P12LL W=420.00n L=60.00n
MM52 net296 D VDD VNW P12LL W=590.00n L=60.00n
MM53 net0370 SE net0418 VNW P12LL W=590.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=450.00n L=60.00n
MM40 QN OS VDD VNW P12LL W=440.00n L=60.00n
MM64 net268 S VDD VNW P12LL W=390.00n L=60.00n
MM65 OS cn net268 VNW P12LL W=390.00n L=60.00n
MM67 net0418 RN VDD VNW P12LL W=450.00n L=60.00n
MM59 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=360.00n L=60.00n
MM26 VDD NET64 net253 VNW P12LL W=300.00n L=60.00n
MM25 net253 c OS VNW P12LL W=300.00n L=60.00n
MM20 Q NET64 VDD VNW P12LL W=440.00n L=60.00n
MM18 NET64 OS VDD VNW P12LL W=390.00n L=60.00n
MM14 net313 cn M VNW P12LL W=300.00n L=60.00n
MM13 VDD S net313 VNW P12LL W=300.00n L=60.00n
MM55 net280 net0370 VDD VNW P12LL W=450.00n L=60.00n
MM56 M c net280 VNW P12LL W=450.00n L=60.00n
MM1 S M VDD VNW P12LL W=450.00n L=60.00n
.ENDS SDGRSNHSV1
****Sub-Circuit for SDGRSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRSNHSV2 CK D Q QN RN SE SI SN VDD VSS
MM45 net0370 SE net201 VPW N12LL W=270.00n L=60.00n
MM46 net201 SI VSS VPW N12LL W=270.00n L=60.00n
MM47 net0172 RN VSS VPW N12LL W=350.00n L=60.00n
MM48 net0370 SEN net213 VPW N12LL W=350.00n L=60.00n
MM49 net213 D net205 VPW N12LL W=350.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=290.00n L=60.00n
MM39 QN OS VSS VPW N12LL W=430.00n L=60.00n
MM62 OS c net181 VPW N12LL W=400.00n L=60.00n
MM63 net181 S VSS VPW N12LL W=400.00n L=60.00n
MM61 M cn net193 VPW N12LL W=260.00n L=60.00n
MM58 SEN SE VSS VPW N12LL W=290.00n L=60.00n
MM70 net205 SN net0172 VPW N12LL W=350.00n L=60.00n
MM60 net193 net0370 VSS VPW N12LL W=260.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net172 cn OS VPW N12LL W=200.00n L=60.00n
MM23 VSS NET64 net172 VPW N12LL W=200.00n L=60.00n
MM69 net213 SNN net0172 VPW N12LL W=300.00n L=60.00n
MM19 Q NET64 VSS VPW N12LL W=430.00n L=60.00n
MM17 NET64 OS VSS VPW N12LL W=300.00n L=60.00n
MM12 net240 c M VPW N12LL W=200.00n L=60.00n
MM11 VSS S net240 VPW N12LL W=200.00n L=60.00n
MM0 S M VSS VPW N12LL W=360.00n L=60.00n
MM66 net0418 SNN net296 VNW P12LL W=590.00n L=60.00n
MM50 net288 SI VDD VNW P12LL W=410.00n L=60.00n
MM51 net0370 SEN net288 VNW P12LL W=410.00n L=60.00n
MM52 net296 D VDD VNW P12LL W=590.00n L=60.00n
MM53 net0370 SE net0418 VNW P12LL W=590.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=440.00n L=60.00n
MM40 QN OS VDD VNW P12LL W=650.00n L=60.00n
MM64 net268 S VDD VNW P12LL W=480.00n L=60.00n
MM65 OS cn net268 VNW P12LL W=480.00n L=60.00n
MM67 net0418 RN VDD VNW P12LL W=400.00n L=60.00n
MM59 SEN SE VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD NET64 net253 VNW P12LL W=300.00n L=60.00n
MM25 net253 c OS VNW P12LL W=300.00n L=60.00n
MM20 Q NET64 VDD VNW P12LL W=650.00n L=60.00n
MM18 NET64 OS VDD VNW P12LL W=450.00n L=60.00n
MM14 net313 cn M VNW P12LL W=300.00n L=60.00n
MM13 VDD S net313 VNW P12LL W=300.00n L=60.00n
MM55 net280 net0370 VDD VNW P12LL W=390.00n L=60.00n
MM56 M c net280 VNW P12LL W=390.00n L=60.00n
MM1 S M VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRSNHSV2
****Sub-Circuit for SDGRSNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRSNHSV4 CK D Q QN RN SE SI SN VDD VSS
MM45 net0370 SE net201 VPW N12LL W=300.00n L=60.00n
MM46 net201 SI VSS VPW N12LL W=300.00n L=60.00n
MM47 net0172 RN VSS VPW N12LL W=350.00n L=60.00n
MM48 net0370 SEN net213 VPW N12LL W=350.00n L=60.00n
MM49 net213 D net205 VPW N12LL W=350.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=290.00n L=60.00n
MM39 QN OS VSS VPW N12LL W=860.00n L=60.00n
MM62 OS c net181 VPW N12LL W=450.00n L=60.00n
MM63 net181 S VSS VPW N12LL W=450.00n L=60.00n
MM61 M cn net193 VPW N12LL W=260.00n L=60.00n
MM58 SEN SE VSS VPW N12LL W=290.00n L=60.00n
MM70 net205 SN net0172 VPW N12LL W=350.00n L=60.00n
MM60 net193 net0370 VSS VPW N12LL W=260.00n L=60.00n
MM30 c cn VSS VPW N12LL W=260.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net172 cn OS VPW N12LL W=200.00n L=60.00n
MM23 VSS NET64 net172 VPW N12LL W=200.00n L=60.00n
MM69 net213 SNN net0172 VPW N12LL W=300.00n L=60.00n
MM19 Q NET64 VSS VPW N12LL W=860.00n L=60.00n
MM17 NET64 OS VSS VPW N12LL W=360.00n L=60.00n
MM12 net240 c M VPW N12LL W=200.00n L=60.00n
MM11 VSS S net240 VPW N12LL W=200.00n L=60.00n
MM0 S M VSS VPW N12LL W=360.00n L=60.00n
MM66 net0418 SNN net296 VNW P12LL W=590.00n L=60.00n
MM50 net288 SI VDD VNW P12LL W=450.00n L=60.00n
MM51 net0370 SEN net288 VNW P12LL W=450.00n L=60.00n
MM52 net296 D VDD VNW P12LL W=590.00n L=60.00n
MM53 net0370 SE net0418 VNW P12LL W=590.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=440.00n L=60.00n
MM40 QN OS VDD VNW P12LL W=1.3u L=60.00n
MM64 net268 S VDD VNW P12LL W=570.00n L=60.00n
MM65 OS cn net268 VNW P12LL W=570.00n L=60.00n
MM67 net0418 RN VDD VNW P12LL W=400.00n L=60.00n
MM59 SEN SE VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=390.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD NET64 net253 VNW P12LL W=300.00n L=60.00n
MM25 net253 c OS VNW P12LL W=300.00n L=60.00n
MM20 Q NET64 VDD VNW P12LL W=1.3u L=60.00n
MM18 NET64 OS VDD VNW P12LL W=540.00n L=60.00n
MM14 net313 cn M VNW P12LL W=300.00n L=60.00n
MM13 VDD S net313 VNW P12LL W=300.00n L=60.00n
MM55 net280 net0370 VDD VNW P12LL W=390.00n L=60.00n
MM56 M c net280 VNW P12LL W=390.00n L=60.00n
MM1 S M VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRSNHSV4
****Sub-Circuit for SDGSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGSNHSV1 CK D Q QN SE SI SN VDD VSS
MM39 QN PS VSS VPW N12LL W=290.00n L=60.00n
MM45 N74 SE net0128 VPW N12LL W=200.00n L=60.00n
MM46 net0128 SI VSS VPW N12LL W=200.00n L=60.00n
MM48 N74 cn PM VPW N12LL W=270.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=200.00n L=60.00n
MM52 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM3 M c PS VPW N12LL W=270.00n L=60.00n
MM42 net69 SNN VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=250.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn PS VPW N12LL W=200.00n L=60.00n
MM23 VSS S net48 VPW N12LL W=200.00n L=60.00n
MM19 Q S VSS VPW N12LL W=290.00n L=60.00n
MM17 S PS VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c PM VPW N12LL W=200.00n L=60.00n
MM11 VSS M net52 VPW N12LL W=200.00n L=60.00n
MM9 N74 SEN net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=250.00n L=60.00n
MM0 M PM VSS VPW N12LL W=270.00n L=60.00n
MM41 net_0231 SNN VDD VNW P12LL W=400.00n L=60.00n
MM40 QN PS VDD VNW P12LL W=440.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=300.00n L=60.00n
MM50 net0207 SI VDD VNW P12LL W=300.00n L=60.00n
MM51 N74 SEN net0207 VNW P12LL W=300.00n L=60.00n
MM54 N74 c PM VNW P12LL W=400.00n L=60.00n
MM4 M cn PS VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=380.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD S net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c PS VNW P12LL W=300.00n L=60.00n
MM20 Q S VDD VNW P12LL W=440.00n L=60.00n
MM18 S PS VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn PM VNW P12LL W=300.00n L=60.00n
MM13 VDD M net117 VNW P12LL W=300.00n L=60.00n
MM10 N74 SE net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=400.00n L=60.00n
MM56 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM1 M PM VDD VNW P12LL W=400.00n L=60.00n
.ENDS SDGSNHSV1
****Sub-Circuit for SDGSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGSNHSV2 CK D Q QN SE SI SN VDD VSS
MM39 QN PS VSS VPW N12LL W=430.00n L=60.00n
MM45 N74 SE net0128 VPW N12LL W=200.00n L=60.00n
MM46 net0128 SI VSS VPW N12LL W=200.00n L=60.00n
MM48 N74 cn PM VPW N12LL W=360.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=200.00n L=60.00n
MM52 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM3 M c PS VPW N12LL W=390.00n L=60.00n
MM42 net69 SNN VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=380.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn PS VPW N12LL W=200.00n L=60.00n
MM23 VSS S net48 VPW N12LL W=200.00n L=60.00n
MM19 Q S VSS VPW N12LL W=430.00n L=60.00n
MM17 S PS VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c PM VPW N12LL W=200.00n L=60.00n
MM11 VSS M net52 VPW N12LL W=200.00n L=60.00n
MM9 N74 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 M PM VSS VPW N12LL W=390.00n L=60.00n
MM41 net_0231 SNN VDD VNW P12LL W=600.0n L=60.00n
MM40 QN PS VDD VNW P12LL W=650.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=300.00n L=60.00n
MM50 net0207 SI VDD VNW P12LL W=300.00n L=60.00n
MM51 N74 SEN net0207 VNW P12LL W=300.00n L=60.00n
MM54 N74 c PM VNW P12LL W=540.00n L=60.00n
MM4 M cn PS VNW P12LL W=580.00n L=60.00n
MM29 c cn VDD VNW P12LL W=570.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD S net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c PS VNW P12LL W=300.00n L=60.00n
MM20 Q S VDD VNW P12LL W=650.00n L=60.00n
MM18 S PS VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn PM VNW P12LL W=300.00n L=60.00n
MM13 VDD M net117 VNW P12LL W=300.00n L=60.00n
MM10 N74 SE net128 VNW P12LL W=600.0n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=600.0n L=60.00n
MM56 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM1 M PM VDD VNW P12LL W=580.00n L=60.00n
.ENDS SDGSNHSV2
****Sub-Circuit for SDGSNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGSNHSV4 CK D Q QN SE SI SN VDD VSS
MM39 QN PS VSS VPW N12LL W=860.00n L=60.00n
MM45 N74 SE net0128 VPW N12LL W=200.00n L=60.00n
MM46 net0128 SI VSS VPW N12LL W=200.00n L=60.00n
MM48 N74 cn PM VPW N12LL W=400.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=200.00n L=60.00n
MM52 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM3 M c PS VPW N12LL W=430.00n L=60.00n
MM42 net69 SNN VSS VPW N12LL W=250.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn PS VPW N12LL W=200.00n L=60.00n
MM23 VSS S net48 VPW N12LL W=200.00n L=60.00n
MM19 Q S VSS VPW N12LL W=860.00n L=60.00n
MM17 S PS VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c PM VPW N12LL W=200.00n L=60.00n
MM11 VSS M net52 VPW N12LL W=200.00n L=60.00n
MM9 N74 SEN net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 M PM VSS VPW N12LL W=430.00n L=60.00n
MM41 net_0231 SNN VDD VNW P12LL W=650.00n L=60.00n
MM40 QN PS VDD VNW P12LL W=1.3u L=60.00n
MM44 SNN SN VDD VNW P12LL W=300.00n L=60.00n
MM50 net0207 SI VDD VNW P12LL W=300.00n L=60.00n
MM51 N74 SEN net0207 VNW P12LL W=300.00n L=60.00n
MM54 N74 c PM VNW P12LL W=600.0n L=60.00n
MM4 M cn PS VNW P12LL W=650.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD S net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c PS VNW P12LL W=300.00n L=60.00n
MM20 Q S VDD VNW P12LL W=1.3u L=60.00n
MM18 S PS VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn PM VNW P12LL W=300.00n L=60.00n
MM13 VDD M net117 VNW P12LL W=300.00n L=60.00n
MM10 N74 SE net128 VNW P12LL W=650.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=650.00n L=60.00n
MM56 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM1 M PM VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDGSNHSV4
****Sub-Circuit for SDHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDHSV1 CK D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=290.00n L=60.00n
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=280.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=280.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=290.00n L=60.00n
MM53 QN s VDD VNW P12LL W=440.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=300.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=300.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDHSV1
****Sub-Circuit for SDHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDHSV2 CK D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=430.00n L=60.00n
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=400.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=400.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM53 QN s VDD VNW P12LL W=650.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDHSV2
****Sub-Circuit for SDHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDHSV4 CK D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=860.00n L=60.00n
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=420.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=300.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=300.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM53 QN s VDD VNW P12LL W=1.3u L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=520.0n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=520.0n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.0n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDHSV4
****Sub-Circuit for SDQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDQHSV1 CK D Q SE SI VDD VSS
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=280.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=280.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=290.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=300.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=300.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDQHSV1
****Sub-Circuit for SDQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDQHSV2 CK D Q SE SI VDD VSS
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=400.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=400.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDQHSV2
****Sub-Circuit for SDQHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SDQHSV4 CK D Q SE SI VDD VSS
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=430.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=300.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=300.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=490.0n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=490.0n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.0n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDQHSV4
****Sub-Circuit for SDRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNHSV1 CK D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=290.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=290.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=290.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=290.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=440.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=330.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=330.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=330.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDRNHSV1
****Sub-Circuit for SDRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNHSV2 CK D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=430.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=320.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=320.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=650.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=350.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=350.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=350.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNHSV2
****Sub-Circuit for SDRNHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SDRNHSV4 CK D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=430.00n L=60.00n m=2
MM45 net_0137 sen net_0133 VPW N12LL W=430.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=400.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=300.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=300.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=650.00n L=60.00n m=2
MM47 net_0137 SE net_0212 VNW P12LL W=500n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=450.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=500n L=60.00n
MM8 net128 SI VDD VNW P12LL W=500n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNHSV4
****Sub-Circuit for SDRNQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNQHSV1 CK D Q RDN SE SI VDD VSS
MM45 net_0137 sen net_0133 VPW N12LL W=290.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=290.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=290.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=330.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=330.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=330.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDRNQHSV1
****Sub-Circuit for SDRNQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNQHSV2 CK D Q RDN SE SI VDD VSS
MM45 net_0137 sen net_0133 VPW N12LL W=320.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=320.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=350.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=350.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=350.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNQHSV2
****Sub-Circuit for SDRNQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNQHSV4 CK D Q RDN SE SI VDD VSS
MM45 net_0137 sen net_0133 VPW N12LL W=430.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=400.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=300.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=300.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=500n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=450.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=500n L=60.00n
MM8 net128 SI VDD VNW P12LL W=500n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNQHSV4
****Sub-Circuit for SDRSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRSNHSV1 CK D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=250.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=290.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=200.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=260.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=260.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=260.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=260.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=280.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=330.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=420.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=380.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=330.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=330.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=330.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=440.00n L=60.00n
.ENDS SDRSNHSV1
****Sub-Circuit for SDRSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRSNHSV2 CK D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=280.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=250.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=360.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=390.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=200.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=220.00n L=60.00n
MM40 net43 R L VPW N12LL W=280.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=220.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=220.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=220.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=380.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=300.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=300.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=600.00n L=60.00n
.ENDS SDRSNHSV2
****Sub-Circuit for SDRSNHSV4, Mon May 30 16:10:14 CST 2011****
.SUBCKT SDRSNHSV4 CK D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=280.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=250.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=320.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=430.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=400.00n L=60.00n
MM40 net43 R L VPW N12LL W=280.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=400.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=400.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=500.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM57 net_0140 c net_0139 VNW P12LL W=580.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=600.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=520.00n L=60.00n
MM29 c cn VDD VNW P12LL W=620.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=380.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=500.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=500.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=500.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=650.00n L=60.00n
.ENDS SDRSNHSV4
****Sub-Circuit for SDSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDSNHSV1 CK D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=300.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=300.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=200.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=400.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=400.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=300.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=450.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=450.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=400.00n L=60.00n
.ENDS SDSNHSV1
****Sub-Circuit for SDSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDSNHSV2 CK D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=300.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=300.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=200.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=420.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=420.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=300.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=450.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=450.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=390.00n L=60.00n
.ENDS SDSNHSV2
****Sub-Circuit for SDSNHSV4, Mon May 30 17:13:17 CST 2011****
.SUBCKT SDSNHSV4 CK D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=300.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=300.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=200.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=360.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=300.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=450.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=450.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM38 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=625.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=480.00n L=60.00n
.ENDS SDSNHSV4
****Sub-Circuit for SDXHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDXHSV1 CK DA DB Q QN SA SE SI VDD VSS
MM5 net41 SB net_0171 VPW N12LL W=240.00n L=60.00n
MM49 net39 DA VSS VPW N12LL W=350.00n L=60.00n
MM48 net39 SA net_0171 VPW N12LL W=240.00n L=60.00n
MM37 SEN SE VSS VPW N12LL W=240.00n L=60.00n
MM41 net41 DB VSS VPW N12LL W=350.00n L=60.00n
MM31 SB SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=350.00n L=60.00n
MM19 QN s VSS VPW N12LL W=350.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM7 m c net43 VPW N12LL W=350.00n L=60.00n
MM12 net52 c net_0157 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM46 net_0169 SE VSS VPW N12LL W=240.00n L=60.00n
MM45 net_0153 sin net_0169 VPW N12LL W=240.00n L=60.00n
MM43 net_0161 SEN VSS VPW N12LL W=300.00n L=60.00n
MM9 net_0157 cn net_0153 VPW N12LL W=300.00n L=60.00n
MM42 net_0153 net_0171 net_0161 VPW N12LL W=300.00n L=60.00n
MM6 sin SI VSS VPW N12LL W=350.00n L=60.00n
MM0 m net_0157 VSS VPW N12LL W=350.00n L=60.00n
MM52 net39 DA VDD VNW P12LL W=440.0n L=60.00n
MM53 sin SI VDD VNW P12LL W=440.0n L=60.00n
MM54 net41 SA net_0171 VNW P12LL W=300.0n L=60.00n
MM55 net41 DB VDD VNW P12LL W=440.0n L=60.00n
MM56 net39 SB net_0171 VNW P12LL W=300.0n L=60.00n
MM38 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM4 m cn net43 VNW P12LL W=440.0n L=60.00n
MM44 net_0236 SE VDD VNW P12LL W=450.00n L=60.00n
MM32 SB SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM20 QN s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM47 net_0233 net_0171 net_0236 VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0157 VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM51 net_0233 sin net_0252 VNW P12LL W=300.00n L=60.00n
MM50 net_0252 SEN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0157 c net_0233 VNW P12LL W=450.00n L=60.00n
MM1 m net_0157 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDXHSV1
****Sub-Circuit for SDXHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDXHSV2 CK DA DB Q QN SA SE SI VDD VSS
MM8 sin SI VSS VPW N12LL W=350.00n L=60.00n
MM41 net41 DB VSS VPW N12LL W=430.00n L=60.00n
MM37 SEN SE VSS VPW N12LL W=240.00n L=60.00n
MM31 SB SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM19 QN s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM2 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0157 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM46 net_0169 SE VSS VPW N12LL W=240.00n L=60.00n
MM45 net_0153 sin net_0169 VPW N12LL W=240.00n L=60.00n
MM43 net_0161 SEN VSS VPW N12LL W=350.00n L=60.00n
MM9 net_0157 cn net_0153 VPW N12LL W=350.00n L=60.00n
MM42 net_0153 net_0152 net_0161 VPW N12LL W=350.00n L=60.00n
MM48 net39 SA net_0152 VPW N12LL W=240.00n L=60.00n
MM5 net41 SB net_0152 VPW N12LL W=240.00n L=60.00n
MM49 net39 DA VSS VPW N12LL W=430.00n L=60.00n
MM0 m net_0157 VSS VPW N12LL W=430.00n L=60.00n
MM38 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM53 sin SI VDD VNW P12LL W=440.0n L=60.00n
MM44 net_0236 SE VDD VNW P12LL W=440.00n L=60.00n
MM32 SB SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=550.00n L=60.00n
MM20 QN s VDD VNW P12LL W=550.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM7 m cn net43 VNW P12LL W=540.00n L=60.00n
MM47 net_0233 net_0152 net_0236 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0157 VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM51 net_0233 sin net_0252 VNW P12LL W=300.00n L=60.00n
MM50 net_0252 SEN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0157 c net_0233 VNW P12LL W=440.00n L=60.00n
MM56 net39 SB net_0152 VNW P12LL W=300.0n L=60.00n
MM54 net41 SA net_0152 VNW P12LL W=300.0n L=60.00n
MM55 net41 DB VDD VNW P12LL W=550.0n L=60.00n
MM52 net39 DA VDD VNW P12LL W=550.0n L=60.00n
MM1 m net_0157 VDD VNW P12LL W=550.00n L=60.00n
.ENDS SDXHSV2
****Sub-Circuit for SDXHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDXHSV4 CK DA DB Q QN SA SE SI VDD VSS
MM8 sin SI VSS VPW N12LL W=350.00n L=60.00n
MM41 net41 DB VSS VPW N12LL W=430.00n L=60.00n
MM37 SEN SE VSS VPW N12LL W=240.00n L=60.00n
MM31 SB SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM19 QN s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM2 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0157 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM46 net_0169 SE VSS VPW N12LL W=240.00n L=60.00n
MM45 net_0153 sin net_0169 VPW N12LL W=240.00n L=60.00n
MM43 net_0161 SEN VSS VPW N12LL W=350.00n L=60.00n
MM9 net_0157 cn net_0153 VPW N12LL W=350.00n L=60.00n
MM42 net_0153 net_0152 net_0161 VPW N12LL W=350.00n L=60.00n
MM49 net39 DA VSS VPW N12LL W=430.00n L=60.00n
MM5 net41 SB net_0152 VPW N12LL W=240.00n L=60.00n
MM48 net39 SA net_0152 VPW N12LL W=240.00n L=60.00n
MM0 m net_0157 VSS VPW N12LL W=430.00n L=60.00n
MM38 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0236 SE VDD VNW P12LL W=440.00n L=60.00n
MM56 net39 SB net_0152 VNW P12LL W=300.0n L=60.00n
MM54 net41 SA net_0152 VNW P12LL W=300.0n L=60.00n
MM52 net39 DA VDD VNW P12LL W=550.0n L=60.00n
MM55 net41 DB VDD VNW P12LL W=550.0n L=60.00n
MM32 SB SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.1u L=60.00n
MM20 QN s VDD VNW P12LL W=1.1u L=60.00n
MM18 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM53 sin SI VDD VNW P12LL W=440.0n L=60.00n
MM7 m cn net43 VNW P12LL W=540.00n L=60.00n
MM47 net_0233 net_0152 net_0236 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0157 VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM51 net_0233 sin net_0252 VNW P12LL W=300.00n L=60.00n
MM50 net_0252 SEN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0157 c net_0233 VNW P12LL W=440.00n L=60.00n
MM1 m net_0157 VDD VNW P12LL W=550.00n L=60.00n
.ENDS SDXHSV4
****Sub-Circuit for SEDGRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNHSV1 CK D E Q QN RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM64 QN s VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=290.00n L=60.00n
MM17 sp s VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM65 QN s VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=440.00n L=60.00n
MM18 sp s VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNHSV1
****Sub-Circuit for SEDGRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNHSV2 CK D E Q QN RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM64 QN s VSS VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=430.00n L=60.00n
MM17 sp s VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM65 QN s VDD VNW P12LL W=650.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=650.00n L=60.00n
MM18 sp s VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNHSV2
****Sub-Circuit for SEDGRNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNHSV4 CK D E Q QN RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM64 QN s VSS VPW N12LL W=860.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=860.00n L=60.00n
MM17 sp s VSS VPW N12LL W=400.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM65 QN s VDD VNW P12LL W=1.3u L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=1.3u L=60.00n
MM18 sp s VDD VNW P12LL W=480.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNHSV4
****Sub-Circuit for SEDGRNQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNQHSV1 CK D E Q RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=290.00n L=60.00n
MM17 sp s VSS VPW N12LL W=220.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=440.00n L=60.00n
MM18 sp s VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNQHSV1
****Sub-Circuit for SEDGRNQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNQHSV2 CK D E Q RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=430.00n L=60.00n
MM17 sp s VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=650.00n L=60.00n
MM18 sp s VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNQHSV2
****Sub-Circuit for SEDGRNQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNQHSV4 CK D E Q RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=860.00n L=60.00n
MM17 sp s VSS VPW N12LL W=310.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=1.3u L=60.00n
MM18 sp s VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNQHSV4
****Sub-Circuit for SEDHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDHSV1 CK D E Q QN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=300.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=300.00n L=60.00n
MM68 QN s VSS VPW N12LL W=290.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=420.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=420.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=420.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=420.00n L=60.00n
MM0 m pm VSS VPW N12LL W=400.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=300.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=300.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM69 QN s VDD VNW P12LL W=440.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=600.00n L=60.00n
.ENDS SEDHSV1
****Sub-Circuit for SEDHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDHSV2 CK D E Q QN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 QN s VSS VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=400.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=400.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM69 QN s VDD VNW P12LL W=650.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDHSV2
****Sub-Circuit for SEDHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDHSV4 CK D E Q QN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 QN s VSS VPW N12LL W=860.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=390.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=440.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=440.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM69 QN s VDD VNW P12LL W=1.3u L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDHSV4
****Sub-Circuit for SEDQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDQHSV1 CK D E Q SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=300.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=300.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=300.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=300.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDQHSV1
****Sub-Circuit for SEDQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDQHSV2 CK D E Q SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=400.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=400.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDQHSV2
****Sub-Circuit for SEDQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDQHSV4 CK D E Q SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=420.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=420.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDQHSV4
****Sub-Circuit for SEDRNHSV1, Fri May 27 10:36:55 CST 2011****
.SUBCKT SEDRNHSV1 CK D E Q QN RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=390.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM73 QN s VSS VPW N12LL W=290.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=250.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=250.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=275.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=250.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=270.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM74 QN s VDD VNW P12LL W=440.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=355.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=390.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=390.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=380.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=400.00n L=60.00n
.ENDS SEDRNHSV1
****Sub-Circuit for SEDRNHSV2, Thu May 26 17:37:04 CST 2011****
.SUBCKT SEDRNHSV2 CK D E Q QN RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=390.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM73 QN s VSS VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=250.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=250.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=275.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM74 QN s VDD VNW P12LL W=650.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=355.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=390.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=390.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SEDRNHSV2
****Sub-Circuit for SEDRNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDRNHSV4 CK D E Q QN RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=360.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=360.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM73 QN s VSS VPW N12LL W=860.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=250.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=250.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=275.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=400.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=400.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=470.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=470.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM74 QN s VDD VNW P12LL W=1.3u L=60.00n
MM53 net0267 SE VDD VNW P12LL W=355.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=390.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=390.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=600.00n L=60.00n
.ENDS SEDRNHSV4
****Sub-Circuit for SEDRNQHSV1, Thu May 26 14:31:08 CST 2011****
.SUBCKT SEDRNQHSV1 CK D E Q RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=390.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=240.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=240.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=300.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=385.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=385.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=370.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=380.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=380.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDRNQHSV1
****Sub-Circuit for SEDRNQHSV2, Thu May 26 13:48:52 CST 2011****
.SUBCKT SEDRNQHSV2 CK D E Q RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=240.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=240.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=290.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=380.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=380.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=380.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDRNQHSV2
****Sub-Circuit for SEDRNQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDRNQHSV4 CK D E Q RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=240.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=240.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=300.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=390.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=380.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=380.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDRNQHSV4
****Sub-Circuit for SNDHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDHSV1 CKN D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=290.00n L=60.00n
MM46 net_0107 SE VSS VPW N12LL W=250.00n L=60.00n
MM45 net_0163 SI net_0107 VPW N12LL W=250.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=230.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=230.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=250.00n L=60.00n
MM30 cn c VSS VPW N12LL W=250.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=250.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=250.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=270.00n L=60.00n
MM53 QN s VDD VNW P12LL W=440.00n L=60.00n
MM51 net128 SI net_0174 VNW P12LL W=650.00n L=60.00n
MM50 net_0174 SEN VDD VNW P12LL W=650.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=380.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=650.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=650.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=650.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=400.00n L=60.00n
.ENDS SNDHSV1
****Sub-Circuit for SNDHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDHSV2 CKN D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=430.00n L=60.00n
MM46 net_0107 SE VSS VPW N12LL W=250.00n L=60.00n
MM45 net_0163 SI net_0107 VPW N12LL W=250.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=230.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=230.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=250.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=250.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=250.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=390.00n L=60.00n
MM53 QN s VDD VNW P12LL W=650.00n L=60.00n
MM51 net128 SI net_0174 VNW P12LL W=650.00n L=60.00n
MM50 net_0174 SEN VDD VNW P12LL W=650.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=650.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=650.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=650.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=580.00n L=60.00n
.ENDS SNDHSV2
****Sub-Circuit for SNDHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDHSV4 CKN D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=860.00n L=60.00n
MM46 net_0107 SE VSS VPW N12LL W=260.00n L=60.00n
MM45 net_0163 SI net_0107 VPW N12LL W=260.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=250.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=250.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=260.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=260.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=260.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM53 QN s VDD VNW P12LL W=1.3u L=60.00n
MM51 net128 SI net_0174 VNW P12LL W=650.00n L=60.00n
MM50 net_0174 SEN VDD VNW P12LL W=650.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=650.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=650.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=650.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SNDHSV4
****Sub-Circuit for SNDRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRNHSV1 CKN D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=290.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=300.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=300.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=300.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=300.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=300.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM39 s ps net_099 VPW N12LL W=360.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=360.00n L=60.00n
MM30 cn c VSS VPW N12LL W=300.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=300.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=440.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=500.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM38 s ps VDD VNW P12LL W=390.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=390.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=450.00n L=60.00n
MM29 cn c VDD VNW P12LL W=450.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=450.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=450.00n L=60.00n
.ENDS SNDRNHSV1
****Sub-Circuit for SNDRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRNHSV2 CKN D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=430.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=350.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=350.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=300.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=290.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=300.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=190.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM39 s ps net_099 VPW N12LL W=360.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=360.00n L=60.00n
MM30 cn c VSS VPW N12LL W=300.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=190.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=190.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=300.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=650.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=450.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=450.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM38 s ps VDD VNW P12LL W=390.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=390.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=445.00n L=60.00n
MM29 cn c VDD VNW P12LL W=450.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=450.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=450.00n L=60.00n
.ENDS SNDRNHSV2
****Sub-Circuit for SNDRNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRNHSV4 CKN D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=860.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=350.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=350.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=300.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=300.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=300.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM39 s ps net_099 VPW N12LL W=380.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=380.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=300.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=1.3u L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=500.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM38 s ps VDD VNW P12LL W=350.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=450.00n L=60.00n
MM29 cn c VDD VNW P12LL W=530.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn ps VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=450.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=450.00n L=60.00n
.ENDS SNDRNHSV4
****Sub-Circuit for SNDRSNHSV1, Mon May 30 19:16:43 CST 2011****
.SUBCKT SNDRSNHSV1 CKN D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=270.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=340.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=300.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=300.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=300.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=300.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=450.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=450.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=500.00n L=60.00n
MM29 cn c VDD VNW P12LL W=540.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=540.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=540.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=500.00n L=60.00n
.ENDS SNDRSNHSV1
****Sub-Circuit for SNDRSNHSV2, Mon May 30 17:13:17 CST 2011****
.SUBCKT SNDRSNHSV2 CKN D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=270.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=340.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=300.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=300.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=300.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=300.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=450.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=450.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=500.00n L=60.00n
MM29 cn c VDD VNW P12LL W=540.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=540.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=540.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=500.00n L=60.00n
.ENDS SNDRSNHSV2
****Sub-Circuit for SNDRSNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRSNHSV4 CKN D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=270.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=350.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=360.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=300.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=320.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=320.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=300.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=450.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=450.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=540.00n L=60.00n
MM29 cn c VDD VNW P12LL W=540.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=540.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=540.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=540.00n L=60.00n
.ENDS SNDRSNHSV4
****Sub-Circuit for SNDSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDSNHSV1 CKN D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=220.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=220.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=220.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=220.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=200.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=250.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=220.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=430.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=480.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=480.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=480.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=480.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=380.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=480.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=500.00n L=60.00n
.ENDS SNDSNHSV1
****Sub-Circuit for SNDSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDSNHSV2 CKN D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=220.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=220.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=220.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=220.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=250.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=220.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=430.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=480.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=480.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=480.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=480.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=480.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=500.00n L=60.00n
.ENDS SNDSNHSV2
****Sub-Circuit for SNDSNHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SNDSNHSV4 CKN D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=250.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=250.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=250.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=250.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=390.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=250.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=430.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=480.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=480.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=480.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=480.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM38 s net43 VDD VNW P12LL W=540.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=470.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=480.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=500.00n L=60.00n
.ENDS SNDSNHSV4