
******************arithmetic************************






******************INV************************

.SUBCKT INV_1 IN1 VDD VSS OUT1
PM1 VDD  IN1  OUT1 VDD pmos l=1 w=1 n=1 ro=5 co=1
NM1 VSS  IN1  OUT1 VSS nmos l=1 w=1 n=1 ro=2 co=1
.ends INV_1


.subckt INV_2 VSS Y VDD A
PM1 OUT1 IN1  VDD  VDD pmos l=1 w=1 n=1 ro=5 co=1
PM2 VDD  IN1  OUT1 VDD pmos l=1 w=1 n=1 ro=5 co=2
NM1 OUT1 IN1  VSS  VSS nmos l=1 w=1 n=1 ro=2 co=1
NM2 VSS  IN1  OUT1 VSS nmos l=1 w=1 n=1 ro=2 co=2
.ends INV_2

.subckt INV_3 VSS Y VDD A
PM1 VDD  IN1  OUT1 VDD pmos l=1 w=1 n=1 ro=5 co=1
PM2 OUT1 IN1  VDD VDD pmos l=1 w=1 n=1 ro=5 co=2
PM3 VDD  IN1  OUT1 VDD pmos l=1 w=1 n=1 ro=5 co=3
NM1 VSS  IN1  OUT1 VSS nmos l=1 w=1 n=1 ro=2 co=1
NM2 OUT1 IN1  VSS VSS nmos l=1 w=1 n=1 ro=2 co=2
NM3 VSS  IN1  OUT1 VSS nmos l=1 w=1 n=1 ro=2 co=3
.ends INV_3

.subckt INV_4 VSS Y VDD A
PM1 OUT1 IN1  VDD  VDD pmos l=1 w=1 n=1 ro=5 co=1
PM2 VDD  IN1  OUT1 VDD pmos l=1 w=1 n=1 ro=5 co=2
PM3 OUT1 IN1  VDD  VDD pmos l=1 w=1 n=1 ro=5 co=3
PM4 VDD  IN1  OUT1 VDD pmos l=1 w=1 n=1 ro=5 co=4
NM1 OUT1 IN1  VSS  VSS nmos l=1 w=1 n=1 ro=2 co=1
NM2 VSS  IN1  OUT1 VSS nmos l=1 w=1 n=1 ro=2 co=2
NM3 OUT1 IN1  VSS  VSS nmos l=1 w=1 n=1 ro=2 co=3
NM4 VSS  IN1  OUT1 VSS nmos l=1 w=1 n=1 ro=2 co=4
.ends INV_4




******************AND************************
.SUBCKT I2_AND2 IN1 IN2 VDD VSS OUT1
pmos_1 VDD  IN1  net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
nmos_1 net1 IN1  net2 VSS nmos l=1 w=1 n=1 ro=1 co=1
pmos_2 net1 IN2  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=2
nmos_2 net2 IN2  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=2
pmos_3 VDD  net1  OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=3
nmos_3 VSS  net1  OUT1  VSS nmos l=1 w=1 n=1 ro=1 co=3
.ends I2_AND2

.subckt I3_AND3 C B A VSS Y VDD

PM1 N_2 A   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD B   N_2 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_2 C   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD N_2 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 N_2  A  N_9  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_9  B  N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_10 C  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS N_2 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends I3_AND3

.subckt I3_AND12 B AN VSS VDD Y
PM1 VDD AN  N_4 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
NM1 VSS AN  N_4 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1

PM2 VDD N_4 N_2 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM3 N_2 B   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM4 VDD N_2 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM2 N_2  N_4 N_14 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM3 N_14 B   VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM4 VSS  N_2 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends I3_AND12


.subckt I3_AND13 C B AN VSS VDD Y
PM1 N_6 C   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD B   N_6 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_6 N_4 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3

PM4 N_4 AN  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 VDD N_6 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 VSS  C   N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_10 B   N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_11 N_4 N_6  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3

NM4 N_4  AN  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 VSS  N_6  Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I4_AND13



.subckt I3_AND23 C BN AN VDD Y VSS

PM1 N_4 AN VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD BN N_3 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2

PM3 N_5 N_4 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM4 VDD N_3 N_5 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 N_5 C   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6
PM6 VDD N_5 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=7


NM1 N_4 AN VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS BN N_3 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2

NM3 N_5  N_4 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM4 N_11 N_3 N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 N_12 C   VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
NM6 VSS  N_5 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=7
.ends I3_AND23

.subckt I4_AND4 VSS Y VDD D C B A
PM1 VDD A N_4 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_4 B VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD C N_4 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_4 D VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD N_4 Y VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 N_4 A N_6 VSS nmos  l=0.5u w=0.58u n=1 ro=1 co=1
NM2 N_6 B N_7 VSS nmos  l=0.5u w=0.58u n=1 ro=1 co=2
NM3 N_7 C N_8 VSS nmos  l=0.5u w=0.58u n=1 ro=1 co=3
NM4 N_8 D VSS VSS nmos  l=0.5u w=0.58u n=1 ro=1 co=4
NM5 VSS N_4 Y VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends I4_AND4



******************OR************************

.SUBCKT I2_OR02 IN1 IN2 VDD VSS OUT1
pmos_1 net1  IN1  net2 VDD pmos l=1 w=1 n=1 ro=1 co=1
nmos_1 VSS   IN1  net1 VSS nmos l=1 w=1 n=1 ro=1 co=1
pmos_2 net2  IN2  VDD  VDD pmos l=1 w=1 n=1 ro=1 co=2
nmos_2 net1  IN2  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=2
pmos_3 VDD  net1  OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=3
nmos_3 VSS  net1  OUT1  VSS nmos l=1 w=1 n=1 ro=1 co=3
.ends I2_OR02


* Top of hierarchy  cell=or03d0
.subckt I3_OR03 B A C VSS VDD Y
PM1 N_3  C   N_13 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_13 B   N_14 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_14 A   VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD  N_3 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 N_3 C   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS B   N_3 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_3 A   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS N_3 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends I3_OR03

* Top of hierarchy  cell=or04d0
.subckt I4_OR04 A B D C VDD Y VSS
PM1 N_3  D N_14 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_14 C N_15 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_15 B N_16 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_16 A VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD  N_3 Y  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 VSS D  N_3 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_3 C  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS B  N_3 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_3 A  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 VSS N_3 Y  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends I4_OR04


* Top of hierarchy  cell=or12d0
.subckt I2_OR12 B AN VDD VSS Y
PM1 N_4  AN  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  N_4 N_14 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_14 B   N_2  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD  N_2 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 N_4 AN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS N_4 N_2 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_2 B   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS N_2 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends I2_OR12

* Top of hierarchy  cell=or13d0
.subckt I3_OR13 C B AN Y VDD VSS
PM1 N_4  AN  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  N_4 N_15 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_15 B   N_16 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_16 C   N_6  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD  N_6 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 N_4 AN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS N_4 N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_6 B   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS C   N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 VSS N_6 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I3_OR13


* Top of hierarchy  cell=or23d0
.subckt I3_OR23 AN C BN Y VDD VSS
PM1 N_3  AN  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  N_3 N_17 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_17 N_7 N_18 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_18 C   N_6  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 N_7  BN  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6
PM6 VDD  N_6 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=7

NM1 N_3 AN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS N_3 N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_6 N_7 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS C   N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_7 BN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
NM6 VSS N_6 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=7
.ends I3_OR23

******************OR AND************************
* Top of hierarchy  cell=ora211d0
.subckt I4_ORA211 C0 B0 A1 A0 VSS Y VDD
PM1 VDD  A0 N_17 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_17 A1 N_6  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_6  B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD  C0 N_6  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD  N_6 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 N_8  A0 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS  A1 N_8  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_8  B0 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_11 C0 N_6  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 VSS  N_6 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I4_ORA211

* Top of hierarchy  cell=ora21d0
.subckt I3_ORA21 B0 A1 A0 Y VDD VSS
PM1 VDD  A0 N_14 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_14 A1 N_5  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_5  B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD  N_5 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 N_6 A0 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS A1 N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_6 B0 N_5 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS N_5 Y  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends I3_ORA21

* Top of hierarchy  cell=ora31d0
.subckt I4_ORA31 B0 A2 A0 A1 Y VDD VSS
PM1 VDD  A1 N_15 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_15 A0 N_16 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_16 A2 N_6  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_6  B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD  N_6 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 VSS A1 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_7 A0 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS A2 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_7 B0 N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 VSS N_6 Y  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I4_ORA31



******************NAND************************

.SUBCKT I2_NAND02 IN1 IN2 VDD VSS OUT1
pmos_1 OUT1 IN2  VDD VDD pmos l=1 w=1 n=1 ro=1 co=1
nmos_1 OUT1 IN2  net1  VSS nmos l=1 w=1 n=1 ro=1 co=1
pmos_2 VDD  IN1  OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=2
nmos_2 net1 IN1  VSS  VSS nmos l=1 w=1 n=1 ro=1 co=2  
.ends I2_NAND02

.subckt I3_NAND03 C B A Y VDD VSS
PM1 VDD C Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 Y   B VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD A Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3

NM1 VSS C N_9 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_9 B N_8 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_8 A Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
.ends I3_NAND03

.subckt I4_NAND04 C B D A VSS VDD Y
PM1 VDD D Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 Y   C VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD B Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 Y   A VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 VSS  D N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_10 C N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_11 B N_9  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_9  A Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends I4_NAND04


* Top of hierarchy  cell=nd12d0
.subckt I2_NAND12 B AN Y VDD VSS
PM1 N_4 AN  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD B   Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 Y   N_4 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3

NM1 N_4  AN  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS  B   N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_12 N_4 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
.ends I2_NAND12


* Top of hierarchy  cell=nd13d0
.subckt I3_NAND13 VSS Y VDD B C AN
PM1 N_4 AN  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD C   Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 Y   B   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD N_4 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 N_4 AN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS C   N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_7 B   N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_6 N_4 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends I3_NAND13


* Top of hierarchy  cell=nd14d0
.subckt I4_NAND14 VSS Y VDD B C D AN

PM1 N_4 AN VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD D   Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 Y   C   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD B   Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 Y   N_4 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 N_4 AN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS D   N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_7 C   N_8 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_8 B   N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_6 N_4 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends I4_NAND14


* Top of hierarchy  cell=nd23d0
.subckt I3_NAND23 AN C BN VSS Y VDD
PM1 N_5 AN VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 Y   C   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM3 VDD N_4 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM4 Y   N_5 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 VDD BN N_4 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=7

NM1 N_5  AN  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS  C   N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM3 N_10 N_4 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM4 N_11 N_5 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 VSS  BN  N_4  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=7
.ends I3_NAND23

* Top of hierarchy  cell=nd24d0
.subckt I4_NAND24 VSS Y VDD D AN C BN
PM1 N_4 AN  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD D   Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 Y   C   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD N_3 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 Y   N_4 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM6 VDD BN  N_3 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=7

NM1 N_4 AN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS D   N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_7 C   N_8 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_8 N_3 N_9 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_9 N_4 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM6 VSS BN  N_3 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=7
.ends I4_NAND24

******************NOR************************
.SUBCKT I2_NOR02 IN1 IN2 VDD VSS OUT1
PM1 VDD  IN1  net1 VDD pmos l=1 w=1 n=1 ro=1 co=1
NM1 VSS  IN1  OUT1  VSS nmos l=1 w=1 n=1 ro=1 co=1
PM2 net1 IN2  OUT1  VDD pmos l=1 w=1 n=1 ro=1 co=2
NM2 OUT1 IN2  VSS  VSS nmos l=1 w=1 n=1  ro=1 co=2
.ends I2_NOR02



* Top of hierarchy  cell=nr03d0
.subckt I3_NOR03 A B C Y VDD VSS

PM1 VDD A N_9 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_9 B N_8 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_8 C Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3

NM1 VSS A Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 Y   B VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS C Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
.ends I3_NOR03


.subckt I4_NOR04 A B C D Y VDD VSS
PM1 VDD  A N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_10 B N_11 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_11 C N_9  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_9  D Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 VSS A  Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 Y   B  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS C  Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 Y   D  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends I4_NOR04

.subckt I2_NOR12 AN B Y VDD VSS
PM1 N_3 AN  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD N_3 N_8 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_8 B   Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3

NM1 N_3 AN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS N_3 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 Y   B   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
.ends I2_NOR12


.subckt I3_NOR13 AN B C Y VDD VSS
PM1 N_3  AN  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  N_3 N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_10 B   N_9  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_9  C   Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 N_3 AN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS N_3 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 Y   B   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS C   Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends I3_NOR13

* Top of hierarchy  cell=nr14d0
.subckt I4_NOR14 D C B AN VSS VDD Y
PM1 N_5  AN  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  N_5 N_15 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_15 B   N_16 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_16 C   N_14 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 N_14 D   Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 N_5 AN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS N_5 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 Y   B   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS C   Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 Y   D   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends I4_NOR14

* Top of hierarchy  cell=nr23d0
.subckt I3_NOR23 C AN BN VSS VDD Y

PM1 N_3  BN  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  AN  N_4  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD  N_4 N_11 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM4 N_11 N_3 N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 N_10 C   Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 N_3 BN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS AN  N_4 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS N_4 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM4 Y   N_3 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 VSS C   Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I3_NOR23

* Top of hierarchy  cell=nr24d0
.subckt I4_NOR24 D C AN BN Y VDD VSS

PM1 N_4  BN  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  AN  N_5  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD  N_5 N_12 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM4 N_12 N_4 N_13 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 N_13 C   N_11 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6
PM6 N_11 D   Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=7

NM1 N_4 BN  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS AN  N_5 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS N_5 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM4 Y   N_4 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 VSS C   Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
NM6 Y   D   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=7
.ends I4_NOR24

******************AOI************************

.subckt I3_AOI21 A0 A1 B0 C0 Y VDD VSS
PM1 N_6  A0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  A1 N_6  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_6  B0 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3

NM1 VSS  A0  N_15 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_15 A1  Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 Y    B0  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3

.ends I3_AOI21

.subckt I3_AOIM21 A1N A0N B0 VSS VDD Y
PM1 VDD  A0N N_14 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_14 A1N N_4  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD  N_4 N_13 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_13 B0  Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 VSS  A0N N_4 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_4  A1N VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  N_4 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 Y    B0  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends I3_AOIM21



.subckt I4_AOI211 A0 A1 B0 C0 Y VDD VSS
PM1 N_6  A0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  A1 N_6  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_6  B0 N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_10 C0 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 VSS  A0  N_15 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_15 A1  Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 Y    B0  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS  C0  Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4

.ends I4_AOI211

.subckt I4_AOI22 B0 B1 A1 A0 VSS VDD Y

PM1 N_8 A0 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD A1 N_8 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_8 B1 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 Y   B0 N_8 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 VSS  A0 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_11 A1 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 Y    B1 N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_10 B0 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends I4_AOI22


.subckt I4_AOI31 A0 A1 A2 B0 VDD Y VSS
PM1 VDD A0 N_7 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_7 A1 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD A2 N_7 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_7 B0 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 VSS  A0 N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_10 A1 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_11 A2 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 Y    B0 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4

.ends I4_AOI31


.subckt I4_AOIM22 B1 B0 A1N A0N VSS VDD Y

PM1 VDD  A0N N_11 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_11 A1N N_2  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_10  B1 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM4 VDD   B0 N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 N_10  N_2 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 VSS  A0N N_2  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_2  A1N VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  B1  N_16 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM4 N_16 B0  Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 Y    N_2 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I4_AOIM22

.subckt I5_AOI221 C0 A0 A1 B1 B0 VDD VSS Y
PM1 N_11 B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  B1 N_11 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_11 A1 N_7  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_7  A0 N_11 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 N_7  C0 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 VSS  B0 N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_12 B1 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 Y    A1 N_13 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_13 A0 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 VSS  C0 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I5_AOI221

.subckt I5_AOI32 VSS Y VDD A1 A0 A2 B1 B0
PM1 VDD  A0 N_12 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_12 A1 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD  A2 N_12 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_12 B1 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 Y    B0 N_12 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 VSS A0 N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_6 A1 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_7 A2 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 Y   B1 N_5 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_5 B0 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends I5_AOI32



******************OAI************************
* Top of hierarchy  cell=oai211d0
.subckt oai211d0 C0 B0 A1 A0 VSS VDD Y

PM1 VDD  A0 N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_10 A1 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 Y    B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD  C0 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 N_9  A0 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS  A1 N_9  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_9  B0 N_16 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_16 C0 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends oai211d0

* Top of hierarchy  cell=oai21d0
.subckt oai21d0 A0 B0 A1 VDD Y VSS
PM1 VDD  A0 N_12 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_12 A1 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 Y    B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3

NM1 N_5  A0 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS  A1 N_5  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_5  B0 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
.ends oai21d0

* Top of hierarchy  cell=oai221d0
.subckt oai221d0 C0 B1 A1 A0 B0 Y VDD VSS

PM1 VDD  A0 N_12 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_12 A1 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 Y    B1 N_13 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_13 B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD  C0 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 N_8 A0 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS A1 N_8 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_8 B1 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_7 B0 N_8 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_7 C0 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends oai221d0

* Top of hierarchy  cell=oai222d0
.subckt oai222d0 B0 A0 A1 B1 C0 C1 Y VDD VSS
PM1 N_9  B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  A0 N_21 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_21 A1 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_9  B1 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 Y    C0 N_20 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6
PM6 N_20 C1 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=7

NM1 N_11 B0 N_8  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_8  A0 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  A1 N_8  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_8  B1 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 N_11 C0 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
NM6 Y    C1 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=7
.ends oai222d0

* Top of hierarchy  cell=oai22d0
.subckt oai22d0 A0 A1 B1 B0 VSS VDD Y
PM1 Y    B1 N_11 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_11 B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD  A0 N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_10 A1 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 N_7 B1 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 Y   B0 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_7 A0 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 VSS A1 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends oai22d0

* Top of hierarchy  cell=oai311d0
.subckt oai311d0 VDD Y VSS C0 B0 A0 A1 A2

PM1 Y   A2 N_7 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_7 A1 N_8 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_8 A0 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD B0 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 Y   C0 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 VSS  A2 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_11 A1 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  A0 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_11 B0 N_20 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_20 C0 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends oai22d0


* Top of hierarchy  cell=oai31d0
.subckt oai31d0 A2 A0 A1 B0 Y VDD VSS
PM1 Y    B0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  A1 N_11 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_11 A0 N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_10 A2 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 Y   B0 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_7 A1 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS A0 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_7 A2 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends oai31d0

* Top of hierarchy  cell=oai321d0
.subckt oai321d0 B1 B0 A0 A1 A2 C0 VDD Y VSS
PM1 Y    A2 N_17 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_17 A1 N_18 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_18 A0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD  B0 N_19 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 N_19 B1 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM6 Y    C0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=7

NM1 VSS  A2 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_11 A1 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  A0 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_11 B0 N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_10 B1 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM6 N_10 C0 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=7
.ends oai321d0

* Top of hierarchy  cell=oai322d0
.subckt oai322d0 VDD Y VSS B0 A0 A1 A2 B1 C0 C1

PM1 VDD  C1 N_8 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_8  C0 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 Y    B1 N_3 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 Y    A2 N_9  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 N_9  A1 N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6
PM6 N_10 A0 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=7
PM7 VDD  B0 N_3  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=9

NM1 N_11 C1 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 Y    C0 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_11 B1 N_13 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_13 A2 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 VSS  A1 N_13 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
NM6 N_13 A0 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=7
NM7 N_13 B0 N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=9
.ends oai322d0

* Top of hierarchy  cell=oai32d0
.subckt oai32d0 A0 B1 A1 A2 B0 Y VDD VSS
PM1 Y    A2 N_16 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_16 A0 N_17 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_17 A1 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD  B0 N_15 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 N_15 B1 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 VSS A2 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_7 A0 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS A1 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_7 B0 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 Y   B1 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends oai32d0

* Top of hierarchy  cell=oai33d0
.subckt oai33d0 VDD Y VSS B2 B1 B0 A1 A0 A2
PM1 Y   A2 N_7 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_7 A0 N_8 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_8 A1 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD B0 N_9 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 N_9 B1 N_6 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM6 N_6 B2 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 VSS  A2 N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_12 A0 VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  A1 N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_12 B0 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 Y    B1 N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM6 N_12 B2 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends oai33d0

* Top of hierarchy  cell=oaim211d0
.subckt oaim211d0 B0 C0 A0N A1N VSS VDD Y

PM1 VDD A1N N_4 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_4 A0N VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD N_4 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 Y   B0  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD C0  Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 N_4  A1N N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_11 A0N VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  N_4 N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_12 B0  N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_10 C0  Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends oaim211d0

* Top of hierarchy  cell=oaim21d0
.subckt oaim21d0 B0 A1N A0N VDD VSS Y

PM1 VDD A0N N_3 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_3 A1N VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD B0  Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 Y   N_3 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4

NM1 N_3  A0N N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_10 A1N VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  B0  N_9  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_9  N_3 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
.ends oaim21d0

* Top of hierarchy  cell=oaim22d0
.subckt oaim22d0 B1 B0 A0N A1N Y VDD VSS

PM1 N_4 A1N VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD A0N N_4 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 Y    N_4 VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM4 VDD  B0  N_18 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 N_18 B1  Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 VSS  A1N N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_11 A0N N_4 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 Y   N_4 N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM4 N_7 B0  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 VSS B1  N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends oaim22d0

* Top of hierarchy  cell=oaim2m11d0
.subckt oaim2m11d0 C0 A0N B0N A1N VDD VSS Y
PM1 N_7 A0N VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD A1N N_7 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_7 B0N N_6 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3

PM4 Y   N_6  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 VDD C0   Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 N_6  A0N N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_12 A1N VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  B0N N_6  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3

NM4 VSS  N_6 N_11 VSS nmos  l=0.5u w=0.6u n=1 ro=1 co=5
NM5 N_11 C0  Y    VSS nmos  l=0.5u w=0.6u n=1 ro=1 co=6
.ends oaim2m11d0

* Top of hierarchy  cell=oaim31d0
.subckt oaim31d0 VSS Y VDD A1N A2N B0 A0N

PM1 VDD N_4 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 Y   B0  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD A2N N_4 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_4 A1N VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD A0N N_4 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 Y   N_4 N_6 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_6 B0  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS A2N N_8 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_8 A1N N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_7 A0N N_4 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends oaim31d0


******************AOR************************

.subckt I3_AOR21 B0 A1 A0 VDD Y VSS
PM1 N_9 A0  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD A1  N_9 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_9 B0  N_2 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM5 VDD N_2 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 VSS  A0  N_10 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_10 A1  N_2  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_2  B0  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM5 VSS  N_2 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends I3_AOR21


.subckt I4_AOR211 C0 B0 A0 A1 VSS Y VDD
PM1 N_9  A1  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD  A0  N_9  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_9  B0  N_18 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_18 C0  N_2  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD  N_2 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 N_2  A1  N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_11 A0  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 VSS  B0  N_2  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_2  C0  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 VSS  N_2 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I4_AOR211

.subckt I4_AOR22 B0 B1 A1 A0 Y VSS VDD

PM1 N_9 A0 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD A1 N_9 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_9 B1 N_6 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_6 B0 N_9 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD N_6 Y  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 VSS  A0  N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_11 A1  N_6  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_6  B1  N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_12 B0  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 VSS  N_6 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6

.ends I4_AOR22

.subckt I4_AOR31 B0 A2 A1 A0 Y VDD VSS
PM1 VDD A0  N_9 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_9 A1  VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 VDD A2  N_9 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 N_9 B0  N_2 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 VDD N_2 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 VSS  A0  N_11 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 N_11 A1  N_12 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_12 A2  N_2  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_2  B0  VSS  VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 VSS  N_2 Y    VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I4_AOR31

.subckt I5_AOR221 VSS Y VDD C0 A0 A1 B1 B0
PM1 N_4  C0  N_12 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_12 A0  N_14 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_14 A1  N_12 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD  B1  N_14 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM5 N_14 B0  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6
PM6 VDD  N_4 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=7

NM1 N_4 C0  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS A0  N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_7 A1  N_4 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_4 B1  N_8 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM5 N_8 B0  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
NM6 VSS N_4 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=7
.ends I5_AOR221

.subckt I5_AOR311 VSS Y VDD A2 A0 A1 B0 C0
PM1 N_4  C0  N_15 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 N_15 B0  N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_10 A1  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=3
PM4 VDD  A0  N_10 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM5 N_10 A2  VDD  VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5
PM6 VDD  N_4 Y    VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=6

NM1 N_4 C0  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS B0  N_4 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_4 A1  N_7 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=3
NM4 N_7 A0  N_8 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM5 N_8 A2  VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
NM6 VSS N_4 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=6
.ends I5_AOR311
******************Logic 4************************






******************Logic 5************************








******************Buffer************************

.subckt BUFF_2 VDD Y VSS A
PM1 N_4 A   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD N_4 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
NM1 N_4 A   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS N_4 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
.ends BUFF_1

.subckt BUFF_3 VDD Y VSS A
PM3 VDD  N_4 Y   VDD pmos  l=0.42u w=0.72u n=1 ro=1 co=1
PM2 Y    N_4 VDD VDD pmos  l=0.42u w=0.72u n=1 ro=1 co=2
PM1 VDD  A   N_4 VDD pmos  l=0.42u w=0.76u n=1 ro=1 co=3
NM3 VSS  N_4 Y   VSS nmos  l=0.5u w=0.34u n=1 ro=1 co=1
NM2 Y    N_4 VSS VSS nmos  l=0.5u w=0.74u n=1 ro=1 co=2
NM1 VSS  A   N_4 VSS nmos  l=0.5u w=0.58u n=1 ro=1 co=3
.ends BUFF_3

******************Delay************************
.subckt DELAY_4 A VSS VDD Y
PM1 N_4 A   VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=1
PM2 VDD N_4 N_3 VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=2
PM3 N_2 N_3 VDD VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=4
PM4 VDD N_2 Y   VDD pmos  l=0.42u w=0.52u n=1 ro=1 co=5

NM1 N_4 A   VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=1
NM2 VSS N_4 N_3 VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=2
NM3 N_2 N_3 VSS VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=4
NM4 VSS N_2 Y   VSS nmos  l=0.5u w=0.5u n=1 ro=1 co=5
.ends DELAY_4