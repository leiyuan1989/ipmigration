* SPICE INPUT		Wed Jul 10 14:00:28 2019	sdbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb1
.subckt sdbfb1 VDD Q QN GND RN SN SI SE D CKN
M1 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M9 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M10 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M11 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_9 N_5 N_29 GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_4 N_55 GND mn5  l=0.5u w=0.5u m=1
M14 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M16 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M17 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_4 N_56 GND mn5  l=0.5u w=0.5u m=1
M20 N_57 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M21 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M23 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M24 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M25 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M26 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M28 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_4 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M34 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M44 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M45 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M46 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M47 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M48 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdbfb1
* SPICE INPUT		Wed Jul 10 14:00:35 2019	sdbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb2
.subckt sdbfb2 VDD Q QN GND RN SN SI SE D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_5 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_4 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_4 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M20 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M21 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M22 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M23 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M24 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M25 N_4 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.52u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M42 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M44 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M45 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M46 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M47 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M48 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdbfb2
* SPICE INPUT		Wed Jul 10 14:00:42 2019	sdbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb1
.subckt sdbrb1 VDD Q QN GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M18 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M19 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M20 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M21 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M22 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M23 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M24 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M42 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M44 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M45 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M46 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M47 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M48 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdbrb1
* SPICE INPUT		Wed Jul 10 14:00:50 2019	sdbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb2
.subckt sdbrb2 VDD Q QN GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M18 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M20 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M21 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M22 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M23 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M24 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M43 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M44 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M45 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M46 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M47 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M48 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
.ends sdbrb2
* SPICE INPUT		Wed Jul 10 14:00:57 2019	sdbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq1
.subckt sdbrq1 VDD Q GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_35 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_35 N_6 N_30 GND mn5  l=0.5u w=0.5u m=1
M6 N_36 SI N_30 GND mn5  l=0.5u w=0.5u m=1
M7 N_36 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_30 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_37 GND mn5  l=0.5u w=0.5u m=1
M10 N_37 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_28 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_28 N_3 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_38 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_38 GND mn5  l=0.5u w=0.5u m=1
M16 Q N_11 N_24 GND mn5  l=0.5u w=0.58u m=1
M17 N_24 N_3 Q GND mn5  l=0.5u w=0.58u m=1
M18 N_24 SN GND GND mn5  l=0.5u w=0.58u m=1
M19 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M20 N_39 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M21 N_39 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_12 N_3 N_26 GND mn5  l=0.5u w=0.5u m=1
M23 N_26 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M24 N_26 SN GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_22 N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M42 Q N_3 N_22 VDD mp5  l=0.42u w=0.76u m=1
M43 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M44 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M45 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M46 N_21 N_3 N_12 VDD mp5  l=0.42u w=0.5u m=1
M47 N_21 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M48 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdbrq1
* SPICE INPUT		Wed Jul 10 14:01:05 2019	sdbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq2
.subckt sdbrq2 VDD Q GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_35 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_35 N_6 N_30 GND mn5  l=0.5u w=0.5u m=1
M6 N_36 SI N_30 GND mn5  l=0.5u w=0.5u m=1
M7 N_36 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_30 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_37 GND mn5  l=0.5u w=0.5u m=1
M10 N_37 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_28 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_28 N_3 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_38 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_12 N_3 N_26 GND mn5  l=0.5u w=0.5u m=1
M16 N_26 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M17 N_26 SN GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 N_24 GND mn5  l=0.5u w=0.72u m=1
M19 N_24 N_3 Q GND mn5  l=0.5u w=0.72u m=1
M20 N_24 SN GND GND mn5  l=0.5u w=0.72u m=1
M21 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M22 N_11 N_5 N_38 GND mn5  l=0.5u w=0.5u m=1
M23 N_39 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M24 N_39 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_21 N_3 N_12 VDD mp5  l=0.42u w=0.5u m=1
M41 N_21 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M42 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M43 N_22 N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M44 Q N_3 N_22 VDD mp5  l=0.42u w=0.96u m=1
M45 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M46 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M47 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M48 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdbrq2
* SPICE INPUT		Wed Jul 10 14:01:12 2019	sdcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb1
.subckt sdcfb1 VDD Q QN GND RN SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_26 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M6 N_47 SI N_26 GND mn5  l=0.5u w=0.5u m=1
M7 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M9 N_48 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_11 N_5 N_49 GND mn5  l=0.5u w=0.5u m=1
M15 N_50 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M16 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M20 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M28 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M32 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M35 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M37 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M38 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M41 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M42 N_14 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M43 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M44 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends sdcfb1
* SPICE INPUT		Wed Jul 10 14:01:19 2019	sdcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb2
.subckt sdcfb2 VDD Q QN GND CKN D SE SI RN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M5 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M10 N_11 N_5 N_49 GND mn5  l=0.5u w=0.5u m=1
M11 N_50 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M12 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_28 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M14 N_47 SI N_28 GND mn5  l=0.5u w=0.5u m=1
M15 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_4 N_28 GND mn5  l=0.5u w=0.5u m=1
M17 N_48 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M25 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 N_14 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M31 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M33 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M35 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M39 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M44 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdcfb2
* SPICE INPUT		Wed Jul 10 14:01:27 2019	sdcfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfq1
.subckt sdcfq1 VDD Q GND CKN D SE SI RN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_5 N_47 GND mn5  l=0.5u w=0.5u m=1
M4 N_48 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M6 N_48 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_44 D GND GND mn5  l=0.5u w=0.5u m=1
M10 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M11 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M13 N_27 N_6 N_44 GND mn5  l=0.5u w=0.5u m=1
M14 N_45 SI N_27 GND mn5  l=0.5u w=0.5u m=1
M15 N_45 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_4 N_27 GND mn5  l=0.5u w=0.5u m=1
M17 N_46 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_47 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M25 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_21 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_12 N_13 N_22 VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M33 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M38 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_10 N_13 N_19 VDD mp5  l=0.42u w=0.52u m=1
M41 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcfq1
* SPICE INPUT		Wed Jul 10 14:01:34 2019	sdcfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfq2
.subckt sdcfq2 VDD Q GND RN SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_48 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_48 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_44 D GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M10 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M12 N_25 N_6 N_44 GND mn5  l=0.5u w=0.5u m=1
M13 N_45 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M14 N_45 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M16 N_46 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_47 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_11 N_5 N_47 GND mn5  l=0.5u w=0.5u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_21 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_12 N_13 N_22 VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M30 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M37 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M38 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_10 N_13 N_19 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
.ends sdcfq2
* SPICE INPUT		Wed Jul 10 14:01:41 2019	sdcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb1
.subckt sdcrb1 VDD Q QN GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M5 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_50 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M13 N_11 N_4 N_49 GND mn5  l=0.5u w=0.5u m=1
M14 N_26 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M15 N_47 SI N_26 GND mn5  l=0.5u w=0.5u m=1
M16 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_5 N_26 GND mn5  l=0.5u w=0.5u m=1
M18 N_48 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M19 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M31 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M35 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M40 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M41 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M44 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrb1
* SPICE INPUT		Wed Jul 10 14:01:49 2019	sdcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb2
.subckt sdcrb2 VDD Q QN GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M5 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_46 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_50 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_50 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M13 N_11 N_4 N_49 GND mn5  l=0.5u w=0.5u m=1
M14 N_26 N_6 N_46 GND mn5  l=0.5u w=0.5u m=1
M15 N_47 SI N_26 GND mn5  l=0.5u w=0.5u m=1
M16 N_47 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_5 N_26 GND mn5  l=0.5u w=0.5u m=1
M18 N_48 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M19 N_48 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_49 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_23 VDD mp5  l=0.42u w=0.52u m=1
M31 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M35 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M40 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M41 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_10 N_13 N_20 VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M44 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrb2
* SPICE INPUT		Wed Jul 10 14:01:56 2019	sdcrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrn1
.subckt sdcrn1 VDD QN GND RN SI SE D CK
M1 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M5 N_42 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M9 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_24 N_6 N_42 GND mn5  l=0.5u w=0.5u m=1
M13 N_43 SI N_24 GND mn5  l=0.5u w=0.5u m=1
M14 N_43 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_5 N_24 GND mn5  l=0.5u w=0.5u m=1
M16 N_44 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_44 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M21 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M28 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_12 N_13 N_21 VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_10 N_13 N_18 VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrn1
* SPICE INPUT		Wed Jul 10 14:02:03 2019	sdcrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrn2
.subckt sdcrn2 VDD QN GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_42 D GND GND mn5  l=0.5u w=0.5u m=1
M5 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_24 N_6 N_42 GND mn5  l=0.5u w=0.5u m=1
M9 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M12 N_43 SI N_24 GND mn5  l=0.5u w=0.5u m=1
M13 N_43 SE GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_5 N_24 GND mn5  l=0.5u w=0.5u m=1
M15 N_44 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M16 N_44 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M26 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_12 N_13 N_21 VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_21 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M36 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 N_13 N_18 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
.ends sdcrn2
* SPICE INPUT		Wed Jul 10 14:02:11 2019	sdcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq1
.subckt sdcrq1 VDD Q GND RN SI SE D CK
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_12 GND GND mn5  l=0.5u w=0.58u m=1
M4 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_13 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_12 RN GND GND mn5  l=0.5u w=0.5u m=1
M8 N_47 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_43 D GND GND mn5  l=0.5u w=0.5u m=1
M10 N_47 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M11 N_11 N_4 N_46 GND mn5  l=0.5u w=0.5u m=1
M12 N_25 N_6 N_43 GND mn5  l=0.5u w=0.5u m=1
M13 N_44 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M14 N_44 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M16 N_45 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M24 Q N_12 N_15 VDD mp5  l=0.42u w=0.76u m=1
M25 N_15 N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M26 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_12 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_21 N_13 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M32 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M33 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M34 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M38 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M39 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_10 N_12 N_19 VDD mp5  l=0.42u w=0.52u m=1
M41 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_22 N_12 N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrq1
* SPICE INPUT		Wed Jul 10 14:02:18 2019	sdcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq2
.subckt sdcrq2 VDD Q GND RN SI SE D CK
M1 N_12 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M4 Q N_12 GND GND mn5  l=0.5u w=0.72u m=1
M5 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_13 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_47 N_13 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_43 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_47 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M12 N_11 N_4 N_46 GND mn5  l=0.5u w=0.5u m=1
M13 N_25 N_6 N_43 GND mn5  l=0.5u w=0.5u m=1
M14 N_44 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M15 N_44 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_45 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 N_10 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_46 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_12 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M25 Q N_12 N_15 VDD mp5  l=0.42u w=0.96u m=1
M26 N_15 N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_22 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_22 N_12 N_13 VDD mp5  l=0.42u w=0.52u m=1
M30 N_21 N_13 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_16 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M33 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M34 N_7 SE N_16 VDD mp5  l=0.42u w=0.52u m=1
M35 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M37 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M38 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M39 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_19 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 N_12 N_19 VDD mp5  l=0.42u w=0.52u m=1
M42 N_20 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdcrq2
* SPICE INPUT		Wed Jul 10 14:02:25 2019	sdnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb1
.subckt sdnfb1 GND QN Q VDD SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M6 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M7 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_17 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_11 N_5 N_18 GND mn5  l=0.5u w=0.5u m=1
M14 N_19 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M15 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M18 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M19 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M24 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M25 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_9 N_5 N_21 VDD mp5  l=0.42u w=0.52u m=1
M27 N_40 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M28 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_41 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M32 N_42 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M33 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M36 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends sdnfb1
* SPICE INPUT		Wed Jul 10 14:02:33 2019	sdnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb2
.subckt sdnfb2 GND QN Q VDD SI SE D CKN
M1 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M3 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M7 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_19 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_5 N_18 GND mn5  l=0.5u w=0.5u m=1
M10 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M14 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_4 N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_17 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M18 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M21 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M22 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M24 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_42 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_41 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M29 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M32 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M33 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_9 N_5 N_21 VDD mp5  l=0.42u w=0.52u m=1
M35 N_40 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M36 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdnfb2
* SPICE INPUT		Wed Jul 10 14:02:40 2019	sdnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb1
.subckt sdnrb1 GND QN Q VDD SI SE D CK
M1 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M3 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_11 N_4 N_18 GND mn5  l=0.5u w=0.5u m=1
M8 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M10 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M13 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M14 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M16 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M18 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M19 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M22 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_42 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M25 N_41 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M26 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M33 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M34 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_9 N_4 N_21 VDD mp5  l=0.42u w=0.52u m=1
M36 N_40 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
.ends sdnrb1
* SPICE INPUT		Wed Jul 10 14:02:47 2019	sdnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb2
.subckt sdnrb2 GND QN Q VDD SI SE D CK
M1 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_19 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_19 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 N_4 N_18 GND mn5  l=0.5u w=0.5u m=1
M6 N_18 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M8 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_17 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_15 GND mn5  l=0.5u w=0.5u m=1
M14 N_16 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M19 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_42 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_42 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M23 N_41 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M24 N_41 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_40 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_38 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_21 SE N_38 VDD mp5  l=0.42u w=0.52u m=1
M31 N_39 N_6 N_21 VDD mp5  l=0.42u w=0.52u m=1
M32 N_39 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_9 N_4 N_21 VDD mp5  l=0.42u w=0.52u m=1
M34 N_40 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdnrb2
* SPICE INPUT		Wed Jul 10 14:02:54 2019	sdnrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrn1
.subckt sdnrn1 GND QN VDD SI SE D CK
M1 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M7 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M9 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M12 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M13 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M14 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M15 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M16 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M18 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M23 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M24 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_20 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_37 N_6 N_20 VDD mp5  l=0.42u w=0.52u m=1
M32 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_9 N_4 N_20 VDD mp5  l=0.42u w=0.52u m=1
M34 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
.ends sdnrn1
* SPICE INPUT		Wed Jul 10 14:03:02 2019	sdnrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrn2
.subckt sdnrn2 GND QN VDD CK D SE SI
M1 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M14 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M21 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M22 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M27 N_9 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M28 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_37 N_6 N_22 VDD mp5  l=0.42u w=0.52u m=1
M30 N_22 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdnrn2
* SPICE INPUT		Wed Jul 10 14:03:09 2019	sdnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq1
.subckt sdnrq1 GND Q VDD CK D SE SI
M1 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M2 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M10 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M12 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M13 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M14 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M19 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M20 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M24 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_9 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M26 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M29 N_37 N_6 N_22 VDD mp5  l=0.42u w=0.52u m=1
M30 N_22 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdnrq1
* SPICE INPUT		Wed Jul 10 14:03:16 2019	sdnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq2
.subckt sdnrq2 GND Q VDD CK D SE SI
M1 N_12 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_18 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_17 GND mn5  l=0.5u w=0.5u m=1
M5 N_18 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_17 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_16 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M10 N_9 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_15 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_15 SI N_7 GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_6 N_14 GND mn5  l=0.5u w=0.5u m=1
M14 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_12 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_40 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M21 N_40 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_39 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M23 N_39 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_10 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_38 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_38 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M27 N_9 N_4 N_19 VDD mp5  l=0.42u w=0.52u m=1
M28 N_37 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_37 N_6 N_19 VDD mp5  l=0.42u w=0.52u m=1
M30 N_19 SE N_36 VDD mp5  l=0.42u w=0.52u m=1
M31 N_36 D VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdnrq2
* SPICE INPUT		Wed Jul 10 14:03:23 2019	sdpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb1
.subckt sdpfb1 VDD Q QN GND CKN D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.58u m=1
M2 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M5 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_46 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_5 N_45 GND mn5  l=0.5u w=0.5u m=1
M9 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M11 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_43 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M15 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M18 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.76u m=1
M23 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M25 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M29 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M30 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M38 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M39 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdpfb1
* SPICE INPUT		Wed Jul 10 14:03:31 2019	sdpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb2
.subckt sdpfb2 VDD Q QN GND CKN D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_46 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M5 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_5 N_45 GND mn5  l=0.5u w=0.5u m=1
M7 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M9 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M10 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_43 N_5 N_9 GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M15 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M18 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CKN GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.96u m=1
M23 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M28 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M32 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_18 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M35 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M38 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M39 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_5 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdpfb2
* SPICE INPUT		Wed Jul 10 14:03:38 2019	sdprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb1
.subckt sdprb1 VDD Q QN GND CK D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M4 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M5 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M10 N_43 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M12 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M13 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M15 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M16 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M17 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M18 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M19 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.76u m=1
M23 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M28 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M29 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M32 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M33 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M35 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M38 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M39 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M40 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M41 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprb1
* SPICE INPUT		Wed Jul 10 14:03:45 2019	sdprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb2
.subckt sdprb2 VDD Q QN GND CK D SE SI SN
M1 Q N_13 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_44 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_46 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_47 SN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_46 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_4 N_45 GND mn5  l=0.5u w=0.5u m=1
M7 N_45 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_10 SN N_44 GND mn5  l=0.5u w=0.5u m=1
M9 N_43 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_43 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M11 N_9 N_5 N_25 GND mn5  l=0.5u w=0.5u m=1
M12 N_42 SE GND GND mn5  l=0.5u w=0.5u m=1
M13 N_42 SI N_25 GND mn5  l=0.5u w=0.5u m=1
M14 N_25 N_6 N_41 GND mn5  l=0.5u w=0.5u m=1
M15 N_41 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_12 GND GND mn5  l=0.5u w=0.72u m=1
M18 N_13 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_12 N_11 N_47 GND mn5  l=0.5u w=0.5u m=1
M20 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M21 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M22 Q N_13 VDD VDD mp5  l=0.42u w=0.96u m=1
M23 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_20 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_19 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M28 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_18 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_18 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M32 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M33 N_17 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M35 N_7 SE N_16 VDD mp5  l=0.42u w=0.5u m=1
M36 N_16 D VDD VDD mp5  l=0.42u w=0.5u m=1
M37 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M38 QN N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M39 N_13 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M41 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprb2
* SPICE INPUT		Wed Jul 10 14:03:53 2019	sdprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq1
.subckt sdprq1 VDD Q GND CK D SN SE SI
M1 N_43 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M2 N_43 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_42 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_44 SN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_41 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_4 N_42 GND mn5  l=0.5u w=0.5u m=1
M7 N_41 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M8 N_12 N_11 N_44 GND mn5  l=0.5u w=0.5u m=1
M9 Q N_11 N_37 GND mn5  l=0.5u w=0.58u m=1
M10 N_40 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_40 N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M12 N_9 N_5 N_24 GND mn5  l=0.5u w=0.5u m=1
M13 N_37 SN GND GND mn5  l=0.5u w=0.58u m=1
M14 N_39 SE GND GND mn5  l=0.5u w=0.5u m=1
M15 N_39 SI N_24 GND mn5  l=0.5u w=0.5u m=1
M16 N_24 N_6 N_38 GND mn5  l=0.5u w=0.5u m=1
M17 N_38 D GND GND mn5  l=0.5u w=0.5u m=1
M18 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M19 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M20 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_18 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_17 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M23 N_17 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_10 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_18 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M27 N_10 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M29 N_12 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_16 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_16 N_5 N_9 VDD mp5  l=0.42u w=0.5u m=1
M32 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M33 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M34 N_15 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_15 N_6 N_7 VDD mp5  l=0.42u w=0.5u m=1
M36 N_7 SE N_14 VDD mp5  l=0.42u w=0.5u m=1
M37 N_14 D VDD VDD mp5  l=0.42u w=0.5u m=1
M38 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_5 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprq1
* SPICE INPUT		Wed Jul 10 14:04:00 2019	sdprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq2
.subckt sdprq2 GND Q VDD CK D SE SI SN
M1 N_20 N_11 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_20 N_4 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 N_3 N_19 GND mn5  l=0.5u w=0.5u m=1
M4 N_19 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_18 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_18 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M7 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_11 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M9 Q N_10 N_14 GND mn5  l=0.5u w=0.72u m=1
M10 N_17 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M12 N_14 SN GND GND mn5  l=0.5u w=0.72u m=1
M13 N_16 SE GND GND mn5  l=0.5u w=0.5u m=1
M14 N_16 SI N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_6 N_5 N_15 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 SE GND GND mn5  l=0.5u w=0.5u m=1
M19 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M20 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M21 N_44 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_44 N_3 N_10 VDD mp5  l=0.42u w=0.5u m=1
M23 N_43 N_4 N_10 VDD mp5  l=0.42u w=0.52u m=1
M24 N_43 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_9 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_42 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 Q N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_11 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_42 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M31 N_8 N_3 N_25 VDD mp5  l=0.42u w=0.5u m=1
M32 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M33 N_41 SI VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_41 N_5 N_25 VDD mp5  l=0.42u w=0.5u m=1
M35 N_11 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M36 N_25 SE N_40 VDD mp5  l=0.42u w=0.5u m=1
M37 N_40 D VDD VDD mp5  l=0.42u w=0.5u m=1
M38 N_5 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdprq2