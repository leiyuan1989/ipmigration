//* No part of this file can be released without the consent of SMIC.
//************************************************************************************************************                                                                                                                                                   
//* SMIC 0.11um Mixed Signal 1P6M(1P5M, 1P7M, 1P8M) 1.2V/3.3V SPICE model (for SPECTRE only) //*                                                                                                                                                     
//************************************************************************************************************                                                                                                                                                   
//*                                                                                                                                                                                                                                                              
//* Release version    : 1.14                                                                                                                                                                                                                                     
//*                                                                                                                                                                                                                                                              
//* Release date       : 03/28/2016                                                                                                                                                                                                                              
//*                                                                                                                                                                                                                                                              
//* Simulation tool    : Cadence spectre V10.1.1                                                                                                                                                                                                 
//*                                                                                                                                                                                                                                                              
//*  Inductor   :                                                                                                                                                                                                                                                
//* *  *------------------------*-----------------------------------------------------------------------------------------------------*
//*    |  Turn, Radius & Width  |T=1~3 step 0.5,W=5~13.5um,R=1.7071*W+16.378~120um;T=3.5~5.0 step 0.5,W=5~8um,R=1.7071*W+16.378~120um |
//* *  *------------------------*-----------------------------------------------------------------------------------------------------*
//*    |        Model Name      |      ind_rf_pgs_n                      										  |            
//* *  *------------------------*-----------------------------------------------------------------------------------------------------*
simulator lang=spectre  insensitive=yes
subckt ind_rf_pgs_n (PLUS MINUS)
parameters r=6e-05 radius_=0.00833333*(r/1e-06-0) w=8e-06 w_=0.0666667*(w/1e-06-0) n=3  \
T0=(n==1.5) \
T1=(radius_>=0.416958) \
T2=(w_+7.291667e-01*radius_>=0.904432) \
T3=(w_>=0.6004) \
T4=(radius_>=0.416375) \
T5=(radius_>=0.708625) \
T6=(w_+7.291667e-01*radius_>=0.903207) \
T7=(w_>=0.5996) \
T8=(radius_>=0.708042) \
T9=(n==1) \
T10=(n==2.5) \
T11=(n==2) \
T12=(n==3.5) \
T13=(n==3) \
T14=(n==4.5) \
T15=(n==4) \
T16=(n==5) \
S0=T0*(1-T1)*(1-T2) \
noS0=(1-S0) \
S1=T0*(1-T3)*T4*(1-T5)*noS0 \
noS1=(1-S1)*noS0 \
S2=T0*T6*T7*(1-T5)*noS1 \
noS2=(1-S2)*noS1 \
S3=T0*(1-T3)*T8*noS2 \
noS3=(1-S3)*noS2 \
S4=T0*T8*T7*noS3 \
noS4=(1-S4)*noS3 \
S5=T9*(1-T1)*(1-T2)*noS4 \
noS5=(1-S5)*noS4 \
S6=T9*(1-T3)*T4*(1-T5)*noS5 \
noS6=(1-S6)*noS5 \
S7=T9*T6*T7*(1-T5)*noS6 \
noS7=(1-S7)*noS6 \
S8=T9*(1-T3)*T8*noS7 \
noS8=(1-S8)*noS7 \
S9=T9*T8*T7*noS8 \
noS9=(1-S9)*noS8 \
S10=T10*(1-T1)*(1-T2)*noS9 \
noS10=(1-S10)*noS9 \
S11=T10*(1-T3)*T4*(1-T5)*noS10 \
noS11=(1-S11)*noS10 \
S12=T10*T6*T7*(1-T5)*noS11 \
noS12=(1-S12)*noS11 \
S13=T10*(1-T3)*T8*noS12 \
noS13=(1-S13)*noS12 \
S14=T10*T8*T7*noS13 \
noS14=(1-S14)*noS13 \
S15=T11*(1-T1)*(1-T2)*noS14 \
noS15=(1-S15)*noS14 \
S16=T11*(1-T3)*T4*(1-T5)*noS15 \
noS16=(1-S16)*noS15 \
S17=T11*T6*T7*(1-T5)*noS16 \
noS17=(1-S17)*noS16 \
S18=T11*(1-T3)*T8*noS17 \
noS18=(1-S18)*noS17 \
S19=T11*T8*T7*noS18 \
noS19=(1-S19)*noS18 \
S20=T12*(1-T1)*noS19 \
noS20=(1-S20)*noS19 \
S21=T12*T4*(1-T5)*noS20 \
noS21=(1-S21)*noS20 \
S22=T12*T8*noS21 \
noS22=(1-S22)*noS21 \
S23=T13*(1-T1)*(1-T2)*noS22 \
noS23=(1-S23)*noS22 \
S24=T13*(1-T3)*T4*(1-T5)*noS23 \
noS24=(1-S24)*noS23 \
S25=T13*T6*T7*(1-T5)*noS24 \
noS25=(1-S25)*noS24 \
S26=T13*(1-T3)*T8*noS25 \
noS26=(1-S26)*noS25 \
S27=T13*T8*T7*noS26 \
noS27=(1-S27)*noS26 \
S28=T14*(1-T1)*noS27 \
noS28=(1-S28)*noS27 \
S29=T14*T4*(1-T5)*noS28 \
noS29=(1-S29)*noS28 \
S30=T14*T8*noS29 \
noS30=(1-S30)*noS29 \
S31=T15*(1-T1)*noS30 \
noS31=(1-S31)*noS30 \
S32=T15*T4*(1-T5)*noS31 \
noS32=(1-S32)*noS31 \
S33=T15*T8*noS32 \
noS33=(1-S33)*noS32 \
S34=T16*(1-T1)*noS33 \
noS34=(1-S34)*noS33 \
S35=T16*T4*(1-T5)*noS34 \
noS35=(1-S35)*noS34 \
S36=T16*T8*noS35 \
noS36=(1-S36)*noS35 \
V0_part1=6.706940e-02*S0+8.771798e-03*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V0_part2=V0_part1+0.000000e+00*S10+(-4.500103e-01)*S11+1.018617e-01*S12+(-1.801514e+00)*S13+0.000000e+00*S14+(-2.480988e+00)*S15+(-4.302653e+00)*S16+0.000000e+00*S17+1.165178e+00*S18+(-2.938107e+01)*S19 \
V0_part3=V0_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+(-8.626834e+00)*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29 \
V0=V0_part3+(-1.205511e+01)*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36 \
V1_part1=2.686316e+01*S0+2.769156e+01*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V1_part2=V1_part1+0.000000e+00*S10+1.277478e+01*S11+3.501357e-01*S12+1.604120e+01*S13+0.000000e+00*S14+3.357469e+01*S15+2.824707e+01*S16+0.000000e+00*S17+3.704576e+01*S18+4.554832e+01*S19 \
V1_part3=V1_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+2.179308e+01*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29 \
V1=V1_part3+4.036215e+01*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36 \
V2_part1=(-1.039065e+01)*S0+(-1.114054e+01)*S1+0.000000e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V2_part2=V2_part1+0.000000e+00*S10+9.563871e-01*S11+5.092456e-02*S12+(-1.354546e+00)*S13+0.000000e+00*S14+1.473535e+00*S15+(-1.700649e+00)*S16+0.000000e+00*S17+(-3.901627e+01)*S18+6.324147e+00*S19 \
V2_part3=V2_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+0.000000e+00*S25+5.708420e-01*S26+0.000000e+00*S27+0.000000e+00*S28+0.000000e+00*S29 \
V2=V2_part3+(-1.016759e+01)*S30+0.000000e+00*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+0.000000e+00*S36 \
V3_part1=(-9.289502e-02)*S0+(-2.423093e-01)*S1+1.786207e+01*S2+(-4.714740e-01)*S3+(-4.906457e-01)*S4+(-1.908046e-01)*S5+(-3.697507e-01)*S6+(-1.288413e-01)*S7+(-7.124345e-01)*S8+(-3.298215e-01)*S9 \
V3_part2=V3_part1+(-8.707372e-02)*S10+(-1.215435e+00)*S11+8.294896e-03*S12+(-5.237036e-01)*S13+(-9.341215e-01)*S14+(-2.868522e-01)*S15+(-4.317691e-01)*S16+(-1.138101e-01)*S17+(-8.963756e-01)*S18+(-5.279721e-01)*S19 \
V3_part3=V3_part2+(-2.424475e-01)*S20+(-6.334610e-01)*S21+(-1.230426e+00)*S22+(-3.186449e-01)*S23+(-4.722558e-01)*S24+6.166916e-02*S25+(-1.322141e+00)*S26+(-5.430105e-01)*S27+(-7.808132e-01)*S28+(-6.813459e-01)*S29 \
V3=V3_part3+(-1.460057e+00)*S30+(-2.201382e+00)*S31+(-6.698481e-01)*S32+(-1.395894e+00)*S33+(-2.591356e-01)*S34+(-5.830727e-01)*S35+(-7.948682e+00)*S36 \
V4_part1=6.296895e-01*S0+6.428929e-01*S1+(-4.310579e-01)*S2+9.272212e-01*S3+4.883327e-01*S4+2.217717e-01*S5+3.399495e-01*S6+1.274319e-01*S7+5.778129e-03*S8+1.955272e-01*S9 \
V4_part2=V4_part1+7.576609e-01*S10+1.277118e+00*S11+5.681789e-01*S12+(-2.301695e+00)*S13+9.048445e-01*S14+6.813941e-01*S15+1.637456e+00*S16+1.216810e+00*S17+1.648160e+00*S18+1.250411e+00*S19 \
V4_part3=V4_part2+2.310374e+00*S20+2.553091e+00*S21+2.995839e+00*S22+2.874484e+00*S23+2.254376e+00*S24+4.252402e-01*S25+5.360258e-01*S26+8.146851e-01*S27+4.579948e+00*S28+3.213587e+00*S29 \
V4=V4_part3+3.293119e+00*S30+(-3.577007e+00)*S31+2.960452e+00*S32+2.990745e+00*S33+3.244294e+00*S34+3.396598e+00*S35+1.384057e+00*S36 \
V5_part1=1.169767e-01*S0+1.851693e-01*S1+5.982505e+00*S2+2.192013e-01*S3+8.441039e-01*S4+2.967490e-01*S5+4.342589e-01*S6+5.474076e-01*S7+1.698185e+00*S8+1.058230e+00*S9 \
V5_part2=V5_part1+8.076078e-01*S10+1.408243e+00*S11+9.936499e-01*S12+4.089479e+00*S13+1.433009e+00*S14+4.650567e-01*S15+1.905050e-01*S16+1.399333e-01*S17+3.164189e-01*S18+3.239662e-01*S19 \
V5_part3=V5_part2+2.441519e-01*S20+3.372593e-01*S21+4.846975e-01*S22+1.996434e-01*S23+2.545152e-01*S24+1.704969e+00*S25+2.563397e+00*S26+1.738104e+00*S27+2.507950e+00*S28+4.291957e-01*S29 \
V5=V5_part3+6.082943e-01*S30+3.707499e+00*S31+3.631538e-01*S32+5.245692e-01*S33+3.123231e-01*S34+4.160737e-01*S35+7.586608e+00*S36 \
V6_part1=(-4.739273e-03)*S0+(-7.592025e-03)*S1+(-4.692337e-02)*S2+(-3.532433e-03)*S3+(-1.310795e-02)*S4+(-5.911782e-03)*S5+(-4.730840e-03)*S6+(-5.857365e-04)*S7+2.286120e-03*S8+1.294234e-02*S9 \
V6_part2=V6_part1+(-1.497430e-02)*S10+(-1.704554e-02)*S11+(-1.182418e-02)*S12+2.453258e-01*S13+(-2.186761e-02)*S14+(-1.829577e-02)*S15+(-5.598186e-02)*S16+(-3.610758e-02)*S17+(-9.844816e-02)*S18+(-1.028756e-01)*S19 \
V6_part3=V6_part2+(-4.237168e-02)*S20+(-1.526212e-01)*S21+(-3.458138e-01)*S22+(-5.825180e-02)*S23+(-1.062814e-01)*S24+3.172584e-02*S25+6.011305e-02*S26+(-2.428761e-02)*S27+3.090677e-02*S28+(-2.340828e-01)*S29 \
V6=V6_part3+(-4.961552e-01)*S30+7.569500e-01*S31+(-1.993801e-01)*S32+(-3.853702e-01)*S33+(-9.996175e-02)*S34+(-2.833185e-01)*S35+(-1.295014e-02)*S36 \
V7_part1=7.116180e-01*S0+7.807401e-01*S1+2.538904e+00*S2+8.278810e-01*S3+7.725477e-01*S4+2.924509e-01*S5+3.129286e-01*S6+2.880087e-01*S7+3.833444e-01*S8+3.261259e-01*S9 \
V7_part2=V7_part1+1.671874e+00*S10+1.848279e+00*S11+1.656505e+00*S12+1.843852e+00*S13+1.854901e+00*S14+1.010962e+00*S15+1.236429e+00*S16+1.152742e+00*S17+1.342242e+00*S18+1.298815e+00*S19 \
V7_part3=V7_part2+3.281753e+00*S20+3.658960e+00*S21+4.080756e+00*S22+2.431126e+00*S23+2.575358e+00*S24+2.129600e+00*S25+2.508239e+00*S26+2.379545e+00*S27+4.821243e+00*S28+5.657376e+00*S29 \
V7=V7_part3+6.252351e+00*S30+3.509719e+00*S31+4.384555e+00*S32+4.800055e+00*S33+5.839553e+00*S34+6.503209e+00*S35+6.566754e+00*S36 \
V8_part1=(-5.446428e-03)*S0+(-6.080998e-02)*S1+1.797027e-01*S2+(-1.356022e-01)*S3+(-6.880945e-02)*S4+(-1.375212e-02)*S5+(-3.146708e-02)*S6+(-1.352583e-02)*S7+(-5.206480e-02)*S8+(-4.152714e-02)*S9 \
V8_part2=V8_part1+(-1.512999e-02)*S10+(-1.602196e-01)*S11+(-5.722022e-03)*S12+(-4.692003e-01)*S13+(-1.629772e-01)*S14+(-2.958944e-02)*S15+(-4.717413e-02)*S16+(-1.128315e-02)*S17+(-1.112002e-01)*S18+(-4.218930e-02)*S19 \
V8_part3=V8_part2+1.330694e-01*S20+3.995494e-02*S21+(-1.434420e-01)*S22+3.683949e-02*S23+(-5.587386e-02)*S24+(-6.680990e-02)*S25+(-4.975247e-01)*S26+(-2.234247e-01)*S27+9.057408e-02*S28+2.593494e-01*S29 \
V8=V8_part3+(-1.434051e-01)*S30+(-4.630265e-01)*S31+7.298007e-02*S32+(-2.404610e-01)*S33+5.187780e-01*S34+2.988594e-01*S35+(-1.232476e+00)*S36 \
V9_part1=7.751124e+00*S0+2.397491e+00*S1+(-9.807390e-02)*S2+(-1.201800e+00)*S3+(-5.174376e-01)*S4+(-2.977978e-01)*S5+(-5.534069e-01)*S6+(-1.855803e-01)*S7+(-5.422862e-01)*S8+(-3.612400e-01)*S9 \
V9_part2=V9_part1+(-4.783310e-01)*S10+(-9.312847e-01)*S11+(-3.252625e-01)*S12+(-1.728913e+00)*S13+(-8.605138e-01)*S14+(-5.155078e-01)*S15+(-1.939915e+00)*S16+(-3.593077e-01)*S17+(-1.890633e+00)*S18+(-9.771018e-01)*S19 \
V9_part3=V9_part2+6.736491e-01*S20+(-6.531415e+00)*S21+(-8.389289e+00)*S22+(-1.717357e-01)*S23+(-3.632447e+00)*S24+(-3.605967e-01)*S25+(-2.219429e+00)*S26+(-1.271501e+00)*S27+(-4.048428e-01)*S28+(-8.084475e+00)*S29 \
V9=V9_part3+(-1.652002e+01)*S30+(-4.312012e-01)*S31+(-6.205910e+00)*S32+(-1.251144e+01)*S33+(-1.466552e+00)*S34+(-1.104714e+01)*S35+(-2.715491e+00)*S36 \
V10_part1=9.476931e+00*S0+6.111834e+00*S1+6.979741e-01*S2+(-4.250540e+00)*S3+1.780199e+00*S4+1.790693e+00*S5+1.586127e+00*S6+7.258931e-01*S7+8.027211e-01*S8+5.960280e-01*S9 \
V10_part2=V10_part1+4.309468e+00*S10+4.111787e+00*S11+2.510700e+00*S12+3.276203e+00*S13+2.860098e+00*S14+4.364785e+00*S15+1.656504e+00*S16+8.816777e-01*S17+6.848594e-01*S18+8.790573e-01*S19 \
V10_part3=V10_part2+5.185822e+00*S20+4.367516e+00*S21+4.188219e+00*S22+2.218726e+00*S23+3.218946e+00*S24+2.400682e+00*S25+4.190576e+00*S26+2.854699e+00*S27+5.616805e+00*S28+6.982942e+00*S29 \
V10=V10_part3+5.224920e-01*S30+5.669122e+00*S31+5.242096e+00*S32+1.292596e+00*S33+8.137485e+00*S34+8.018648e+00*S35+6.843527e+00*S36 \
V11_part1=8.909352e-01*S0+3.959053e+00*S1+3.029481e-01*S2+6.081374e+00*S3+4.574577e-01*S4+1.554572e-01*S5+2.473651e-01*S6+2.132166e-01*S7+3.290281e-01*S8+3.416173e-01*S9 \
V11_part2=V11_part1+3.411958e-01*S10+4.825211e-01*S11+5.079478e-01*S12+7.495833e-01*S13+7.296555e-01*S14+2.517451e-01*S15+2.085019e+00*S16+1.296095e+00*S17+2.917370e+00*S18+1.981609e+00*S19 \
V11_part3=V11_part2+2.518205e+00*S20+6.141167e+00*S21+6.431519e+00*S22+1.302054e+00*S23+3.724322e+00*S24+5.296305e-01*S25+9.384876e-01*S26+9.980297e-01*S27+5.634377e-01*S28+7.300617e+00*S29 \
V11=V11_part3+1.563778e+01*S30+3.846250e-01*S31+5.544469e+00*S32+1.159924e+01*S33+4.756099e+00*S34+8.914700e+00*S35+1.274704e+00*S36 \
V12_part1=(-3.577463e-02)*S0+(-9.256965e-02)*S1+8.049946e-03*S2+9.056658e-01*S3+(-8.749147e-02)*S4+(-1.040380e-02)*S5+(-2.642379e-02)*S6+(-1.520850e-02)*S7+(-4.747235e-02)*S8+(-3.536408e-02)*S9 \
V12_part2=V12_part1+(-6.263984e-02)*S10+(-1.613166e-01)*S11+(-1.115672e-01)*S12+(-2.620911e-01)*S13+(-2.942665e-01)*S14+(-5.948992e-02)*S15+(-2.773394e-02)*S16+(-2.903326e-02)*S17+2.889849e-02*S18+(-2.674676e-02)*S19 \
V12_part3=V12_part2+(-2.591100e-02)*S20+1.255788e-01*S21+(-8.873569e-02)*S22+(-6.464781e-02)*S23+(-4.839156e-02)*S24+(-1.263540e-01)*S25+(-3.681345e-01)*S26+(-3.394479e-01)*S27+(-1.427899e-01)*S28+2.673966e-02*S29 \
V12=V12_part3+9.836086e-01*S30+(-1.853872e-02)*S31+(-6.276313e-03)*S32+5.724359e-01*S33+2.839127e-02*S34+1.217368e-02*S35+(-9.227734e-01)*S36 \
V13_part1=2.330734e+00*S0+2.609357e+00*S1+1.396846e+00*S2+1.575905e+00*S3+1.780724e+00*S4+6.510387e-01*S5+6.911042e-01*S6+6.265905e-01*S7+7.167472e-01*S8+6.870031e-01*S9 \
V13_part2=V13_part1+3.731723e+00*S10+4.104539e+00*S11+3.768018e+00*S12+4.365816e+00*S13+4.288957e+00*S14+2.309483e+00*S15+2.214317e+00*S16+2.000167e+00*S17+2.345857e+00*S18+2.212401e+00*S19 \
V13_part3=V13_part2+6.122053e+00*S20+6.732712e+00*S21+7.393934e+00*S22+4.285396e+00*S23+4.702337e+00*S24+4.704423e+00*S25+5.634007e+00*S26+5.387294e+00*S27+1.007708e+01*S28+1.053492e+01*S29 \
V13=V13_part3+1.108651e+01*S30+7.216084e+00*S31+8.093918e+00*S32+8.636174e+00*S33+1.109132e+01*S34+1.217124e+01*S35+1.432041e+01*S36 \
V14_part1=1.444372e-01*S0+5.009751e-02*S1+(-1.523184e-02)*S2+(-9.666590e-01)*S3+(-1.086537e-01)*S4+(-1.249719e-02)*S5+(-2.007722e-02)*S6+(-1.121271e-02)*S7+(-6.158413e-02)*S8+(-4.495382e-02)*S9 \
V14_part2=V14_part1+5.910561e-02*S10+(-7.996590e-02)*S11+1.017180e-01*S12+(-3.973623e-01)*S13+(-3.241576e-02)*S14+(-4.678003e-03)*S15+(-2.290458e-01)*S16+(-5.975714e-02)*S17+(-4.515763e-01)*S18+(-2.293367e-01)*S19 \
V14_part3=V14_part2+2.631907e-02*S20+(-8.236196e-01)*S21+(-1.487003e+00)*S22+(-7.200195e-02)*S23+(-4.498803e-01)*S24+9.139253e-02*S25+(-4.741281e-01)*S26+(-1.667234e-01)*S27+8.731918e-01*S28+(-7.608085e-01)*S29 \
V14=V14_part3+(-3.152057e+00)*S30+5.107840e-02*S31+(-8.146088e-01)*S32+(-2.595040e+00)*S33+1.690856e-01*S34+(-9.553339e-01)*S35+(-9.921976e-01)*S36 \
V15_part1=1.307742e+00*S0+1.296546e+00*S1+3.598787e-01*S2+(-3.518191e-01)*S3+2.270946e+00*S4+3.049234e-01*S5+8.827302e-01*S6+9.163181e-01*S7+6.594643e-01*S8+6.403707e-01*S9 \
V15_part2=V15_part1+1.257224e+00*S10+9.546523e-01*S11+1.105548e+00*S12+(-4.447668e-01)*S13+1.254015e+00*S14+1.159837e+00*S15+7.462046e-01*S16+1.330943e+00*S17+3.751647e-01*S18+1.405297e+00*S19 \
V15_part3=V15_part2+1.042797e+00*S20+2.095157e-01*S21+8.662223e-01*S22+1.495626e+00*S23+6.251655e-01*S24+3.582023e-01*S25+3.035965e-01*S26+1.063137e+00*S27+5.992943e-01*S28+7.156160e-01*S29 \
V15=V15_part3+(-6.171904e-01)*S30+(-5.824140e-02)*S31+5.477193e-01*S32+(-5.592391e-01)*S33+6.747078e-01*S34+5.362591e-01*S35+(-1.537855e-01)*S36 \
V16_part1=(-1.370037e-01)*S0+(-1.727206e-01)*S1+(-7.561592e-02)*S2+1.390068e+00*S3+(-3.434252e-01)*S4+2.130890e+00*S5+1.146053e+00*S6+5.322099e-01*S7+9.867898e-02*S8+2.223594e-01*S9 \
V16_part2=V16_part1+1.659125e+00*S10+1.285092e+00*S11+7.151121e-01*S12+1.689066e+00*S13+4.096876e-01*S14+1.975322e+00*S15+1.651248e+00*S16+6.151373e-01*S17+1.461130e+00*S18+5.144222e-01*S19 \
V16_part3=V16_part2+1.383585e+00*S20+1.759201e+00*S21+1.575817e+00*S22+1.386591e+00*S23+1.827779e+00*S24+1.127174e+00*S25+1.289875e+00*S26+5.207719e-01*S27+1.709245e+00*S28+1.742772e+00*S29 \
V16=V16_part3+2.313266e+00*S30+2.798172e+00*S31+1.785027e+00*S32+2.044150e+00*S33+2.090951e+00*S34+1.896995e+00*S35+2.857290e+00*S36 \
V17_part1=(-3.989884e-01)*S0+(-4.577185e-01)*S1+(-7.217999e-02)*S2+1.087649e+00*S3+4.513530e-01*S4+1.305547e+00*S5+(-6.724217e-02)*S6+9.037756e-02*S7+(-4.049434e-01)*S8+(-8.834163e-02)*S9 \
V17_part2=V17_part1+3.452572e-01*S10+4.329651e-01*S11+1.575463e-01*S12+3.774640e-01*S13+7.637779e-03*S14+8.913676e-01*S15+3.886114e-01*S16+5.165487e-01*S17+(-1.709497e-01)*S18+(-2.096461e-01)*S19 \
V17_part3=V17_part2+(-3.831012e-01)*S20+6.609266e-01*S21+(-1.696100e-01)*S22+8.589805e-02*S23+7.275795e-01*S24+2.017367e-01*S25+1.123879e-01*S26+(-1.568522e-01)*S27+(-5.640837e-02)*S28+1.361940e-01*S29 \
V17=V17_part3+6.835730e-01*S30+1.312543e+00*S31+4.297228e-01*S32+1.060935e+00*S33+(-1.293243e-01)*S34+7.528523e-01*S35+7.545436e-01*S36 \
V18_part1=(-5.456904e-01)*S0+(-1.452313e+00)*S1+(-1.851381e+00)*S2+6.113579e-01*S3+(-1.437075e+00)*S4+(-4.920300e+01)*S5+(-1.441278e+01)*S6+(-5.716984e+00)*S7+(-3.040550e+01)*S8+(-3.748293e+00)*S9 \
V18_part2=V18_part1+(-1.395382e+00)*S10+(-1.497044e+00)*S11+(-2.919557e+00)*S12+(-1.931752e+00)*S13+(-2.787009e+00)*S14+(-2.541776e-01)*S15+(-1.899330e-01)*S16+(-1.486988e+00)*S17+(-1.916124e+00)*S18+3.093284e+00*S19 \
V18_part3=V18_part2+(-1.973750e+00)*S20+(-1.312415e+00)*S21+(-2.132076e+00)*S22+(-1.578094e+00)*S23+(-1.282793e+00)*S24+(-2.225450e+00)*S25+(-9.608144e-01)*S26+(-2.714117e+00)*S27+(-1.704528e+00)*S28+(-2.308929e+00)*S29 \
V18=V18_part3+(-9.346961e-01)*S30+(-3.586042e+00)*S31+(-1.483306e+00)*S32+(-2.261530e+00)*S33+(-1.783179e+00)*S34+(-2.123020e+00)*S35+(-3.335822e+00)*S36 \
V19_part1=1.460053e+00*S0+1.520751e+00*S1+9.142988e+00*S2+2.161668e+01*S3+6.752977e+00*S4+1.425578e+01*S5+2.355393e+01*S6+3.443974e+01*S7+3.027850e+01*S8+7.923439e+00*S9 \
V19_part2=V19_part1+8.997682e+00*S10+6.284541e+00*S11+1.193903e+01*S12+5.843808e+00*S13+9.144980e+00*S14+1.382596e+00*S15+2.299435e+00*S16+9.218756e+00*S17+9.491084e-01*S18+7.466201e-02*S19 \
V19_part3=V19_part2+1.039116e+01*S20+8.270420e+00*S21+9.122730e+00*S22+9.448116e+00*S23+9.129488e+00*S24+1.089746e+01*S25+5.569080e+00*S26+9.394180e+00*S27+1.011072e+01*S28+1.001663e+01*S29 \
V19=V19_part3+1.593624e+00*S30+2.329013e+01*S31+9.156837e+00*S32+9.162154e+00*S33+1.004937e+01*S34+1.020184e+01*S35+9.747134e+00*S36 \
V20_part1=5.445980e+00*S0+7.386807e+00*S1+4.303885e+00*S2+1.009686e+01*S3+5.788542e+00*S4+1.611026e+02*S5+3.002534e+01*S6+(-7.656726e-01)*S7+5.851291e+01*S8+9.517763e+00*S9 \
V20_part2=V20_part1+7.485159e+00*S10+7.592379e+00*S11+8.374113e+00*S12+8.982189e+00*S13+1.063205e+01*S14+4.144060e+00*S15+5.599124e+00*S16+5.182955e+00*S17+1.396399e+01*S18+5.851709e+00*S19 \
V20_part3=V20_part2+1.083291e+01*S20+1.076820e+01*S21+1.118420e+01*S22+8.488361e+00*S23+6.918040e+00*S24+8.823002e+00*S25+9.112589e+00*S26+1.111889e+01*S27+1.252534e+01*S28+1.337112e+01*S29 \
V20=V20_part3+1.823605e+01*S30+2.993995e+01*S31+1.033891e+01*S32+1.240944e+01*S33+1.312825e+01*S34+1.255251e+01*S35+1.614563e+01*S36 \
V21_part1=4.659939e-01*S0+1.314149e+00*S1+4.531666e-01*S2+1.000000e+04*S3+2.806292e-01*S4+1.367659e+02*S5+1.285027e+02*S6+2.569182e+01*S7+1.596592e+02*S8+9.742963e+01*S9 \
V21_part2=V21_part1+3.748924e-01*S10+2.156257e+00*S11+8.531187e-01*S12+1.086533e+01*S13+4.281221e-03*S14+9.416375e-01*S15+3.460650e-01*S16+2.724990e-01*S17+1.384087e+00*S18+(-4.707743e-01)*S19 \
V21_part3=V21_part2+2.356716e-01*S20+8.500216e-01*S21+2.895944e+00*S22+1.981434e-01*S23+2.958536e-01*S24+3.155801e-01*S25+4.359593e-01*S26+2.804147e-01*S27+3.258652e-01*S28+2.736132e-01*S29 \
V21=V21_part3+8.677640e-01*S30+2.368956e+03*S31+9.337059e-01*S32+(-3.333135e+03)*S33+3.623110e-01*S34+2.092545e-01*S35+4.025291e+00*S36 \
V22_part1=1.948701e+00*S0+9.633530e-01*S1+(-1.375805e-01)*S2+9.646952e+02*S3+(-2.174640e-01)*S4+5.556796e+01*S5+7.323826e+00*S6+9.245893e+01*S7+(-2.306778e+01)*S8+1.981090e+00*S9 \
V22_part2=V22_part1+5.677823e-01*S10+(-7.885912e-01)*S11+2.171777e-01*S12+(-7.168509e+00)*S13+(-2.530213e-01)*S14+1.466658e+00*S15+1.225579e-01*S16+(-3.110697e-01)*S17+2.660360e-02*S18+2.239781e+00*S19 \
V22_part3=V22_part2+7.497187e-02*S20+4.098636e-02*S21+2.854330e-01*S22+(-6.184207e-02)*S23+(-3.368640e-01)*S24+8.393687e-02*S25+(-2.734967e-01)*S26+(-1.757087e-01)*S27+(-2.897189e-01)*S28+1.677804e-01*S29 \
V22=V22_part3+(-6.808402e-01)*S30+3.857229e+02*S31+2.076738e+00*S32+8.368711e-01*S33+(-4.333246e-01)*S34+4.824308e-02*S35+3.815841e+01*S36 \
V23_part1=(-1.019941e+00)*S0+(-1.313381e+00)*S1+1.759519e-01*S2+1.377262e+02*S3+3.499562e-01*S4+(-1.062172e+02)*S5+(-1.100103e+02)*S6+(-1.910736e+01)*S7+(-1.323562e+02)*S8+(-6.117874e+01)*S9 \
V23_part2=V23_part1+(-2.423258e-01)*S10+(-1.720243e+00)*S11+(-4.576922e-01)*S12+(-5.291537e+00)*S13+1.094384e+00*S14+(-5.920735e-01)*S15+6.551917e-01*S16+2.810896e-01*S17+(-9.770630e-01)*S18+(-4.688945e-02)*S19 \
V23_part3=V23_part2+1.555633e-01*S20+(-5.812307e-01)*S21+(-4.796199e+00)*S22+2.451517e-01*S23+6.245170e-01*S24+2.513817e-01*S25+5.103610e-01*S26+4.341919e-01*S27+5.083513e-01*S28+1.997432e-01*S29 \
V23=V23_part3+(-8.582048e-02)*S30+1.007324e+02*S31+(-1.995307e+00)*S32+1.000000e+04*S33+7.863970e-01*S34+3.744624e-01*S35+4.310572e+02*S36 \
V24_part1=(-2.050492e+00)*S0+0.000000e+00*S1+(-9.611695e+01)*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+(-2.986037e+00)*S6+(-4.834384e+00)*S7+(-9.337762e+00)*S8+(-1.269940e+01)*S9 \
V24_part2=V24_part1+0.000000e+00*S10+(-4.711676e+02)*S11+(-1.707345e+02)*S12+(-7.224588e+02)*S13+0.000000e+00*S14+0.000000e+00*S15+(-2.627679e+01)*S16+1.561365e+01*S17+0.000000e+00*S18+0.000000e+00*S19 \
V24_part3=V24_part2+1.495444e+02*S20+(-1.120318e+02)*S21+(-1.471098e+02)*S22+1.006927e+02*S23+0.000000e+00*S24+0.000000e+00*S25+(-2.626714e+02)*S26+(-9.915910e+01)*S27+0.000000e+00*S28+6.469577e+01*S29 \
V24=V24_part3+(-3.472751e+03)*S30+0.000000e+00*S31+2.336341e+02*S32+(-6.189568e+02)*S33+0.000000e+00*S34+0.000000e+00*S35+4.912425e+02*S36 \
V25_part1=3.184610e+01*S0+0.000000e+00*S1+7.429615e+02*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+2.373825e+01*S6+2.914266e+01*S7+2.839173e+01*S8+3.187711e+01*S9 \
V25_part2=V25_part1+0.000000e+00*S10+1.586759e+03*S11+5.470479e+02*S12+2.162736e+03*S13+0.000000e+00*S14+0.000000e+00*S15+1.076273e+02*S16+5.806951e+02*S17+0.000000e+00*S18+0.000000e+00*S19 \
V25_part3=V25_part2+(-4.285948e+01)*S20+7.698605e+02*S21+7.601704e+02*S22+2.304709e+02*S23+0.000000e+00*S24+0.000000e+00*S25+6.999643e+02*S26+7.424581e+02*S27+0.000000e+00*S28+4.235915e+02*S29 \
V25=V25_part3+5.891802e+03*S30+0.000000e+00*S31+4.047335e+02*S32+1.271518e+03*S33+0.000000e+00*S34+0.000000e+00*S35+3.630916e+01*S36 \
V26_part1=2.463342e+01*S0+0.000000e+00*S1+3.365444e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+(-4.612957e+00)*S6+(-5.436564e+00)*S7+1.344959e+00*S8+1.469240e+01*S9 \
V26_part2=V26_part1+0.000000e+00*S10+1.461829e+02*S11+2.269066e+01*S12+3.067936e+01*S13+0.000000e+00*S14+0.000000e+00*S15+(-1.435190e+01)*S16+(-3.220237e+01)*S17+0.000000e+00*S18+0.000000e+00*S19 \
V26_part3=V26_part2+3.284180e+01*S20+1.753480e-01*S21+3.388173e+02*S22+(-5.220491e+01)*S23+0.000000e+00*S24+0.000000e+00*S25+4.503689e+00*S26+(-1.126246e+02)*S27+0.000000e+00*S28+(-1.954619e+01)*S29 \
V26=V26_part3+1.685417e+03*S30+0.000000e+00*S31+(-5.087332e+02)*S32+(-4.354797e+02)*S33+0.000000e+00*S34+0.000000e+00*S35+4.394091e+02*S36 \
V27_part1=(-4.907766e-01)*S0+(-1.416786e+00)*S1+(-1.913161e+00)*S2+(-8.317363e+00)*S3+(-1.670695e+00)*S4+(-2.799643e+01)*S5+(-9.973332e+00)*S6+(-1.154946e+00)*S7+(-1.779006e+01)*S8+(-3.406407e+00)*S9 \
V27_part2=V27_part1+(-1.613930e+00)*S10+(-1.516919e+00)*S11+(-3.339524e+00)*S12+(-2.028725e+00)*S13+(-2.918594e+00)*S14+(-3.061131e-01)*S15+(-2.872921e-01)*S16+(-1.618635e+00)*S17+(-1.865712e+00)*S18+2.964196e+00*S19 \
V27_part3=V27_part2+(-2.027532e+00)*S20+(-1.400339e+00)*S21+(-2.264082e+00)*S22+(-1.610634e+00)*S23+(-1.404242e+00)*S24+(-2.489379e+00)*S25+(-1.189124e+00)*S26+(-2.875907e+00)*S27+(-1.822029e+00)*S28+(-2.346500e+00)*S29 \
V27=V27_part3+(-5.291872e-01)*S30+(-1.598199e+00)*S31+(-1.811318e+00)*S32+(-1.997702e+00)*S33+(-1.730522e+00)*S34+(-2.148906e+00)*S35+(-3.292094e+00)*S36 \
V28_part1=1.345826e+00*S0+1.550261e+00*S1+9.110657e+00*S2+2.059542e+01*S3+6.778732e+00*S4+1.356070e+01*S5+1.647474e+01*S6+2.321505e+01*S7+1.966124e+01*S8+7.977425e+00*S9 \
V28_part2=V28_part1+8.642479e+00*S10+6.212244e+00*S11+1.156010e+01*S12+5.864625e+00*S13+9.001148e+00*S14+1.434180e+00*S15+2.321498e+00*S16+9.521647e+00*S17+9.273163e-01*S18+1.743811e-01*S19 \
V28_part3=V28_part2+1.016107e+01*S20+8.278014e+00*S21+9.097161e+00*S22+9.334735e+00*S23+9.121397e+00*S24+1.087088e+01*S25+5.702061e+00*S26+9.439805e+00*S27+9.833953e+00*S28+9.895596e+00*S29 \
V28=V28_part3+1.216903e+00*S30+1.006340e+01*S31+9.189404e+00*S32+9.259134e+00*S33+9.821300e+00*S34+1.000074e+01*S35+9.573181e+00*S36 \
V29_part1=6.059926e+00*S0+7.873066e+00*S1+5.103809e+00*S2+1.286490e+01*S3+6.762460e+00*S4+9.486666e+01*S5+2.538211e+01*S6+9.323823e+00*S7+3.986367e+01*S8+9.497885e+00*S9 \
V29_part2=V29_part1+8.397823e+00*S10+8.008126e+00*S11+9.544603e+00*S12+9.323635e+00*S13+1.136214e+01*S14+4.273917e+00*S15+5.847381e+00*S16+5.286147e+00*S17+1.390995e+01*S18+6.031328e+00*S19 \
V29_part3=V29_part2+1.101487e+01*S20+1.081955e+01*S21+1.133192e+01*S22+8.278306e+00*S23+6.905375e+00*S24+8.929647e+00*S25+9.008601e+00*S26+1.100088e+01*S27+1.251017e+01*S28+1.301304e+01*S29 \
V29=V29_part3+1.719444e+01*S30+7.967395e+00*S31+1.028180e+01*S32+1.089829e+01*S33+1.198986e+01*S34+1.176730e+01*S35+1.496082e+01*S36 \
V30_part1=1.921147e-01*S0+8.080166e-01*S1+5.052821e-01*S2+4.037982e+03*S3+(-1.313757e-01)*S4+1.014340e+02*S5+1.178312e+02*S6+4.512374e+01*S7+1.355042e+02*S8+6.199962e+01*S9 \
V30_part2=V30_part1+3.593295e-01*S10+2.132304e+00*S11+4.627973e-01*S12+5.147220e+00*S13+(-1.089291e-02)*S14+4.546673e-02*S15+1.811269e+00*S16+9.015618e-01*S17+2.124157e+01*S18+(-4.779342e-01)*S19 \
V30_part3=V30_part2+(-9.788725e-02)*S20+6.511456e+00*S21+1.186118e+00*S22+8.847437e-02*S23+1.626406e-01*S24+(-5.876088e-01)*S25+5.670479e-01*S26+2.633887e-01*S27+3.450568e-01*S28+1.162722e+00*S29 \
V30=V30_part3+1.352868e+00*S30+7.104231e-02*S31+1.908997e-01*S32+1.000000e+04*S33+2.551744e-01*S34+1.022113e+00*S35+1.416331e+01*S36 \
V31_part1=1.297254e+00*S0+6.307078e-01*S1+(-1.015222e-01)*S2+3.905220e+01*S3+(-2.511771e-01)*S4+7.567857e+01*S5+3.478676e+01*S6+1.758640e+02*S7+(-6.608865e+00)*S8+1.930041e+01*S9 \
V31_part2=V31_part1+(-2.302945e-01)*S10+(-5.108907e-01)*S11+(-3.173191e-02)*S12+(-2.191776e+00)*S13+(-2.487653e-01)*S14+6.820714e+00*S15+5.454933e-01*S16+(-8.790911e-02)*S17+2.129571e+00*S18+1.194204e+00*S19 \
V31_part3=V31_part2+(-5.058514e-01)*S20+2.289783e-02*S21+1.186736e-01*S22+(-8.675803e-01)*S23+(-1.926278e-01)*S24+(-4.068525e-01)*S25+(-3.148183e-01)*S26+(-1.292614e-01)*S27+(-4.107680e-01)*S28+9.977752e-01*S29 \
V31=V31_part3+(-7.700674e-01)*S30+(-2.440281e-02)*S31+2.564307e-01*S32+1.000000e+04*S33+(-8.194695e-01)*S34+9.176249e-01*S35+6.840586e-01*S36 \
V32_part1=(-3.521929e-01)*S0+(-6.062316e-01)*S1+(-3.294175e-03)*S2+(-5.026926e+03)*S3+1.239291e+00*S4+(-7.339912e+01)*S5+(-1.211152e+02)*S6+(-5.169713e+01)*S7+(-1.256154e+02)*S8+(-4.786081e+01)*S9 \
V32_part2=V32_part1+1.621439e-01*S10+(-1.947757e+00)*S11+5.658718e-02*S12+(-3.580015e+00)*S13+1.104832e+00*S14+(-9.091701e-01)*S15+(-1.684917e+00)*S16+(-5.009641e-01)*S17+4.250120e-01*S18+4.709118e-01*S19 \
V32_part3=V32_part2+2.021728e+00*S20+(-9.881392e+00)*S21+(-1.369285e+00)*S22+1.676508e+00*S23+7.669074e-01*S24+2.785887e+00*S25+2.725414e-01*S26+4.574314e-01*S27+6.716988e-01*S28+(-2.189088e+00)*S29 \
V32=V32_part3+(-4.218831e-01)*S30+3.879153e-01*S31+8.138608e-01*S32+5.322916e+03*S33+2.006824e+00*S34+(-1.889875e+00)*S35+(-2.643946e+01)*S36 \
V33_part1=(-4.146251e+01)*S0+(-4.007854e+01)*S1+(-1.032521e+02)*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+(-5.079812e+00)*S9 \
V33_part2=V33_part1+2.579271e+01*S10+(-4.216204e+02)*S11+5.709017e+01*S12+(-2.957257e+02)*S13+0.000000e+00*S14+0.000000e+00*S15+(-1.854066e+00)*S16+(-1.478990e+02)*S17+0.000000e+00*S18+0.000000e+00*S19 \
V33_part3=V33_part2+4.631222e+01*S20+(-1.894504e+02)*S21+(-1.041988e+02)*S22+1.028942e+02*S23+(-2.442379e-01)*S24+0.000000e+00*S25+(-3.691279e+02)*S26+(-1.128350e+02)*S27+0.000000e+00*S28+0.000000e+00*S29 \
V33=V33_part3+(-6.276574e+02)*S30+1.900447e+02*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+3.420882e+01*S36 \
V34_part1=1.273665e+02*S0+6.448046e+01*S1+8.186402e+02*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+3.049179e+01*S9 \
V34_part2=V34_part1+2.671002e+02*S10+1.467830e+03*S11+5.037270e+02*S12+1.065054e+03*S13+0.000000e+00*S14+0.000000e+00*S15+1.014817e+02*S16+7.396003e+02*S17+0.000000e+00*S18+0.000000e+00*S19 \
V34_part3=V34_part2+1.530697e+02*S20+1.023470e+03*S21+7.776920e+02*S22+1.184018e+02*S23+4.580011e+02*S24+0.000000e+00*S25+7.823248e+02*S26+6.893211e+02*S27+0.000000e+00*S28+0.000000e+00*S29 \
V34=V34_part3+1.139548e+03*S30+(-9.967858e+01)*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+(-2.194216e+01)*S36 \
V35_part1=2.229082e+02*S0+2.525143e+02*S1+2.778641e+00*S2+0.000000e+00*S3+0.000000e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+8.835403e-01*S9 \
V35_part2=V35_part1+(-5.260696e+01)*S10+1.299066e+02*S11+(-1.457400e+02)*S12+1.273437e+02*S13+0.000000e+00*S14+0.000000e+00*S15+(-3.095445e+01)*S16+1.521095e+02*S17+0.000000e+00*S18+0.000000e+00*S19 \
V35_part3=V35_part2+(-3.594785e+01)*S20+(-6.947368e+01)*S21+(-4.801235e-01)*S22+(-6.017577e+01)*S23+7.339642e+01*S24+0.000000e+00*S25+(-1.487661e+02)*S26+(-1.206327e+02)*S27+0.000000e+00*S28+0.000000e+00*S29 \
V35=V35_part3+9.949639e+02*S30+(-2.882499e+01)*S31+0.000000e+00*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+5.618057e+00*S36 \
V36_part1=(-2.061684e+00)*S0+(-8.362754e-01)*S1+(-2.283160e+00)*S2+(-1.372575e+00)*S3+(-7.830364e+00)*S4+(-1.280722e+00)*S5+(-1.405127e+00)*S6+(-4.047131e+00)*S7+(-1.178621e+00)*S8+(-3.403899e+00)*S9 \
V36_part2=V36_part1+0.000000e+00*S10+(-2.627016e+00)*S11+(-1.756198e+00)*S12+(-3.502260e+00)*S13+(-1.184584e+01)*S14+(-1.806286e+00)*S15+(-3.476001e+00)*S16+(-5.687384e+00)*S17+(-2.675548e+00)*S18+(-1.547486e+01)*S19 \
V36_part3=V36_part2+0.000000e+00*S20+(-6.341264e+00)*S21+(-7.514292e+00)*S22+0.000000e+00*S23+(-4.270579e+00)*S24+(-8.987726e+00)*S25+(-6.874741e+00)*S26+(-1.644585e+01)*S27+(-3.071488e+00)*S28+(-6.074809e+00)*S29 \
V36=V36_part3+(-1.255988e+01)*S30+(-5.438574e+00)*S31+(-5.637102e+00)*S32+(-7.883545e+00)*S33+(-3.575984e+00)*S34+(-7.306876e+00)*S35+(-8.745375e+00)*S36 \
V37_part1=1.130761e+01*S0+8.883288e+00*S1+8.172183e-01*S2+(-1.480129e+00)*S3+5.043052e+00*S4+6.406283e+00*S5+5.259301e+00*S6+7.650503e+00*S7+4.542693e+00*S8+7.475375e+00*S9 \
V37_part2=V37_part1+0.000000e+00*S10+6.017207e+00*S11+2.693843e-01*S12+5.991275e+00*S13+7.379745e+00*S14+1.036246e+01*S15+9.063003e+00*S16+2.670915e+00*S17+1.106842e+01*S18+1.734254e+01*S19 \
V37_part3=V37_part2+0.000000e+00*S20+7.858195e+00*S21+4.395941e+00*S22+0.000000e+00*S23+1.899701e+00*S24+7.625057e+00*S25+7.654149e+00*S26+1.317203e+01*S27+5.806513e+00*S28+7.583737e+00*S29 \
V37=V37_part3+2.222373e+01*S30+6.197019e+00*S31+6.379361e+00*S32+4.050557e+00*S33+6.963254e+00*S34+8.941113e+00*S35+9.607550e+00*S36 \
V38_part1=(-4.623696e-02)*S0+6.331533e-02*S1+4.301664e+00*S2+9.866379e+00*S3+7.504428e+00*S4+6.298961e+00*S5+7.425044e+00*S6+7.978933e+00*S7+7.556285e+00*S8+6.733021e+00*S9 \
V38_part2=V38_part1+0.000000e+00*S10+6.364392e+00*S11+4.425345e+00*S12+1.109392e+01*S13+1.166302e+01*S14+4.135528e+00*S15+5.601277e+00*S16+8.096676e+00*S17+(-2.042886e+00)*S18+1.112613e+01*S19 \
V38_part3=V38_part2+0.000000e+00*S20+9.922035e+00*S21+1.881337e+01*S22+0.000000e+00*S23+1.173948e+01*S24+1.125652e+01*S25+1.507553e+01*S26+1.536889e+01*S27+7.727631e+00*S28+1.539674e+01*S29 \
V38=V38_part3+1.844839e+01*S30+2.938158e+01*S31+1.329992e+01*S32+2.494842e+01*S33+9.866465e+00*S34+2.044654e+01*S35+2.487261e+01*S36 \
V39_part1=0.000000e+00*S0+0.000000e+00*S1+(-5.471594e-01)*S2+2.034005e-02*S3+0.000000e+00*S4+2.158858e-02*S5+1.714407e-02*S6+2.458605e-02*S7+0.000000e+00*S8+1.823278e-03*S9 \
V39_part2=V39_part1+(-8.021978e-02)*S10+(-5.002396e-01)*S11+(-6.413453e-02)*S12+3.889892e+00*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+1.028572e-02*S17+0.000000e+00*S18+0.000000e+00*S19 \
V39_part3=V39_part2+0.000000e+00*S20+(-1.701494e-01)*S21+(-2.061171e-01)*S22+1.133085e+00*S23+6.596759e-01*S24+(-1.799628e-01)*S25+9.612874e+00*S26+1.004453e+01*S27+8.011002e-02*S28+(-1.758201e-02)*S29 \
V39=V39_part3+(-5.549608e+00)*S30+(-1.680640e+03)*S31+0.000000e+00*S32+2.693170e-01*S33+1.896699e-01*S34+(-1.945441e-01)*S35+3.094709e-01*S36 \
V40_part1=0.000000e+00*S0+0.000000e+00*S1+2.550041e+00*S2+(-3.144428e-02)*S3+0.000000e+00*S4+(-1.307085e-02)*S5+(-8.512993e-03)*S6+(-1.541154e-02)*S7+0.000000e+00*S8+1.509380e-02*S9 \
V40_part2=V40_part1+(-1.738703e-01)*S10+2.433931e+00*S11+(-1.999941e-02)*S12+1.786558e+00*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+(-3.885510e-01)*S17+0.000000e+00*S18+0.000000e+00*S19 \
V40_part3=V40_part2+0.000000e+00*S20+4.493598e-01*S21+(-1.405065e-01)*S22+2.002920e+00*S23+9.169274e-01*S24+2.588973e-01*S25+6.155600e-01*S26+1.371214e+00*S27+2.094974e+00*S28+(-4.237010e-01)*S29 \
V40=V40_part3+6.277860e+00*S30+1.000000e+04*S31+0.000000e+00*S32+(-1.219109e-01)*S33+8.407348e-01*S34+(-7.510748e-01)*S35+(-2.806951e-01)*S36 \
V41_part1=0.000000e+00*S0+0.000000e+00*S1+(-2.559034e-01)*S2+1.479411e-01*S3+0.000000e+00*S4+2.521794e-02*S5+1.035783e-02*S6+2.891988e-02*S7+0.000000e+00*S8+2.739178e-02*S9 \
V41_part2=V41_part1+9.113120e-01*S10+(-1.492443e-01)*S11+5.511272e-01*S12+(-5.753022e+00)*S13+0.000000e+00*S14+0.000000e+00*S15+0.000000e+00*S16+1.041740e+00*S17+0.000000e+00*S18+0.000000e+00*S19 \
V41_part3=V41_part2+0.000000e+00*S20+1.998567e-01*S21+1.623985e+00*S22+(-1.919531e+00)*S23+(-1.087145e+00)*S24+1.504778e-01*S25+(-1.215004e+01)*S26+(-1.091882e+01)*S27+(-6.626048e-01)*S28+2.074739e+00*S29 \
V41=V41_part3+6.285481e+00*S30+1.365430e+02*S31+0.000000e+00*S32+3.427903e-02*S33+(-3.586405e-01)*S34+3.684692e+00*S35+3.718300e-01*S36 \
V42_part1=0.000000e+00*S0+8.748653e+03*S1+0.000000e+00*S2+3.244148e+02*S3+0.000000e+00*S4+2.986493e+03*S5+0.000000e+00*S6+2.040513e+02*S7+9.803207e+02*S8+0.000000e+00*S9 \
V42_part2=V42_part1+6.772774e+02*S10+0.000000e+00*S11+1.601227e+03*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+4.873814e-01*S16+0.000000e+00*S17+3.723532e+03*S18+0.000000e+00*S19 \
V42_part3=V42_part2+1.736003e+03*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+(-4.167481e+01)*S24+2.516046e+03*S25+1.275568e+03*S26+9.579891e+02*S27+6.651936e+02*S28+(-3.578615e+01)*S29 \
V42=V42_part3+0.000000e+00*S30+(-2.897087e+01)*S31+0.000000e+00*S32+3.735068e+02*S33+0.000000e+00*S34+(-3.339961e+01)*S35+(-1.859816e+02)*S36 \
V43_part1=0.000000e+00*S0+(-1.205859e+02)*S1+0.000000e+00*S2+7.817777e+02*S3+0.000000e+00*S4+(-2.272111e+03)*S5+0.000000e+00*S6+1.158123e+03*S7+6.861187e+02*S8+0.000000e+00*S9 \
V43_part2=V43_part1+(-8.923262e+02)*S10+0.000000e+00*S11+(-1.559763e+03)*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+2.310868e+01*S16+0.000000e+00*S17+4.982709e+03*S18+0.000000e+00*S19 \
V43_part3=V43_part2+1.696099e+02*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+6.543535e+02*S24+1.330919e+02*S25+(-6.740187e+02)*S26+(-7.163746e+02)*S27+(-5.286072e+02)*S28+9.499082e+02*S29 \
V43=V43_part3+0.000000e+00*S30+4.157829e+01*S31+0.000000e+00*S32+(-1.526472e+02)*S33+0.000000e+00*S34+1.280251e+03*S35+2.139525e+02*S36 \
V44_part1=0.000000e+00*S0+(-3.219348e+03)*S1+0.000000e+00*S2+6.223837e+02*S3+0.000000e+00*S4+(-2.782881e+03)*S5+0.000000e+00*S6+(-2.810931e+02)*S7+(-2.275523e+03)*S8+0.000000e+00*S9 \
V44_part2=V44_part1+2.383571e+02*S10+0.000000e+00*S11+(-3.229664e+02)*S12+0.000000e+00*S13+0.000000e+00*S14+0.000000e+00*S15+(-3.669428e+00)*S16+0.000000e+00*S17+(-1.000000e+04)*S18+0.000000e+00*S19 \
V44_part3=V44_part2+7.295041e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+5.283056e+01*S24+(-1.919737e+03)*S25+(-3.050420e+01)*S26+1.157012e+02*S27+(-5.051938e+01)*S28+(-3.645669e+01)*S29 \
V44=V44_part3+0.000000e+00*S30+1.141503e+02*S31+0.000000e+00*S32+1.377200e+03*S33+0.000000e+00*S34+(-3.799838e+01)*S35+2.636527e+02*S36 \
V45_part1=1.000000e+04*S0+1.000000e+04*S1+1.000000e+04*S2+1.843085e+01*S3+1.000000e+04*S4+2.478665e+01*S5+1.913893e+01*S6+2.372327e+01*S7+1.771945e+01*S8+1.250153e+01*S9 \
V45_part2=V45_part1+1.000000e+04*S10+(-7.338417e-01)*S11+1.000000e+04*S12+(-9.420890e-02)*S13+3.023296e+03*S14+5.637035e+03*S15+1.825683e+00*S16+1.000000e+04*S17+1.000000e+04*S18+1.000000e+04*S19 \
V45_part3=V45_part2+4.781103e+03*S20+3.472444e+02*S21+1.000000e+04*S22+1.000000e+04*S23+2.027957e-01*S24+1.000000e+04*S25+(-8.367960e+01)*S26+(-4.787067e+02)*S27+3.598011e+02*S28+(-1.601326e-02)*S29 \
V45=V45_part3+1.000000e+04*S30+(-6.794786e+01)*S31+3.584362e-01*S32+5.317364e-01*S33+1.000000e+04*S34+1.748198e-01*S35+1.661911e+01*S36 \
V46_part1=1.000000e+04*S0+5.259215e+03*S1+1.000000e+04*S2+2.441735e+01*S3+1.000000e+04*S4+3.037686e+00*S5+2.925026e+00*S6+3.076312e-01*S7+3.120172e+00*S8+8.635582e-01*S9 \
V46_part2=V46_part1+1.000000e+04*S10+(-1.908664e+00)*S11+1.000000e+04*S12+(-7.986076e-01)*S13+1.617113e+01*S14+(-1.000000e+04)*S15+(-7.382987e-01)*S16+1.000000e+04*S17+1.000000e+04*S18+1.000000e+04*S19 \
V46_part3=V46_part2+5.319043e+03*S20+3.472444e+02*S21+(-1.026629e+03)*S22+5.539315e+03*S23+(-2.991360e-01)*S24+1.000000e+04*S25+(-1.290638e+00)*S26+(-2.205145e-01)*S27+4.437944e+00*S28+(-1.150206e+00)*S29 \
V46=V46_part3+1.000000e+04*S30+6.326434e+02*S31+(-1.470117e+00)*S32+8.665323e-01*S33+1.000000e+04*S34+(-4.527656e-01)*S35+(-1.971763e+01)*S36 \
V47_part1=1.000000e+04*S0+1.000000e+04*S1+1.000000e+04*S2+(-2.224044e+01)*S3+1.000000e+04*S4+(-4.364945e+00)*S5+(-1.917575e+00)*S6+(-8.883997e+00)*S7+1.407026e-01*S8+(-2.520060e-01)*S9 \
V47_part2=V47_part1+1.000000e+04*S10+6.956734e+00*S11+1.000000e+04*S12+3.074218e+00*S13+(-2.863730e+02)*S14+(-1.410071e+01)*S15+6.141329e+01*S16+1.000000e+04*S17+1.000000e+04*S18+1.000000e+04*S19 \
V47_part3=V47_part2+1.000000e+04*S20+4.861222e+02*S21+(-1.050932e+02)*S22+1.000000e+04*S23+3.380071e-01*S24+1.000000e+04*S25+2.561200e+02*S26+1.197913e+03*S27+(-3.102281e+00)*S28+2.835180e+00*S29 \
V47=V47_part3+9.895944e+03*S30+1.993983e+02*S31+2.662421e+00*S32+(-1.518950e+00)*S33+(-4.105377e+03)*S34+6.884249e-01*S35+9.504105e+00*S36 \
V48_part1=(-9.435244e-02)*S0+0.000000e+00*S1+0.000000e+00*S2+0.000000e+00*S3+(-1.287048e+00)*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V48_part2=V48_part1+0.000000e+00*S10+0.000000e+00*S11+(-1.748030e-01)*S12+0.000000e+00*S13+(-2.457217e+00)*S14+(-1.975355e-01)*S15+2.311028e-02*S16+9.868242e-02*S17+0.000000e+00*S18+1.880615e-01*S19 \
V48_part3=V48_part2+(-1.988390e+00)*S20+(-2.382366e-01)*S21+0.000000e+00*S22+(-9.312159e-01)*S23+0.000000e+00*S24+1.698282e+00*S25+0.000000e+00*S26+1.785969e+00*S27+0.000000e+00*S28+(-1.890448e+00)*S29 \
V48=V48_part3+0.000000e+00*S30+(-2.549410e-01)*S31+(-1.298235e+00)*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+(-1.098144e+02)*S36 \
V49_part1=4.660224e-01*S0+0.000000e+00*S1+0.000000e+00*S2+0.000000e+00*S3+1.629664e+00*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V49_part2=V49_part1+0.000000e+00*S10+0.000000e+00*S11+8.343175e-02*S12+0.000000e+00*S13+6.352435e+00*S14+2.872495e-01*S15+2.975944e-01*S16+2.376824e+00*S17+0.000000e+00*S18+(-3.041365e-01)*S19 \
V49_part3=V49_part2+1.214013e+01*S20+7.876352e+00*S21+0.000000e+00*S22+7.043262e+00*S23+0.000000e+00*S24+2.796612e-01*S25+0.000000e+00*S26+2.646033e+00*S27+0.000000e+00*S28+1.909588e+01*S29 \
V49=V49_part3+0.000000e+00*S30+1.706578e+00*S31+1.249985e+01*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+3.440019e+02*S36 \
V50_part1=(-4.843345e-02)*S0+0.000000e+00*S1+0.000000e+00*S2+0.000000e+00*S3+7.425505e-01*S4+0.000000e+00*S5+0.000000e+00*S6+0.000000e+00*S7+0.000000e+00*S8+0.000000e+00*S9 \
V50_part2=V50_part1+0.000000e+00*S10+0.000000e+00*S11+4.952255e-01*S12+0.000000e+00*S13+7.596755e-01*S14+5.982515e-01*S15+3.118543e-01*S16+(-1.523119e-01)*S17+0.000000e+00*S18+8.846338e-01*S19 \
V50_part3=V50_part2+1.615769e+00*S20+(-1.650702e-01)*S21+0.000000e+00*S22+1.514866e+00*S23+0.000000e+00*S24+(-5.811191e-01)*S25+0.000000e+00*S26+(-5.501870e-01)*S27+0.000000e+00*S28+(-4.450929e+00)*S29 \
V50=V50_part3+0.000000e+00*S30+1.188969e+00*S31+(-1.505801e+00)*S32+0.000000e+00*S33+0.000000e+00*S34+0.000000e+00*S35+(-1.361615e+01)*S36 \
V51_part1=(-1.846268e+01)*S0+(-1.801214e+01)*S1+1.000000e+04*S2+8.029359e+03*S3+1.000000e+04*S4+(-8.028947e+02)*S5+1.843948e+03*S6+(-8.498657e+02)*S7+4.520405e+03*S8+(-1.545015e+02)*S9 \
V51_part2=V51_part1+1.000000e+04*S10+1.861715e+00*S11+1.000000e+04*S12+2.998523e+00*S13+3.876471e+00*S14+(-5.327085e+01)*S15+1.761270e+00*S16+1.000000e+04*S17+(-1.712885e+01)*S18+(-1.082185e+00)*S19 \
V51_part3=V51_part2+(-4.671337e+00)*S20+2.591960e-03*S21+1.696560e-01*S22+1.000000e+04*S23+0.000000e+00*S24+(-1.461236e+02)*S25+3.266248e+00*S26+1.945250e+02*S27+7.280348e-01*S28+3.818328e+03*S29 \
V51=V51_part3+3.268545e+00*S30+9.417760e+00*S31+(-4.339835e-02)*S32+4.576351e+00*S33+7.285898e+03*S34+1.000000e+04*S35+5.981163e+00*S36 \
V52_part1=(-4.483473e+00)*S0+(-3.626141e+00)*S1+1.000000e+04*S2+5.280795e+01*S3+1.000000e+04*S4+6.099404e+03*S5+1.000000e+04*S6+3.774542e+03*S7+6.506036e+03*S8+9.479047e+03*S9 \
V52_part2=V52_part1+1.000000e+04*S10+(-6.790355e+00)*S11+1.000000e+04*S12+(-1.656216e+00)*S13+(-8.289130e-01)*S14+(-4.168467e+02)*S15+(-9.053643e+01)*S16+1.000000e+04*S17+2.746496e+00*S18+1.463431e-01*S19 \
V52_part3=V52_part2+(-2.198022e+01)*S20+(-1.110957e+00)*S21+(-1.517796e-01)*S22+9.316204e+03*S23+0.000000e+00*S24+(-1.124584e+00)*S25+1.232872e+02*S26+3.687271e+00*S27+9.180128e+02*S28+8.918742e+00*S29 \
V52=V52_part3+1.300109e-01*S30+3.025543e+01*S31+(-4.081685e-01)*S32+(-4.458676e+00)*S33+7.285898e+03*S34+1.000000e+04*S35+1.502795e+02*S36 \
V53_part1=6.699149e+01*S0+7.146223e+01*S1+1.000000e+04*S2+(-1.000000e+04)*S3+1.000000e+04*S4+(-1.153220e+03)*S5+3.682463e+03*S6+(-3.455782e+02)*S7+(-1.000000e+04)*S8+(-6.210460e+03)*S9 \
V53_part2=V53_part1+1.000000e+04*S10+1.820951e+01*S11+1.000000e+04*S12+(-8.574348e-01)*S13+(-1.955740e+00)*S14+7.275498e+02*S15+1.938538e+02*S16+1.000000e+04*S17+5.471442e+01*S18+3.406417e+00*S19 \
V53_part3=V53_part2+4.611664e+01*S20+2.619868e+00*S21+(-5.594097e-02)*S22+1.000000e+04*S23+0.000000e+00*S24+3.679375e+02*S25+(-9.046212e+01)*S26+(-1.806569e+02)*S27+1.807730e+01*S28+4.272753e+02*S29 \
V53=V53_part3+(-5.113383e+00)*S30+(-1.683329e+01)*S31+2.518076e+00*S32+1.139841e-01*S33+(-2.595258e+03)*S34+3.460806e+03*S35+1.231576e+01*S36 \
V54_part1=(-4.200138e-01)*S0+(-4.426629e-01)*S1+0.000000e+00*S2+(-3.495701e-01)*S3+1.850109e+00*S4+2.288497e-04*S5+0.000000e+00*S6+2.243959e-02*S7+0.000000e+00*S8+0.000000e+00*S9 \
V54_part2=V54_part1+(-1.803077e+00)*S10+2.569117e+00*S11+(-1.893049e+00)*S12+(-2.042207e+00)*S13+2.903107e+00*S14+3.802131e-01*S15+1.018092e+00*S16+0.000000e+00*S17+(-1.199848e+00)*S18+4.945736e+00*S19 \
V54_part3=V54_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+(-2.390301e+00)*S25+3.969294e+00*S26+0.000000e+00*S27+(-1.251130e+00)*S28+0.000000e+00*S29 \
V54=V54_part3+8.245426e+00*S30+0.000000e+00*S31+0.000000e+00*S32+(-6.574870e+00)*S33+(-7.458432e-02)*S34+0.000000e+00*S35+7.616648e+01*S36 \
V55_part1=9.104523e-01*S0+6.048455e-01*S1+0.000000e+00*S2+1.090376e+00*S3+5.710490e+00*S4+2.226341e-01*S5+0.000000e+00*S6+3.695050e-02*S7+0.000000e+00*S8+0.000000e+00*S9 \
V55_part2=V55_part1+1.859484e+01*S10+(-2.859857e+00)*S11+1.024818e+01*S12+3.332762e+00*S13+4.286990e+00*S14+2.475983e-02*S15+6.970494e-02*S16+0.000000e+00*S17+1.104657e+00*S18+(-6.332224e-01)*S19 \
V55_part3=V55_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+1.081505e+01*S25+2.018173e+00*S26+0.000000e+00*S27+2.589118e+01*S28+0.000000e+00*S29 \
V55=V55_part3+7.200680e+00*S30+0.000000e+00*S31+0.000000e+00*S32+2.077853e+01*S33+2.056130e+01*S34+0.000000e+00*S35+(-3.002118e+01)*S36 \
V56_part1=1.776604e+00*S0+2.348537e+00*S1+0.000000e+00*S2+4.759139e-01*S3+(-2.468723e+00)*S4+(-8.243522e-02)*S5+0.000000e+00*S6+4.689853e-02*S7+0.000000e+00*S8+0.000000e+00*S9 \
V56_part2=V56_part1+1.726904e+00*S10+(-1.473227e-01)*S11+2.268353e+00*S12+2.301456e+00*S13+(-2.166710e+00)*S14+2.455002e-01*S15+1.564877e-01*S16+0.000000e+00*S17+6.348913e+00*S18+(-2.254053e+00)*S19 \
V56_part3=V56_part2+0.000000e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+7.405348e-01*S25+(-3.830314e+00)*S26+0.000000e+00*S27+(-4.369668e-01)*S28+0.000000e+00*S29 \
V56=V56_part3+(-1.691514e+01)*S30+0.000000e+00*S31+0.000000e+00*S32+1.504145e+01*S33+(-1.267894e+00)*S34+0.000000e+00*S35+(-7.736725e+01)*S36 \
V57_part1=4.004720e+03*S0+9.999176e+03*S1+(-1.606258e+00)*S2+(-4.317310e+01)*S3+1.830649e+00*S4+(-1.414170e+03)*S5+9.253100e+03*S6+(-9.216679e+02)*S7+9.913172e+03*S8+8.122543e+03*S9 \
V57_part2=V57_part1+(-3.331052e+03)*S10+(-1.649933e+03)*S11+(-3.828002e+03)*S12+2.156012e+03*S13+3.664295e+00*S14+5.274827e+00*S15+(-1.741243e+00)*S16+0.000000e+00*S17+9.561906e-01*S18+(-3.402730e+00)*S19 \
V57_part3=V57_part2+1.218184e+00*S20+3.161260e-01*S21+1.032459e-02*S22+0.000000e+00*S23+3.205245e+02*S24+1.840104e+00*S25+(-3.065351e+00)*S26+(-1.120450e+02)*S27+1.549465e+01*S28+0.000000e+00*S29 \
V57=V57_part3+5.494080e+03*S30+1.500533e+02*S31+(-3.146610e+00)*S32+2.956357e+03*S33+1.305973e+01*S34+0.000000e+00*S35+2.993397e+00*S36 \
V58_part1=3.082828e+03*S0+8.094366e+03*S1+(-2.546244e+01)*S2+1.026692e+02*S3+(-6.236833e-01)*S4+1.000000e+04*S5+9.247851e+03*S6+9.316326e+03*S7+2.027205e+02*S8+1.688325e+03*S9 \
V58_part2=V58_part1+(-4.987214e+00)*S10+(-1.226926e+03)*S11+(-5.126017e+01)*S12+7.994346e+02*S13+(-3.759595e-01)*S14+(-7.268016e+00)*S15+(-6.201343e-02)*S16+0.000000e+00*S17+7.520931e-02*S18+(-7.578809e-01)*S19 \
V58_part3=V58_part2+8.209430e-01*S20+(-6.513450e-01)*S21+(-1.164389e-01)*S22+0.000000e+00*S23+9.636335e+02*S24+(-4.778241e-01)*S25+3.691296e+02*S26+1.421238e+03*S27+3.043770e+01*S28+0.000000e+00*S29 \
V58=V58_part3+(-7.114478e+03)*S30+1.221370e+02*S31+(-1.855377e+00)*S32+(-2.954439e+03)*S33+(-1.021629e+00)*S34+0.000000e+00*S35+(-2.605195e+00)*S36 \
V59_part1=1.000000e+04*S0+1.000000e+04*S1+3.982935e+01*S2+7.549593e+00*S3+(-6.436671e-01)*S4+(-1.739018e+03)*S5+(-7.591160e+03)*S6+2.312215e+03*S7+(-8.081858e+03)*S8+(-7.524834e+03)*S9 \
V59_part2=V59_part1+1.000000e+04*S10+8.557476e+03*S11+9.752606e+03*S12+(-2.577634e+03)*S13+(-2.184993e+00)*S14+2.722488e-02*S15+7.298070e+00*S16+0.000000e+00*S17+(-5.401968e-01)*S18+1.123378e+01*S19 \
V59_part3=V59_part2+(-1.652495e+00)*S20+6.294154e-01*S21+4.020307e-01*S22+0.000000e+00*S23+1.662101e+02*S24+(-8.676561e-01)*S25+(-2.554181e+02)*S26+(-8.576211e+02)*S27+1.584353e+03*S28+0.000000e+00*S29 \
V59=V59_part3+5.388038e+03*S30+2.532905e+03*S31+1.940995e+01*S32+(-2.990705e+00)*S33+(-2.189395e+01)*S34+0.000000e+00*S35+3.940037e-01*S36 \
V60_part1=0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+(-1.268048e-01)*S3+1.167351e+00*S4+(-2.743252e-03)*S5+(-1.277520e-02)*S6+(-1.034683e-02)*S7+(-8.135445e-02)*S8+(-6.017969e-02)*S9 \
V60_part2=V60_part1+(-9.351939e-01)*S10+2.155392e+00*S11+(-3.746837e+00)*S12+0.000000e+00*S13+3.107565e+00*S14+3.840151e-01*S15+7.950417e-01*S16+0.000000e+00*S17+(-1.285700e+00)*S18+4.738439e+00*S19 \
V60_part3=V60_part2+1.199924e+00*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+(-4.234838e+00)*S25+(-5.667031e+00)*S26+0.000000e+00*S27+(-1.081660e+00)*S28+0.000000e+00*S29 \
V60=V60_part3+0.000000e+00*S30+0.000000e+00*S31+5.000521e-01*S32+(-1.065983e+01)*S33+(-2.501007e+00)*S34+0.000000e+00*S35+0.000000e+00*S36 \
V61_part1=0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+1.132099e+00*S3+6.826562e+00*S4+2.347120e-01*S5+2.484211e-01*S6+3.330280e-01*S7+3.035998e-01*S8+1.697019e-02*S9 \
V61_part2=V61_part1+8.188970e+00*S10+(-2.099477e+00)*S11+9.286864e+00*S12+0.000000e+00*S13+3.851418e+00*S14+1.197330e-02*S15+2.089905e-02*S16+0.000000e+00*S17+1.007450e+00*S18+(-6.414786e-01)*S19 \
V61_part3=V61_part2+(-2.463848e+00)*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+1.282044e+01*S25+1.034210e+01*S26+0.000000e+00*S27+2.342274e+01*S28+0.000000e+00*S29 \
V61=V61_part3+0.000000e+00*S30+0.000000e+00*S31+2.920546e+00*S32+3.928789e+01*S33+2.322065e+01*S34+0.000000e+00*S35+0.000000e+00*S36 \
V62_part1=0.000000e+00*S0+0.000000e+00*S1+0.000000e+00*S2+5.154937e-01*S3+(-1.975579e+00)*S4+(-3.409442e-02)*S5+(-1.308381e-02)*S6+1.939379e-02*S7+4.835651e-02*S8+2.013896e-01*S9 \
V62_part2=V62_part1+2.552550e+00*S10+(-3.902051e-01)*S11+3.608417e+00*S12+0.000000e+00*S13+(-1.939739e+00)*S14+2.356758e-01*S15+3.937623e-01*S16+0.000000e+00*S17+6.902282e+00*S18+(-2.171540e+00)*S19 \
V62_part3=V62_part2+6.453709e-01*S20+0.000000e+00*S21+0.000000e+00*S22+0.000000e+00*S23+0.000000e+00*S24+1.930498e+00*S25+9.341119e+00*S26+0.000000e+00*S27+(-1.695156e-02)*S28+0.000000e+00*S29 \
V62=V62_part3+0.000000e+00*S30+0.000000e+00*S31+(-8.604619e-01)*S32+(-1.064561e+01)*S33+2.570867e+00*S34+0.000000e+00*S35+0.000000e+00*S36 \
_P0=V0+V1*radius_+V2*w_ \
_P1=0.5*(_P0+sqrt(_P0*_P0+0.001)) \
_P2=1e-15*_P1 \
_P3=V3+V4*radius_+V5/w_ \
_P4=0.5*(_P3+sqrt(_P3*_P3+0.001)) \
_P5=V6+V7*radius_+V8*w_ \
_P6=0.5*(_P5+sqrt(_P5*_P5+0.001)) \
_P7=1e-09*_P6 \
_P8=1e-09*_P6 \
_P9=V9+V10*radius_+V11/w_ \
_P10=0.5*(_P9+sqrt(_P9*_P9+0.001)) \
_P11=V12+V13*radius_+V14*w_ \
_P12=0.5*(_P11+sqrt(_P11*_P11+0.001)) \
_P13=1e-09*_P12 \
_P14=V15+V16*radius_+V17*w_ \
_P15=0.5*(atan(2*_P14)/1.5708+1) \
_P16=0.7064*_P15 \
_P17=0.7064*_P15 \
_P18=V18+V19*radius_+V20*w_ \
_P19=0.5*(_P18+sqrt(_P18*_P18+0.001)) \
_P20=V21+V22*radius_+V23*w_ \
_P21=0.5*(_P20+sqrt(_P20*_P20+0.001)) \
_P22=V24+V25*radius_+V26*w_ \
_P23=0.5*(_P22+sqrt(_P22*_P22+0.001)) \
_P24=V27+V28*radius_+V29*w_ \
_P25=0.5*(_P24+sqrt(_P24*_P24+0.001)) \
_P26=V30+V31*radius_+V32*w_ \
_P27=0.5*(_P26+sqrt(_P26*_P26+0.001)) \
_P28=V33+V34*radius_+V35*w_ \
_P29=0.5*(_P28+sqrt(_P28*_P28+0.001)) \
_P30=V36+V37*radius_+V38*w_ \
_P31=0.5*(_P30+sqrt(_P30*_P30+0.001)) \
_P32=V39+V40*radius_+V41*w_ \
_P33=0.5*(_P32+sqrt(_P32*_P32+0.001)) \
_P34=V42+V43*radius_+V44*w_ \
_P35=0.5*(_P34+sqrt(_P34*_P34+0.001)) \
_P36=1e-14*_P19 \
_P37=100*_P21 \
_P38=1e-15*_P23 \
_P39=1e-14*_P25 \
_P40=100*_P27 \
_P41=1e-15*_P29 \
_P42=1e-14*_P31 \
_P43=100*_P33 \
_P44=1e-15*_P35 \
_P45=V45+V46*radius_+V47*w_ \
_P46=0.5*(_P45+sqrt(_P45*_P45+0.001)) \
_P47=V48+V49*radius_+V50*w_ \
_P48=0.5*(_P47+sqrt(_P47*_P47+0.001)) \
_P49=100*_P46 \
_P50=1e-13*_P48 \
_P51=V51+V52*radius_+V53*w_ \
_P52=0.5*(_P51+sqrt(_P51*_P51+0.001)) \
_P53=V54+V55*radius_+V56*w_ \
_P54=0.5*(_P53+sqrt(_P53*_P53+0.001)) \
_P55=100*_P52 \
_P56=1e-13*_P54 \
_P57=V57+V58*radius_+V59*w_ \
_P58=0.5*(_P57+sqrt(_P57*_P57+0.001)) \
_P59=V60+V61*radius_+V62*w_ \
_P60=0.5*(_P59+sqrt(_P59*_P59+0.001)) \
_P61=100*_P58 \
_P62=1e-13*_P60
cs (PLUS MINUS) capacitor c=_P2
rs1_1 (PLUS n1_1) resistor r=_P4*(1+drs_rf_pgs_n) tc1=0.003
ls1_1 (n1_1 ni_1) inductor l=_P7*(1+dls_rf_pgs_n)
rs2_1 (ni_1 n2_1) resistor r=_P4*(1+drs_rf_pgs_n) tc1=0.003
ls2_1 (n2_1 MINUS) inductor l=_P8*(1+dls_rf_pgs_n)
rs1_2 (PLUS n1_2) resistor r=_P10*(1+drs_rf_pgs_n) tc1=0.003
ls1_2 (n1_2 MINUS) inductor l=_P13*(1+dls_rf_pgs_n)
k1 mutual_inductor coupling=_P16 ind1=ls1_1 ind2=ls1_2
k2 mutual_inductor coupling=_P17 ind1=ls2_1 ind2=ls1_2
c_1_sub (PLUS _n1_1_sub) capacitor c=_P36
rs_1_sub (_n1_1_sub 0) resistor r=_P37
cs_1_sub (_n1_1_sub 0) capacitor c=_P38
c_2_sub (MINUS _n1_2_sub) capacitor c=_P39
rs_2_sub (_n1_2_sub 0) resistor r=_P40
cs_2_sub (_n1_2_sub 0) capacitor c=_P41
c_3_sub (ni_1 _n1_3_sub) capacitor c=_P42
rs_3_sub (_n1_3_sub 0) resistor r=_P43
cs_3_sub (_n1_3_sub 0) capacitor c=_P44
rx_1_2_sub (_n1_1_sub _n1_2_sub) resistor r=_P49
cx_1_2_sub (_n1_1_sub _n1_2_sub) capacitor c=_P50
rx_1_3_sub (_n1_1_sub _n1_3_sub) resistor r=_P55
cx_1_3_sub (_n1_1_sub _n1_3_sub) capacitor c=_P56
rx_2_3_sub (_n1_2_sub _n1_3_sub) resistor r=_P61
cx_2_3_sub (_n1_2_sub _n1_3_sub) capacitor c=_P62
ends ind_rf_pgs_n
