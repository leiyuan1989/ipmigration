

*01 Top of hierarchy  cell=an02d0
.subckt an02d0 B A VDD Y GND
M1 N_8 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an02d0

*02 Top of hierarchy  cell=an03d0
.subckt an03d0 C B A GND Y VDD
M1 N_9 A N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.5u m=1
M3 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_2 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 C VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an03d0

*03 Top of hierarchy  cell=an04d0
.subckt an04d0 GND Y VDD D C B A
M1 N_6 A N_4 GND mn5  l=0.5u w=0.58u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.58u m=1
M3 N_8 C N_7 GND mn5  l=0.5u w=0.58u m=1
M4 N_8 D GND GND mn5  l=0.5u w=0.58u m=1
M5 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 C VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 D VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an04d0


*04 Top of hierarchy  cell=an12d0
.subckt an12d0 B AN GND VDD Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_14 N_4 N_2 GND mn5  l=0.5u w=0.5u m=1
M3 N_14 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_2 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an12d0

*05 Top of hierarchy  cell=an13d0
.subckt an13d0 C B AN GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an13d0

*06 Top of hierarchy  cell=an23d0
.subckt an23d0 C BN AN VDD Y GND
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 N_3 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 N_12 C GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_5 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends an23d0

*7 Top of hierarchy  cell=aoi211d0
.subckt aoi211d0 A0 A1 B0 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 Y A1 N_15 GND mn5  l=0.5u w=0.5u m=1
M4 N_15 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M6 N_6 B0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M7 N_6 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi211d0

*11 Top of hierarchy  cell=aoi21d0
.subckt aoi21d0 A0 A1 B0 GND Y VDD
M1 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_12 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y B0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M5 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi21d0

*12 Top of hierarchy  cell=aoi221d0
.subckt aoi221d0 C0 A0 A1 B1 B0 VDD GND Y
M1 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B1 N_12 GND mn5  l=0.5u w=0.5u m=1
M3 N_13 A1 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_13 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y C0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_11 A1 N_7 VDD mp5  l=0.42u w=0.52u m=1
M10 N_11 A0 N_7 VDD mp5  l=0.42u w=0.52u m=1
.ends aoi221d0

*13 Top of hierarchy  cell=aoi22d0
.subckt aoi22d0 B0 B1 A1 A0 GND VDD Y
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 Y B1 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_8 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_8 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 B0 Y VDD mp5  l=0.42u w=0.52u m=1
.ends aoi22d0

*14 Top of hierarchy  cell=aoi31d0
.subckt aoi31d0 A0 A1 A2 B0 VDD Y GND
M1 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A2 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_11 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M6 N_7 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_7 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_7 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi31d0

*15 Top of hierarchy  cell=aoi32d0
.subckt aoi32d0 GND Y VDD A1 A0 A2 B1 B0
M1 N_5 B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B1 N_5 GND mn5  l=0.5u w=0.5u m=1
M3 Y A2 N_7 GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A1 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_6 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_12 B0 Y VDD mp5  l=0.42u w=0.52u m=1
M7 N_12 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_12 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aoi32d0

*16 Top of hierarchy  cell=aoim21d0
.subckt aoim21d0 A1N A0N B0 GND VDD Y
M1 Y B0 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 A0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1N GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 N_13 VDD mp5  l=0.42u w=0.52u m=1
M6 N_13 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_14 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A1N N_14 VDD mp5  l=0.42u w=0.52u m=1
.ends aoim21d0

*17 Top of hierarchy  cell=aoim22d0
.subckt aoim22d0 B1 B0 A1N A0N GND VDD Y
M1 N_2 A0N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_16 B0 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_16 B1 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 A1N N_11 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_10 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends aoim22d0

*18 Top of hierarchy  cell=aor211d0
.subckt aor211d0 C0 B0 A0 A1 GND Y VDD
M1 N_11 A1 N_2 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 C0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 C0 N_18 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor211d0

*19 Top of hierarchy  cell=aor21d0
.subckt aor21d0 B0 A1 A0 VDD Y GND
M1 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 A1 N_10 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor21d0

*20 Top of hierarchy  cell=aor221d0
.subckt aor221d0 GND Y VDD C0 A0 A1 B1 B0
M1 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 B1 N_4 GND mn5  l=0.5u w=0.5u m=1
M4 N_4 A1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_14 A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M8 N_12 A0 N_14 VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_14 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_14 B1 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor221d0

*21 Top of hierarchy  cell=aor22d0
.subckt aor22d0 B0 B1 A1 A0 Y GND VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M4 N_12 B1 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B1 N_9 VDD mp5  l=0.42u w=0.52u m=1
M10 N_9 B0 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends aor22d0


*22 Top of hierarchy  cell=aor311d0
.subckt aor311d0 GND Y VDD A2 A0 A1 B0 C0
M1 N_7 A1 N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_4 C0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A0 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A2 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 B0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_15 C0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M10 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_10 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor311d0


*23 Top of hierarchy  cell=aor31d0
.subckt aor31d0 B0 A2 A1 A0 Y VDD GND
M1 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_2 A2 N_12 GND mn5  l=0.5u w=0.5u m=1
M4 N_2 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_9 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_9 A2 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_2 B0 N_9 VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends aor31d0


*24 Top of hierarchy  cell=buffd0
.subckt buffd0 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends buffd0

*25 Top of hierarchy  cell=buffd1
.subckt buffd1 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.76u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends buffd1


*26 Top of hierarchy  cell=buffd2
.subckt buffd2 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.58u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends buffd2


*27 Top of hierarchy  cell=buffd3
.subckt buffd3 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.74u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.34u m=1
M3 N_4 A GND GND mn5  l=0.5u w=0.58u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.72u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.72u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.76u m=1
.ends buffd3


*28 Top of hierarchy  cell=dfbfb1
.subckt dfbfb1 VDD QN Q GND RN SN CKN D
M1 N_4 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_26 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_27 N_6 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_6 CKN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_23 N_5 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_23 N_10 N_7 GND mn5  l=0.5u w=0.5u m=1
M9 N_23 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_8 N_6 N_28 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_21 SN GND GND mn5  l=0.5u w=0.5u m=1
M15 N_9 N_10 N_21 GND mn5  l=0.5u w=0.5u m=1
M16 N_21 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M18 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M20 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M21 N_4 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_6 N_5 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_4 N_5 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_6 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_16 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_8 N_4 N_17 VDD mp5  l=0.42u w=0.52u m=1
M32 N_18 N_6 N_8 VDD mp5  l=0.42u w=0.5u m=1
M33 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M36 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M37 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M38 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfbfb1


*29 Top of hierarchy  cell=dfcfb1
.subckt dfcfb1 GND QN Q VDD RN D CKN
M1 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_14 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 N_15 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_8 N_4 N_16 GND mn5  l=0.5u w=0.5u m=1
M11 N_17 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_17 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M16 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M18 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M19 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_22 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M23 N_21 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M24 N_22 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M25 N_23 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M27 N_24 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_24 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M29 N_25 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M30 N_25 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M31 N_26 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_26 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M33 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M35 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M36 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends dfcfb1

*30 Top of hierarchy  cell=dfcfq1
.subckt dfcfq1 GND Q VDD CKN D RN
M1 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_16 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M3 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_16 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_15 GND mn5  l=0.5u w=0.5u m=1
M9 N_15 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_14 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_14 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_13 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_25 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_24 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 N_24 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_25 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_23 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_23 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_22 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_22 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_21 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_20 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_21 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_20 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcfq1


*31 Top of hierarchy  cell=dfcrb1
.subckt dfcrb1 VDD QN Q GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_26 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_26 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M9 N_8 N_4 N_25 GND mn5  l=0.5u w=0.5u m=1
M10 N_25 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_24 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_24 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_23 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M16 N_23 D GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M18 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M21 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_19 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M24 N_19 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_18 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_18 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M27 N_17 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_15 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_14 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M33 N_15 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M34 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M35 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrb1


*32 Top of hierarchy  cell=dfcrn1
.subckt dfcrn1 VDD QN GND CK D RN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_10 RN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_34 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_34 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_33 GND mn5  l=0.5u w=0.5u m=1
M8 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_7 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 N_10 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_17 N_10 N_9 VDD mp5  l=0.42u w=0.52u m=1
M20 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_14 N_10 N_7 VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrn1


*33 Top of hierarchy  cell=dfcrq1
.subckt dfcrq1 VDD Q GND CK D RN
M1 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 Q N_3 GND GND mn5  l=0.5u w=0.58u m=1
M4 N_9 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_7 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_33 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_33 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_32 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_32 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_18 N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_17 N_3 N_9 VDD mp5  l=0.42u w=0.52u m=1
M21 N_18 N_3 Q VDD mp5  l=0.42u w=0.76u m=1
M22 N_17 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_14 N_3 N_7 VDD mp5  l=0.42u w=0.52u m=1
M28 N_14 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_4 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfcrq1

*34 Top of hierarchy  cell=dfnfb1
.subckt dfnfb1 VDD QN Q GND D CKN
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_31 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_30 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M10 N_6 N_5 N_28 GND mn5  l=0.5u w=0.5u m=1
M11 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M12 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_15 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M20 N_14 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_13 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M24 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M25 N_12 D VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnfb1

*35 Top of hierarchy  cell=dfnrb1
.subckt dfnrb1 VDD QN Q GND CK D
M1 QN N_10 GND GND mn5  l=0.5u w=0.58u m=1
M2 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_10 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_32 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M6 N_31 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_31 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_30 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_30 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M11 N_6 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M12 N_29 D GND GND mn5  l=0.5u w=0.5u m=1
M13 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M14 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M15 QN N_10 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M17 N_10 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 VDD N_10 N_16 VDD mp5  l=0.42u w=0.5u m=1
M19 N_15 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M20 N_16 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M21 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_14 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M25 N_13 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M26 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dfnrb1

*36 Top of hierarchy  cell=dfnrn1
.subckt dfnrn1 VDD QN GND CK D
M1 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrn1


*37 Top of hierarchy  cell=dfnrq1
.subckt dfnrq1 VDD Q GND CK D
M1 Q N_8 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_9 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_29 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_28 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_28 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_27 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_27 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_6 N_4 N_26 GND mn5  l=0.5u w=0.5u m=1
M10 N_26 D GND GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_4 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M14 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M17 N_14 N_5 N_8 VDD mp5  l=0.42u w=0.5u m=1
M18 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M19 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_12 N_4 N_6 VDD mp5  l=0.42u w=0.5u m=1
M22 N_11 N_5 N_6 VDD mp5  l=0.42u w=0.52u m=1
M23 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_4 N_8 VDD mp5  l=0.42u w=0.52u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_4 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfnrq1


*38 Top of hierarchy  cell=dfpfb1
.subckt dfpfb1 VDD Q QN GND CKN D SN
M1 Q N_11 GND GND mn5  l=0.5u w=0.58u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_11 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_36 N_8 N_9 GND mn5  l=0.5u w=0.5u m=1
M5 N_36 SN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_35 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_35 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M8 N_8 N_4 N_34 GND mn5  l=0.5u w=0.5u m=1
M9 N_34 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_33 SN N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_33 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_32 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_32 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_31 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M15 N_31 D GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M17 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M18 Q N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M19 QN N_9 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_11 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_9 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M22 N_9 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_16 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M24 N_16 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M25 N_15 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M26 N_15 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_7 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_14 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M30 N_13 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M31 N_14 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M32 N_13 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_5 N_4 VDD VDD mp5  l=0.42u w=0.5u m=1
M34 N_4 CKN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfpfb1


*39 Top of hierarchy  cell=dfprb1
.subckt dfprb1 VDD Q QN GND SN D CK
M1 N_4 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_33 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_33 N_12 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_34 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_34 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_10 GND GND mn5  l=0.5u w=0.58u m=1
M7 QN N_8 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_10 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_35 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_35 SN N_6 GND mn5  l=0.5u w=0.5u m=1
M11 N_38 N_7 N_8 GND mn5  l=0.5u w=0.5u m=1
M12 N_36 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M13 N_7 N_4 N_36 GND mn5  l=0.5u w=0.5u m=1
M14 N_37 N_12 N_7 GND mn5  l=0.5u w=0.5u m=1
M15 N_37 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_38 SN GND GND mn5  l=0.5u w=0.5u m=1
M17 N_12 CK GND GND mn5  l=0.5u w=0.5u m=1
M18 N_4 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M19 N_14 D VDD VDD mp5  l=0.42u w=0.52u m=1
M20 N_15 N_12 N_5 VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M22 N_15 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M23 Q N_10 VDD VDD mp5  l=0.42u w=0.76u m=1
M24 QN N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M25 N_10 N_8 VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_6 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_6 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_16 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_12 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_17 N_4 N_7 VDD mp5  l=0.42u w=0.5u m=1
M32 N_17 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M33 N_8 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M34 N_12 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprb1


*40 Top of hierarchy  cell=dfprq1
.subckt dfprq1 VDD Q GND CK D SN
M1 Q N_8 N_27 GND mn5  l=0.5u w=0.58u m=1
M2 N_27 SN GND GND mn5  l=0.5u w=0.58u m=1
M3 N_33 SN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_9 N_8 N_33 GND mn5  l=0.5u w=0.5u m=1
M5 N_32 N_9 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_32 N_5 N_8 GND mn5  l=0.5u w=0.5u m=1
M7 N_8 N_4 N_31 GND mn5  l=0.5u w=0.5u m=1
M8 N_31 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_30 SN GND GND mn5  l=0.5u w=0.5u m=1
M10 N_30 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M11 N_29 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_29 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M14 N_28 D GND GND mn5  l=0.5u w=0.5u m=1
M15 N_4 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M16 N_5 CK GND GND mn5  l=0.5u w=0.5u m=1
M17 Q N_8 VDD VDD mp5  l=0.42u w=0.76u m=1
M18 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M19 N_9 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M20 N_9 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_9 VDD VDD mp5  l=0.42u w=0.5u m=1
M22 N_14 N_4 N_8 VDD mp5  l=0.42u w=0.5u m=1
M23 N_13 N_5 N_8 VDD mp5  l=0.42u w=0.52u m=1
M24 N_13 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M25 N_7 SN VDD VDD mp5  l=0.42u w=0.5u m=1
M26 N_7 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M27 N_12 N_7 VDD VDD mp5  l=0.42u w=0.5u m=1
M28 N_11 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M29 N_12 N_5 N_6 VDD mp5  l=0.42u w=0.5u m=1
M30 N_11 D VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_4 N_5 VDD VDD mp5  l=0.42u w=0.5u m=1
M32 N_5 CK VDD VDD mp5  l=0.42u w=0.5u m=1
.ends dfprq1


*41 Top of hierarchy  cell=dl01d0
.subckt dl01d0 A GND VDD Y
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dl01d0

*42 Top of hierarchy  cell=dl02d0
.subckt dl02d0 A Y VDD GND
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=1u w=0.5u m=1
M3 N_4 N_3 GND GND mn5  l=1u w=0.5u m=1
M4 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_5 N_4 VDD VDD mp5  l=0.84u w=0.52u m=1
M7 N_4 N_3 VDD VDD mp5  l=0.84u w=0.52u m=1
M8 N_3 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends dl02d0


* Top of hierarchy  cell=inv0d0
.subckt inv0d0 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.5u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends inv0d0

* Top of hierarchy  cell=inv0d2
.subckt inv0d2 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d2

* Top of hierarchy  cell=inv0d4
.subckt inv0d4 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d4

* Top of hierarchy  cell=inv0d5
.subckt inv0d5 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.6u m=1
M2 Y A GND GND mn5  l=0.5u w=0.6u m=1
M3 Y A GND GND mn5  l=0.5u w=0.6u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.8u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.8u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.8u m=1
.ends inv0d5

* Top of hierarchy  cell=inv0d6
.subckt inv0d6 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d6

*48 Top of hierarchy  cell=inv0d8
.subckt inv0d8 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A GND GND mn5  l=0.5u w=0.72u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d8

* Top of hierarchy  cell=mi02d0
.subckt mi02d0 VDD Y GND S0 B A
M1 N_4 A GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 N_3 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_5 S0 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 S0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y S0 N_4 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M9 N_5 B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 S0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends mi02d0




* Top of hierarchy  cell=nd02d0
.subckt nd02d0 VDD Y GND B A
M1 Y A N_8 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd02d0


* Top of hierarchy  cell=nd03d0
.subckt nd03d0 C B A Y VDD GND
M1 Y A N_8 GND mn5  l=0.5u w=0.5u m=1
M2 N_9 B N_8 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 C GND GND mn5  l=0.5u w=0.5u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
M5 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd03d0


* Top of hierarchy  cell=nd04d0
.subckt nd04d0 C B D A GND VDD Y
M1 Y A N_9 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B N_9 GND mn5  l=0.5u w=0.5u m=1
M4 N_11 C N_10 GND mn5  l=0.5u w=0.5u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y D VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd04d0


* Top of hierarchy  cell=nd12d0
.subckt nd12d0 B AN Y VDD GND
M1 Y N_4 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd12d0


* Top of hierarchy  cell=nd13d0
.subckt nd13d0 GND Y VDD B C AN
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 B N_6 GND mn5  l=0.5u w=0.5u m=1
M3 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 C GND GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd13d0


* Top of hierarchy  cell=nd14d0
.subckt nd14d0 GND Y VDD B C D AN
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 C N_7 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 B N_6 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y D VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y B VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd14d0


* Top of hierarchy  cell=nd23d0
.subckt nd23d0 AN C BN GND Y VDD
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 N_4 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd23d0

* Top of hierarchy  cell=nd24d0
.subckt nd24d0 GND Y VDD D AN C BN
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_4 N_9 GND mn5  l=0.5u w=0.5u m=1
M3 N_9 N_3 N_8 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 C N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y C VDD VDD mp5  l=0.42u w=0.52u m=1
M11 Y D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nd24d0


* Top of hierarchy  cell=nr02d0
.subckt nr02d0 GND Y VDD B A
M1 Y A GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A VDD VDD mp5  l=0.42u w=0.52u m=1
M4 Y B N_7 VDD mp5  l=0.42u w=0.52u m=1
.ends nr02d0

* Top of hierarchy  cell=nr03d0
.subckt nr03d0 A B C Y VDD GND
M1 Y C GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y A GND GND mn5  l=0.5u w=0.5u m=1
M4 Y C N_8 VDD mp5  l=0.42u w=0.52u m=1
M5 N_9 B N_8 VDD mp5  l=0.42u w=0.52u m=1
M6 N_9 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr03d0

* Top of hierarchy  cell=nr04d0
.subckt nr04d0 A B C D Y VDD GND
M1 Y D GND GND mn5  l=0.5u w=0.5u m=1
M2 Y C GND GND mn5  l=0.5u w=0.5u m=1
M3 Y B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y A GND GND mn5  l=0.5u w=0.5u m=1
M5 Y D N_9 VDD mp5  l=0.42u w=0.52u m=1
M6 N_11 C N_9 VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 B N_10 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr04d0

* Top of hierarchy  cell=nr12d0
.subckt nr12d0 AN B Y VDD GND
M1 Y B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 AN GND GND mn5  l=0.5u w=0.5u m=1
M4 Y B N_8 VDD mp5  l=0.42u w=0.52u m=1
M5 N_8 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr12d0

* Top of hierarchy  cell=nr13d0
.subckt nr13d0 AN B C Y VDD GND
M1 Y C GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_3 AN GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C N_9 VDD mp5  l=0.42u w=0.52u m=1
M6 N_10 B N_9 VDD mp5  l=0.42u w=0.52u m=1
M7 N_10 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_3 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends nr13d0

* Top of hierarchy  cell=nr14d0
.subckt nr14d0 D C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M3 Y B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y C GND GND mn5  l=0.5u w=0.5u m=1
M5 Y D GND GND mn5  l=0.5u w=0.5u m=1
M6 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_16 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M10 Y D N_14 VDD mp5  l=0.42u w=0.52u m=1
.ends nr14d0

* Top of hierarchy  cell=nr23d0
.subckt nr23d0 C AN BN GND VDD Y
M1 N_3 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C GND GND mn5  l=0.5u w=0.5u m=1
M6 N_3 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_11 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_11 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M10 Y C N_10 VDD mp5  l=0.42u w=0.52u m=1
.ends nr23d0

* Top of hierarchy  cell=nr24d0
.subckt nr24d0 D C AN BN Y VDD GND
M1 N_4 BN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y D GND GND mn5  l=0.5u w=0.5u m=1
M7 N_4 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_12 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_13 N_4 N_12 VDD mp5  l=0.42u w=0.52u m=1
M11 N_13 C N_11 VDD mp5  l=0.42u w=0.52u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=0.52u m=1
.ends nr24d0

* Top of hierarchy  cell=oai211d0
.subckt oai211d0 C0 B0 A1 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_9 B0 N_16 GND mn5  l=0.5u w=0.5u m=1
M4 Y C0 N_16 GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 Y A1 N_10 VDD mp5  l=0.42u w=0.52u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai211d0

* Top of hierarchy  cell=oai21d0
.subckt oai21d0 A0 B0 A1 VDD Y GND
M1 N_5 A1 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y B0 N_5 GND mn5  l=0.5u w=0.5u m=1
M3 N_5 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 A1 Y VDD mp5  l=0.42u w=0.52u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_12 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai21d0

* Top of hierarchy  cell=oai221d0
.subckt oai221d0 C0 B1 A1 A0 B0 Y VDD GND
M1 N_7 B0 N_8 GND mn5  l=0.5u w=0.5u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 B1 N_7 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_7 GND mn5  l=0.5u w=0.5u m=1
M6 N_13 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_12 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y A1 N_12 VDD mp5  l=0.42u w=0.52u m=1
M10 N_13 B1 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oai221d0

* Top of hierarchy  cell=oai222d0
.subckt oai222d0 B0 A0 A1 B1 C0 C1 Y VDD GND
M1 N_11 C1 Y GND mn5  l=0.5u w=0.5u m=1
M2 N_11 C0 Y GND mn5  l=0.5u w=0.5u m=1
M3 N_11 B1 N_8 GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_8 B0 N_11 GND mn5  l=0.5u w=0.5u m=1
M7 N_20 C1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y C0 N_20 VDD mp5  l=0.42u w=0.52u m=1
M9 Y B1 N_9 VDD mp5  l=0.42u w=0.52u m=1
M10 Y A1 N_21 VDD mp5  l=0.42u w=0.52u m=1
M11 N_21 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_9 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai222d0

* Top of hierarchy  cell=oai22d0
.subckt oai22d0 A0 A1 B1 B0 GND VDD Y
M1 Y B0 N_7 GND mn5  l=0.5u w=0.5u m=1
M2 Y B1 N_7 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_11 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M7 Y A1 N_10 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai22d0

* Top of hierarchy  cell=oai311d0
.subckt oai311d0 VDD Y GND C0 B0 A0 A1 A2
M1 N_11 A2 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_20 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_20 GND mn5  l=0.5u w=0.5u m=1
M6 N_7 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M7 N_8 A1 N_7 VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 VDD C0 Y VDD mp5  l=0.42u w=0.52u m=1

* Top of hierarchy  cell=oai31d0
.subckt oai31d0 A2 A0 A1 B0 Y VDD GND
M1 Y B0 N_7 GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_11 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_11 A0 N_10 VDD mp5  l=0.42u w=0.52u m=1
M8 N_10 A2 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oai31d0

* Top of hierarchy  cell=oai321d0
.subckt oai321d0 B1 B0 A0 A1 A2 C0 VDD Y GND
M1 Y C0 N_10 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A2 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_11 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 A0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_11 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_10 B1 N_11 GND mn5  l=0.5u w=0.5u m=1
M7 N_17 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_18 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_19 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_19 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M12 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai321d0

* Top of hierarchy  cell=oai322d0
.subckt oai322d0 VDD Y GND B0 A0 A1 A2 B1 C0 C1
M1 N_11 B0 N_13 GND mn5  l=0.5u w=0.5u m=1
M2 Y C1 N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_11 C0 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_13 B1 N_11 GND mn5  l=0.5u w=0.5u m=1
M5 N_13 A2 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_13 A1 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_13 A0 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_8 C1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y C0 N_8 VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 B1 Y VDD mp5  l=0.42u w=0.52u m=1
M11 Y A2 N_9 VDD mp5  l=0.42u w=0.52u m=1
M12 N_10 A1 N_9 VDD mp5  l=0.42u w=0.52u m=1
M13 N_10 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_3 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oai322d0

* Top of hierarchy  cell=oai32d0
.subckt oai32d0 A0 B1 A1 A2 B0 Y VDD GND
M1 N_7 B0 Y GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A2 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 B1 Y GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_16 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M8 N_17 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y B1 N_15 VDD mp5  l=0.42u w=0.52u m=1
M10 N_17 A0 N_16 VDD mp5  l=0.42u w=0.52u m=1
.ends oai32d0

* Top of hierarchy  cell=oai33d0
.subckt oai33d0 VDD Y GND B2 B1 B0 A1 A0 A2
M1 Y B0 N_12 GND mn5  l=0.5u w=0.5u m=1
M2 N_12 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 Y B2 N_12 GND mn5  l=0.5u w=0.5u m=1
M6 Y B1 N_12 GND mn5  l=0.5u w=0.5u m=1
M7 N_9 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_8 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_8 A0 N_7 VDD mp5  l=0.42u w=0.52u m=1
M10 N_7 A2 Y VDD mp5  l=0.42u w=0.52u m=1
M11 Y B2 N_6 VDD mp5  l=0.42u w=0.52u m=1
M12 N_9 B1 N_6 VDD mp5  l=0.42u w=0.52u m=1
.ends oai33d0

* Top of hierarchy  cell=oaim211d0
.subckt oaim211d0 B0 C0 A0N A1N GND VDD Y
M1 N_11 A1N N_4 GND mn5  l=0.5u w=0.5u m=1
M2 N_11 A0N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_12 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 Y C0 N_10 GND mn5  l=0.5u w=0.5u m=1
M5 N_12 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim211d0

* Top of hierarchy  cell=oaim21d0
.subckt oaim21d0 B0 A1N A0N VDD GND Y
M1 N_10 A0N N_3 GND mn5  l=0.5u w=0.5u m=1
M2 N_10 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 N_9 GND mn5  l=0.5u w=0.5u m=1
M4 N_9 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim21d0

* Top of hierarchy  cell=oaim22d0
.subckt oaim22d0 B1 B0 A0N A1N Y VDD GND
M1 N_11 A1N GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 A0N N_11 GND mn5  l=0.5u w=0.5u m=1
M3 N_7 N_4 Y GND mn5  l=0.5u w=0.5u m=1
M4 N_7 B0 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_7 B1 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_18 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_18 B1 Y VDD mp5  l=0.42u w=0.52u m=1
.ends oaim22d0

* Top of hierarchy  cell=oaim2m11d0
.subckt oaim2m11d0 C0 A0N B0N A1N VDD GND Y
M1 N_11 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_12 A1N GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 A0N N_12 GND mn5  l=0.5u w=0.5u m=1
M5 Y C0 N_11 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_7 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B0N N_7 VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim2m11d0

* Top of hierarchy  cell=oaim31d0
.subckt oaim31d0 GND Y VDD A1N A2N B0 A0N
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M2 N_6 B0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A2N GND GND mn5  l=0.5u w=0.5u m=1
M4 N_8 A1N N_7 GND mn5  l=0.5u w=0.5u m=1
M5 N_7 A0N N_4 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_4 A2N VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_4 A1N VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 A0N VDD VDD mp5  l=0.42u w=0.52u m=1
.ends oaim31d0

* Top of hierarchy  cell=or02d0
.subckt or02d0 A B VDD GND Y
M1 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M4 N_12 B N_3 VDD mp5  l=0.42u w=0.52u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or02d0

* Top of hierarchy  cell=or03d0
.subckt or03d0 B A C GND VDD Y
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_13 C N_3 VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A VDD VDD mp5  l=0.42u w=0.52u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_14 B N_13 VDD mp5  l=0.42u w=0.52u m=1
.ends or03d0

* Top of hierarchy  cell=or04d0
.subckt or04d0 A B D C VDD Y GND
M1 N_3 C GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 D GND GND mn5  l=0.5u w=0.5u m=1
M3 N_3 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_3 A GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 C N_14 VDD mp5  l=0.42u w=0.52u m=1
M7 N_14 D N_3 VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_16 A VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or04d0

* Top of hierarchy  cell=or12d0
.subckt or12d0 B AN VDD GND Y
M1 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M2 N_2 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_2 B GND GND mn5  l=0.5u w=0.5u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_14 B N_2 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or12d0

* Top of hierarchy  cell=or13d0
.subckt or13d0 C B AN Y VDD GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 AN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 B GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 C GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_15 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_16 B N_15 VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C N_16 VDD mp5  l=0.42u w=0.52u m=1
.ends or13d0


* Top of hierarchy  cell=or23d0
.subckt or23d0 AN C BN Y VDD GND
M1 N_6 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M2 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 BN GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 C GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_3 AN GND GND mn5  l=0.5u w=0.5u m=1
M7 N_18 N_7 N_17 VDD mp5  l=0.42u w=0.52u m=1
M8 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_7 BN VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C N_18 VDD mp5  l=0.42u w=0.52u m=1
M11 N_17 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_3 AN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends or23d0

* Top of hierarchy  cell=ora211d0
.subckt ora211d0 C0 B0 A1 A0 GND Y VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_8 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_11 B0 N_8 GND mn5  l=0.5u w=0.5u m=1
M5 N_6 C0 N_11 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_17 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 A1 N_17 VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 C0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora211d0

* Top of hierarchy  cell=ora21d0
.subckt ora21d0 B0 A1 A0 Y VDD GND
M1 Y N_5 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_6 A0 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 A1 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_5 B0 N_6 GND mn5  l=0.5u w=0.5u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M6 N_14 A0 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_5 A1 N_14 VDD mp5  l=0.42u w=0.52u m=1
M8 N_5 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora21d0

* Top of hierarchy  cell=ora31d0
.subckt ora31d0 B0 A2 A0 A1 Y VDD GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_7 A0 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_7 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_6 B0 N_7 GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M7 N_15 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_16 A0 N_15 VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A2 N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_6 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends ora31d0
* SPICE INPUT		Wed Jul 10 14:00:13 2019	ora31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d1
.subckt ora31d1 A0 A2 B0 A1 GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.58u m=1
M2 N_10 A1 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 B0 N_10 GND mn5  l=0.5u w=0.5u m=1
M4 N_10 A2 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_10 A0 GND GND mn5  l=0.5u w=0.5u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M7 N_15 A1 VDD VDD mp5  l=0.42u w=0.52u m=1
M8 N_6 B0 VDD VDD mp5  l=0.42u w=0.52u m=1
M9 N_6 A2 N_16 VDD mp5  l=0.42u w=0.52u m=1
M10 N_16 A0 N_15 VDD mp5  l=0.42u w=0.52u m=1
.ends ora31d1

* Top of hierarchy  cell=sdbfb1
.subckt sdbfb1 VDD Q QN GND RN SN SI SE D CKN
M1 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M2 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M3 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_4 CKN GND GND mn5  l=0.5u w=0.5u m=1
M6 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M7 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M9 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M10 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M11 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M12 N_9 N_5 N_29 GND mn5  l=0.5u w=0.5u m=1
M13 N_9 N_4 N_55 GND mn5  l=0.5u w=0.5u m=1
M14 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M16 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M17 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M18 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M19 N_11 N_4 N_56 GND mn5  l=0.5u w=0.5u m=1
M20 N_57 N_5 N_11 GND mn5  l=0.5u w=0.5u m=1
M21 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M23 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M24 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M25 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M26 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M27 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M28 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_4 CKN VDD VDD mp5  l=0.42u w=0.52u m=1
M30 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M31 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M33 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M34 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M35 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_9 N_4 N_7 VDD mp5  l=0.42u w=0.52u m=1
M37 N_19 N_5 N_9 VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M41 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M42 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_21 N_5 N_11 VDD mp5  l=0.42u w=0.52u m=1
M44 N_22 N_4 N_11 VDD mp5  l=0.42u w=0.5u m=1
M45 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M46 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M47 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M48 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdbfb1


* Top of hierarchy  cell=sdbrb1
.subckt sdbrb1 VDD Q QN GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_53 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_53 N_6 N_29 GND mn5  l=0.5u w=0.5u m=1
M6 N_54 SI N_29 GND mn5  l=0.5u w=0.5u m=1
M7 N_54 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_29 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_55 GND mn5  l=0.5u w=0.5u m=1
M10 N_55 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_27 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_27 N_13 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_27 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_56 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_56 GND mn5  l=0.5u w=0.5u m=1
M16 N_57 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M17 N_12 N_13 N_25 GND mn5  l=0.5u w=0.5u m=1
M18 N_25 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M19 N_13 RN GND GND mn5  l=0.5u w=0.5u m=1
M20 N_14 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M21 QN N_12 GND GND mn5  l=0.5u w=0.58u m=1
M22 Q N_14 GND GND mn5  l=0.5u w=0.58u m=1
M23 N_57 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M24 N_25 SN GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_17 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_17 VDD mp5  l=0.42u w=0.52u m=1
M30 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_18 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_19 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_19 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_20 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_20 N_13 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_21 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_21 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_22 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.52u m=1
M42 N_23 N_11 VDD VDD mp5  l=0.42u w=0.52u m=1
M43 N_13 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M44 QN N_12 VDD VDD mp5  l=0.42u w=0.76u m=1
M45 N_14 N_12 VDD VDD mp5  l=0.42u w=0.52u m=1
M46 Q N_14 VDD VDD mp5  l=0.42u w=0.76u m=1
M47 N_22 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M48 N_12 SN VDD VDD mp5  l=0.42u w=0.52u m=1
.ends sdbrb1

* Top of hierarchy  cell=sdbrq1
.subckt sdbrq1 VDD Q GND RN SN SI SE D CK
M1 N_4 CK GND GND mn5  l=0.5u w=0.5u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M3 N_6 SE GND GND mn5  l=0.5u w=0.5u m=1
M4 N_35 D GND GND mn5  l=0.5u w=0.5u m=1
M5 N_35 N_6 N_30 GND mn5  l=0.5u w=0.5u m=1
M6 N_36 SI N_30 GND mn5  l=0.5u w=0.5u m=1
M7 N_36 SE GND GND mn5  l=0.5u w=0.5u m=1
M8 N_9 N_4 N_30 GND mn5  l=0.5u w=0.5u m=1
M9 N_9 N_5 N_37 GND mn5  l=0.5u w=0.5u m=1
M10 N_37 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M11 N_28 N_9 N_10 GND mn5  l=0.5u w=0.5u m=1
M12 N_28 N_3 N_10 GND mn5  l=0.5u w=0.5u m=1
M13 N_28 SN GND GND mn5  l=0.5u w=0.5u m=1
M14 N_38 N_10 GND GND mn5  l=0.5u w=0.5u m=1
M15 N_11 N_5 N_38 GND mn5  l=0.5u w=0.5u m=1
M16 Q N_11 N_24 GND mn5  l=0.5u w=0.58u m=1
M17 N_24 N_3 Q GND mn5  l=0.5u w=0.58u m=1
M18 N_24 SN GND GND mn5  l=0.5u w=0.58u m=1
M19 N_3 RN GND GND mn5  l=0.5u w=0.5u m=1
M20 N_39 N_4 N_11 GND mn5  l=0.5u w=0.5u m=1
M21 N_39 N_12 GND GND mn5  l=0.5u w=0.5u m=1
M22 N_12 N_3 N_26 GND mn5  l=0.5u w=0.5u m=1
M23 N_26 N_11 N_12 GND mn5  l=0.5u w=0.5u m=1
M24 N_26 SN GND GND mn5  l=0.5u w=0.5u m=1
M25 N_4 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M26 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M27 N_6 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M28 N_15 D VDD VDD mp5  l=0.42u w=0.52u m=1
M29 N_7 SE N_15 VDD mp5  l=0.42u w=0.52u m=1
M30 N_16 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M31 N_16 SI VDD VDD mp5  l=0.42u w=0.52u m=1
M32 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.52u m=1
M33 N_17 N_4 N_9 VDD mp5  l=0.42u w=0.5u m=1
M34 N_17 N_10 VDD VDD mp5  l=0.42u w=0.5u m=1
M35 N_18 N_9 VDD VDD mp5  l=0.42u w=0.52u m=1
M36 N_18 N_3 N_10 VDD mp5  l=0.42u w=0.52u m=1
M37 N_10 SN VDD VDD mp5  l=0.42u w=0.52u m=1
M38 N_19 N_10 VDD VDD mp5  l=0.42u w=0.52u m=1
M39 N_19 N_4 N_11 VDD mp5  l=0.42u w=0.52u m=1
M40 N_20 N_5 N_11 VDD mp5  l=0.42u w=0.5u m=1
M41 N_22 N_11 VDD VDD mp5  l=0.42u w=0.76u m=1
M42 Q N_3 N_22 VDD mp5  l=0.42u w=0.76u m=1
M43 Q SN VDD VDD mp5  l=0.42u w=0.76u m=1
M44 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M45 N_20 N_12 VDD VDD mp5  l=0.42u w=0.5u m=1
M46 N_21 N_3 N_12 VDD mp5  l=0.42u w=0.5u m=1
M47 N_21 N_11 VDD VDD mp5  l=0.42u w=0.5u m=1
M48 N_12 SN VDD VDD mp5  l=0.42u w=0.5u m=1
.ends sdbrq1


* Top of hierarchy  cell=tlatncad1
.subckt tlatncad1 VDD ECK GND CK E
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_21 E GND GND mn5  l=0.5u w=0.5u m=1
M3 N_21 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M4 N_22 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M5 N_22 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 ECK N_5 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_6 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M8 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_3 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_9 E VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_10 N_3 N_5 VDD mp5  l=0.42u w=0.5u m=1
M13 N_9 N_4 N_5 VDD mp5  l=0.42u w=0.52u m=1
M14 N_10 N_6 VDD VDD mp5  l=0.42u w=0.5u m=1
M15 N_11 N_5 ECK VDD mp5  l=0.42u w=0.76u m=1
M16 N_6 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_11 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
.ends tlatncad1

* Top of hierarchy  cell=tlatntscad1
.subckt tlatntscad1 VDD ECK GND CK SE E
M1 N_4 E GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 SE GND GND mn5  l=0.5u w=0.5u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M5 N_27 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_27 N_3 N_7 GND mn5  l=0.5u w=0.5u m=1
M7 N_28 N_6 N_7 GND mn5  l=0.5u w=0.5u m=1
M8 N_28 N_8 GND GND mn5  l=0.5u w=0.5u m=1
M9 ECK N_7 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_8 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M11 ECK N_3 GND GND mn5  l=0.5u w=0.58u m=1
M12 N_3 CK GND GND mn5  l=0.5u w=0.5u m=1
M13 N_11 E N_4 VDD mp5  l=0.42u w=0.52u m=1
M14 N_11 SE VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M16 N_6 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_12 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M18 N_13 N_3 N_7 VDD mp5  l=0.42u w=0.5u m=1
M19 N_12 N_6 N_7 VDD mp5  l=0.42u w=0.52u m=1
M20 N_13 N_8 VDD VDD mp5  l=0.42u w=0.5u m=1
M21 N_14 N_7 ECK VDD mp5  l=0.42u w=0.76u m=1
M22 N_8 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M23 N_14 N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M24 N_3 CK VDD VDD mp5  l=0.42u w=0.52u m=1
.ends tlatntscad1





* Top of hierarchy  cell=lachb1
.subckt lachb1 RN D G GND QN Q VDD
M1 N_5 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_7 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.5u m=1
M5 N_19 N_5 N_3 GND mn5  l=0.5u w=0.5u m=1
M6 N_21 RN N_20 GND mn5  l=0.5u w=0.5u m=1
M7 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M8 N_2 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M9 Q N_3 GND GND mn5  l=0.5u w=0.58u m=1
M10 N_20 N_7 N_3 GND mn5  l=0.5u w=0.5u m=1
M11 N_21 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M12 N_5 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_7 G VDD VDD mp5  l=0.42u w=0.52u m=1
M14 N_31 D VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_3 N_7 N_31 VDD mp5  l=0.42u w=0.52u m=1
M16 N_3 RN VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_32 N_5 N_3 VDD mp5  l=0.42u w=0.52u m=1
M18 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M19 Q N_3 VDD VDD mp5  l=0.42u w=0.76u m=1
M20 N_2 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M21 N_32 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lachb1



* Top of hierarchy  cell=lanhb1
.subckt lanhb1 D G GND QN Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_15 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_5 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_16 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M9 N_16 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_25 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_5 N_4 N_25 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 Q N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_26 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M18 N_26 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhb1

* Top of hierarchy  cell=lanhn1
.subckt lanhn1 D G GND QN VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhn1

* Top of hierarchy  cell=lanhq1
.subckt lanhq1 D G GND Q VDD
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_3 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_4 G VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanhq1



* Top of hierarchy  cell=lanlb1
.subckt lanlb1 GND QN Q VDD D GN
M1 N_5 N_4 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_4 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_10 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_7 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_7 N_6 GND GND mn5  l=0.5u w=0.5u m=1
M6 Q N_6 GND GND mn5  l=0.5u w=0.58u m=1
M7 N_11 N_5 N_6 GND mn5  l=0.5u w=0.5u m=1
M8 N_10 N_4 N_6 GND mn5  l=0.5u w=0.5u m=1
M9 N_11 N_7 GND GND mn5  l=0.5u w=0.5u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_4 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M13 N_6 N_5 N_22 VDD mp5  l=0.42u w=0.52u m=1
M14 QN N_7 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 Q N_6 VDD VDD mp5  l=0.42u w=0.76u m=1
M16 N_7 N_6 VDD VDD mp5  l=0.42u w=0.52u m=1
M17 N_23 N_4 N_6 VDD mp5  l=0.42u w=0.52u m=1
M18 N_23 N_7 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlb1


* Top of hierarchy  cell=lanln1
.subckt lanln1 D GN GND QN VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_14 D GND GND mn5  l=0.5u w=0.5u m=1
M4 QN N_2 GND GND mn5  l=0.5u w=0.58u m=1
M5 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M6 N_15 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_14 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_15 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_23 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_23 VDD mp5  l=0.42u w=0.52u m=1
M13 QN N_2 VDD VDD mp5  l=0.42u w=0.76u m=1
M14 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M15 N_24 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_24 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanln1

* Top of hierarchy  cell=lanlq1
.subckt lanlq1 D GN GND Q VDD
M1 N_4 N_3 GND GND mn5  l=0.5u w=0.5u m=1
M2 N_3 GN GND GND mn5  l=0.5u w=0.5u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.5u m=1
M4 N_2 N_5 GND GND mn5  l=0.5u w=0.5u m=1
M5 Q N_5 GND GND mn5  l=0.5u w=0.58u m=1
M6 N_14 N_4 N_5 GND mn5  l=0.5u w=0.5u m=1
M7 N_13 N_3 N_5 GND mn5  l=0.5u w=0.5u m=1
M8 N_14 N_2 GND GND mn5  l=0.5u w=0.5u m=1
M9 N_4 N_3 VDD VDD mp5  l=0.42u w=0.52u m=1
M10 N_3 GN VDD VDD mp5  l=0.42u w=0.52u m=1
M11 N_22 D VDD VDD mp5  l=0.42u w=0.52u m=1
M12 N_5 N_4 N_22 VDD mp5  l=0.42u w=0.52u m=1
M13 N_2 N_5 VDD VDD mp5  l=0.42u w=0.52u m=1
M14 Q N_5 VDD VDD mp5  l=0.42u w=0.76u m=1
M15 N_23 N_3 N_5 VDD mp5  l=0.42u w=0.52u m=1
M16 N_23 N_2 VDD VDD mp5  l=0.42u w=0.52u m=1
.ends lanlq1
