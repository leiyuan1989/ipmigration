

.SUBCKT DFFHQNX1MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFHQNX2MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQNX4MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=6.1e-07
.ends


.SUBCKT DFFHQNX8MTR QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm nmin net063 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net063 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.4e-07
mXI43_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_3 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g9_MXNA1_4 QN s VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net051 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net051 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5e-07
MXP2 net050 c VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm nmin net050 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI43_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_3 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g9_MXPA1_4 QN s VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQX1MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=3.4e-07
MXN3 net87 cn VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP4 net061 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm nmin net62 VNW p12 l=1.3e-07 w=4.1e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.4e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.4e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFHQX2MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=4.8e-07
MXN4 net87 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP6 net061 c cn VNW p12 l=1.3e-07 w=4.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP7 pm nmin net62 VNW p12 l=1.3e-07 w=5.9e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.4e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQX4MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net87 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=7.4e-07
MXP8 net061 c cn VNW p12 l=1.3e-07 w=7.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP9 pm nmin net62 VNW p12 l=1.3e-07 w=8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI36_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHQX8MTR Q VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=4.4e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net87 VPW n12 l=1.3e-07 w=6.9e-07
MXN5 net87 cn VSS VPW n12 l=1.3e-07 w=6.9e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNOE pm c XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.2e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=7.2e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=6.9e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP0 net061 CK VDD VNW p12 l=1.3e-07 w=7.3e-07
MXP10 net061 c cn VNW p12 l=1.3e-07 w=7.3e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.5e-07
mX_g10_MXPA1_2 c nck VDD VNW p12 l=1.3e-07 w=8.5e-07
MXP2 net62 c VDD VNW p12 l=1.3e-07 w=8e-07
MXP9 pm nmin net62 VNW p12 l=1.3e-07 w=8e-07
mXI12_MXPOEN pm cn XI12_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI36_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=7.3e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.4e-07
.ends


.SUBCKT DFFHX1MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=3.6e-07
MXN3 net42 cn VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP5 net63 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.3e-07
MXP2 net53 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP6 pm nmin net53 VNW p12 l=1.3e-07 w=4.4e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.9e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFHX2MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=5.1e-07
MXN4 net42 cn VSS VPW n12 l=1.3e-07 w=5.1e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP7 net63 c cn VNW p12 l=1.3e-07 w=4.6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8e-07
MXP8 net53 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP10 pm nmin net53 VNW p12 l=1.3e-07 w=6.2e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=5.8e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI32_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.1e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT DFFHX4MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=7e-07
MXN5 net42 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP11 net63 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP8 net53 c VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP12 pm nmin net53 VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI32_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT DFFHX8MTR Q QN VDD VNW VPW VSS CK D
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.2e-07
MXN1 pm nmin net42 VPW n12 l=1.3e-07 w=7e-07
MXN5 net42 cn VSS VPW n12 l=1.3e-07 w=7e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI32_MXNOE bm c m VPW n12 l=1.3e-07 w=7.3e-07
mXI1_MXNOE bm cn XI1_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA1 XI1_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net63 CK VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP11 net63 c cn VNW p12 l=1.3e-07 w=6.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP8 net53 c VDD VNW p12 l=1.3e-07 w=8.6e-07
MXP12 pm nmin net53 VNW p12 l=1.3e-07 w=8.6e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI32_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.4e-07
mXI32_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=8.2e-07
mXI1_MXPOEN bm c XI1_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA1 XI1_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=2.3e-07
.ends


.SUBCKT DFFNHX1MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=4.3e-07
MXN2 net67 cn VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net56 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=6.8e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP3 pm net150 net42 VNW p12 l=1.3e-07 w=3.3e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=4.8e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.8e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNHX2MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=6.1e-07
MXN3 net67 cn VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=5.7e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP1 net56 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1_2 cn nckn VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP4 pm net150 net42 VNW p12 l=1.3e-07 w=4.6e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNHX4MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=5.4e-07
MXN3 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN3_2 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 pm net150 net67 VPW n12 l=1.3e-07 w=5.4e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=5.4e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI37_MXNOE_2 bm c m VPW n12 l=1.3e-07 w=5.1e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP5 net56 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=6.6e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g10_MXPA1_2 cn nckn VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 pm net150 net42 VNW p12 l=1.3e-07 w=6.9e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI37_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.3e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mXI52_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNHX8MTR Q QN VDD VNW VPW VSS CKN D
mX_g14_MXNA1 nckn CKN VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN0 c CKN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g13_MXNA1 net150 D VSS VPW n12 l=1.3e-07 w=5e-07
mX_g13_MXNA1_2 net150 D VSS VPW n12 l=1.3e-07 w=5e-07
mX_g10_MXNA1 cn nckn VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN1 pm net150 net67 VPW n12 l=1.3e-07 w=7.4e-07
MXN3 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN3_2 net67 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MXN1_2 pm net150 net67 VPW n12 l=1.3e-07 w=5.7e-07
mXI10_MXNOE pm c XI10_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI10_MXNA1 XI10_n1 m VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=7.4e-07
mXI37_MXNOE bm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI37_MXNOE_2 bm c m VPW n12 l=1.3e-07 w=6.1e-07
mXI11_MXNOE bm cn XI11_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI52_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI52_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI54_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXPA1 nckn CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP0 net56 CKN VDD VNW p12 l=1.3e-07 w=6.4e-07
MXP7 net56 cn c VNW p12 l=1.3e-07 w=6.4e-07
mX_g13_MXPA1 net150 D VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g13_MXPA1_2 net150 D VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g10_MXPA1 cn nckn VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g10_MXPA1_2 cn nckn VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP2 net42 c VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 pm net150 net42 VNW p12 l=1.3e-07 w=6.9e-07
mXI10_MXPOEN pm cn XI10_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI10_MXPA1 XI10_p1 m VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI37_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI37_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
mXI11_MXPOEN bm c XI11_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=4.1e-07
mXI52_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI52_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI52_MXPA1_5 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI54_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.6e-07
.ends


.SUBCKT DFFNSRHX1MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS SN net68 VPW n12 l=1.3e-07 w=4.3e-07
MXN11 net68 cn net72 VPW n12 l=1.3e-07 w=4.3e-07
MXN0 pm nmin net72 VPW n12 l=1.3e-07 w=4.3e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 m pm net80 VPW n12 l=1.3e-07 w=4.5e-07
MXN13 VSS RN net80 VPW n12 l=1.3e-07 w=4.5e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
MXN7 bm cn net91 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net91 RN net88 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net88 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net152 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP13 net152 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmin net118 VNW p12 l=1.3e-07 w=3.3e-07
MXP9 net118 c VDD VNW p12 l=1.3e-07 w=3.3e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=4.8e-07
MXP1 net142 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net142 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.8e-07
MXP16 bm nmset net154 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net154 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP18 bm c net110 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net110 nmset net114 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net114 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT DFFNSRHX2MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=3e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS SN net70 VPW n12 l=1.3e-07 w=6e-07
MXN16 net70 cn net66 VPW n12 l=1.3e-07 w=6e-07
MXN0 pm nmin net66 VPW n12 l=1.3e-07 w=6e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 m pm net78 VPW n12 l=1.3e-07 w=6.3e-07
MXN18 VSS RN net78 VPW n12 l=1.3e-07 w=6.3e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.6e-07
MXN7 bm cn net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net89 RN net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net154 CKN VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP13 net154 cn c VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 pm nmin net120 VNW p12 l=1.3e-07 w=4.6e-07
MXP9 net120 c VDD VNW p12 l=1.3e-07 w=4.6e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP1 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP20 bm nmset net104 VNW p12 l=1.3e-07 w=2.8e-07
MXP4 net104 RN VDD VNW p12 l=1.3e-07 w=2.8e-07
MXP18 bm c net112 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net112 nmset net116 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net116 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFNSRHX4MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=3e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=4.6e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN20 VSS SN net67 VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net67 cn net71 VPW n12 l=1.3e-07 w=7.5e-07
MXN0 pm nmin net71 VPW n12 l=1.3e-07 w=7.5e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN4 m pm net79 VPW n12 l=1.3e-07 w=8.4e-07
MXN21 VSS RN net79 VPW n12 l=1.3e-07 w=8.4e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN7 bm cn net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net90 RN net87 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net87 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net155 CKN VDD VNW p12 l=1.3e-07 w=5e-07
MXP21 net155 cn c VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.6e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP22 pm nmin net121 VNW p12 l=1.3e-07 w=6.9e-07
MXP9 net121 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP11_2 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP1 net145 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net145 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP23 bm nmset net105 VNW p12 l=1.3e-07 w=3.6e-07
MXP4 net105 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP18 bm c net113 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net113 nmset net117 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net117 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFNSRHX8MTR Q QN VDD VNW VPW VSS CKN D RN SN
mX_g14_MXNA1 nck CKN VSS VPW n12 l=1.3e-07 w=5.4e-07
MXN2 c CKN VSS VPW n12 l=1.3e-07 w=3.8e-07
mX_g10_MXNA1 cn nck VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g10_MXNA1_2 cn nck VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.4e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN20 VSS SN net66 VPW n12 l=1.3e-07 w=7.5e-07
MXN19 net66 cn net70 VPW n12 l=1.3e-07 w=7.5e-07
MXN0 pm nmin net70 VPW n12 l=1.3e-07 w=7.5e-07
mXI19_MXNOE pm c XI19_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI19_MXNA1 XI19_n1 m VSS VPW n12 l=1.3e-07 w=2.5e-07
MXN4 m pm net78 VPW n12 l=1.3e-07 w=8.7e-07
MXN22 VSS RN net78 VPW n12 l=1.3e-07 w=8.7e-07
MXN6 m nmset VSS VPW n12 l=1.3e-07 w=2e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN7 bm cn net89 VPW n12 l=1.3e-07 w=1.8e-07
MXN14 net89 RN net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN15 VSS s net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 bm nmset VSS VPW n12 l=1.3e-07 w=3e-07
mX_g11_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CKN VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP2 net154 CKN VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP24 net154 cn c VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 cn nck VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g10_MXPA1_2 cn nck VDD VNW p12 l=1.3e-07 w=8.4e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=1.03e-06
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=3.3e-07
MXP12 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP22 pm nmin net120 VNW p12 l=1.3e-07 w=6.9e-07
MXP9 net120 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI19_MXPOEN pm cn XI19_p1 VNW p12 l=1.3e-07 w=3.1e-07
mXI19_MXPA1 XI19_p1 m VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP11 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP11_2 m pm VDD VNW p12 l=1.3e-07 w=5.2e-07
MXP1 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP15 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP25 bm nmset net104 VNW p12 l=1.3e-07 w=3.5e-07
MXP4 net104 RN VDD VNW p12 l=1.3e-07 w=3.5e-07
MXP18 bm c net112 VNW p12 l=1.3e-07 w=2.3e-07
MXP17 net112 nmset net116 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net116 VNW p12 l=1.3e-07 w=2.3e-07
mX_g11_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=3.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQNX1MTR QN VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE nm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE nm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN nm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN nm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFQNX2MTR QN VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE nm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE nm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN nm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN nm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQNX4MTR QN VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNOE nm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI7_MXNOE nm cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g1_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN nm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI7_MXPOEN nm c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g1_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQX1MTR Q VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI6_MXNOE ns c XI6_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI7_MXNOE ns cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI6_MXPOEN ns cn XI6_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI7_MXPOEN ns c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFQX2MTR Q VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI6_MXNOE ns c XI6_n1 VPW n12 l=1.3e-07 w=3.6e-07
mXI7_MXNOE ns cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI6_MXPOEN ns cn XI6_p1 VNW p12 l=1.3e-07 w=4.9e-07
mXI7_MXPOEN ns c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g1_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFQX4MTR Q VDD VNW VPW VSS CK D
mXI4_MXNA1 XI4_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=4.2e-07
mXI6_MXNOE ns c XI6_n1 VPW n12 l=1.3e-07 w=4.2e-07
mXI7_MXNOE ns cn XI7_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI7_MXNA1 XI7_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s ns VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q ns VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI4_MXPA1 XI4_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm c XI4_p1 VNW p12 l=1.3e-07 w=3e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI6_MXPOEN ns cn XI6_p1 VNW p12 l=1.3e-07 w=6.1e-07
mXI7_MXPOEN ns c XI7_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI7_MXPA1 XI7_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s ns VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g1_MXPA1 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q ns VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRHQX1MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.2e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net89 cn VSS VPW n12 l=1.3e-07 w=3.5e-07
MXN2 pm nmin net89 VPW n12 l=1.3e-07 w=3.5e-07
MXN3 pm c net66 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net66 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net73 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
MXN11 m pm net73 VPW n12 l=1.3e-07 w=4.9e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=3.7e-07
MXN7 bm cn net85 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net85 RN net82 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net82 VPW n12 l=1.3e-07 w=1.5e-07
mXI52_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net126 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP11 net126 c cn VNW p12 l=1.3e-07 w=4.2e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6.1e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP2 net134 c VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP12 pm nmin net134 VNW p12 l=1.3e-07 w=4.2e-07
MXP14 pm cn net104 VNW p12 l=1.3e-07 w=2.3e-07
MXP5 VDD m net104 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.3e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=2.3e-07
MXP16 bm c net120 VNW p12 l=1.3e-07 w=2.3e-07
MXP15 VDD s net120 VNW p12 l=1.3e-07 w=2.3e-07
mXI52_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFRHQX2MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN15 net90 cn VSS VPW n12 l=1.3e-07 w=5.1e-07
MXN2 pm nmin net90 VPW n12 l=1.3e-07 w=5.1e-07
MXN3 pm c net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 net74 RN VSS VPW n12 l=1.3e-07 w=6.8e-07
MXN11 m pm net74 VPW n12 l=1.3e-07 w=6.8e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=5.4e-07
MXN7 bm cn net86 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net86 RN net83 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net83 VPW n12 l=1.3e-07 w=1.5e-07
mXI50_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI51_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=3.4e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net131 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP18 net131 c cn VNW p12 l=1.3e-07 w=4.5e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP19 pm nmin net105 VNW p12 l=1.3e-07 w=6.2e-07
MXP20 pm cn net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP5 VDD m net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=8.5e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.1e-07
mXI58_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=5.3e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=2.7e-07
MXP21 bm c net125 VNW p12 l=1.3e-07 w=1.5e-07
MXP15 VDD s net125 VNW p12 l=1.3e-07 w=1.5e-07
mXI50_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRHQX4MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MXN15 net90 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm nmin net90 VPW n12 l=1.3e-07 w=5.1e-07
MXN3 pm c net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net74 RN VSS VPW n12 l=1.3e-07 w=5.9e-07
MXN11 m pm net74 VPW n12 l=1.3e-07 w=5.9e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MXN7 bm cn net86 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net86 RN net83 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net83 VPW n12 l=1.3e-07 w=1.5e-07
mXI50_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net131 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP18 net131 c cn VNW p12 l=1.3e-07 w=4.5e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
MXP2 net105 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP19 pm nmin net105 VNW p12 l=1.3e-07 w=6.2e-07
MXP20 pm cn net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP5 VDD m net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP6_2 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI58_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=3e-07
MXP21 bm c net125 VNW p12 l=1.3e-07 w=1.5e-07
MXP15 VDD s net125 VNW p12 l=1.3e-07 w=1.5e-07
mXI50_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRHQX8MTR Q VDD VNW VPW VSS CK D RN
mXI47_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mXI48_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI49_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MXN15 net90 cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 pm nmin net90 VPW n12 l=1.3e-07 w=5.1e-07
MXN3 pm c net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS m net67 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 net74 RN VSS VPW n12 l=1.3e-07 w=5.9e-07
MXN11 m pm net74 VPW n12 l=1.3e-07 w=5.9e-07
mXI58_MXNOE bm c m VPW n12 l=1.3e-07 w=4.6e-07
MXN7 bm cn net86 VPW n12 l=1.3e-07 w=1.5e-07
MXN13 net86 RN net83 VPW n12 l=1.3e-07 w=1.5e-07
MXN14 VSS s net83 VPW n12 l=1.3e-07 w=1.5e-07
mXI50_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI51_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI51_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI47_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP0 net131 CK VDD VNW p12 l=1.3e-07 w=4.5e-07
MXP18 net131 c cn VNW p12 l=1.3e-07 w=4.5e-07
mXI48_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.8e-07
mXI49_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7.1e-07
MXP2 net105 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP19 pm nmin net105 VNW p12 l=1.3e-07 w=6.2e-07
MXP20 pm cn net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP5 VDD m net109 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 m pm VDD VNW p12 l=1.3e-07 w=5.5e-07
MXP6_2 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
MXP7 m RN VDD VNW p12 l=1.3e-07 w=2.7e-07
mXI58_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4e-07
mXI58_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP17 VDD RN bm VNW p12 l=1.3e-07 w=3e-07
MXP21 bm c net125 VNW p12 l=1.3e-07 w=1.5e-07
MXP15 VDD s net125 VNW p12 l=1.3e-07 w=1.5e-07
mXI50_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI51_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI51_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRQX1MTR Q VDD VNW VPW VSS CK D RN
MXN5 net86 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net78 D net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 pm cn net78 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 pm c net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net66 m net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net66 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI37_MXNOE net119 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE net119 cn XI4_n1 VPW n12 l=1.3e-07 w=2.3e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=2.3e-07
mXI0_MXNA1 s net119 XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA2 XI0_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP4 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 D VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP6 pm c net105 VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI37_MXPOEN net119 cn m VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN net119 c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 s net119 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFRQX2MTR Q VDD VNW VPW VSS CK D RN
MXN5 net86 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net78 D net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 pm cn net78 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 pm c net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net66 m net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net66 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI37_MXNOE net119 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE net119 cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 s net119 XI0_n1 VPW n12 l=1.3e-07 w=2.7e-07
mXI0_MXNA2 XI0_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 D VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP6 pm c net105 VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3e-07
mXI37_MXPOEN net119 cn m VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN net119 c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 s net119 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRQX4MTR Q VDD VNW VPW VSS CK D RN
MXN5 net86 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net78 D net86 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 pm cn net78 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 pm c net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN9 net66 m net71 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net66 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g4_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI37_MXNOE net119 c m VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE net119 cn XI4_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI0_MXNA1 s net119 XI0_n1 VPW n12 l=1.3e-07 w=4.9e-07
mXI0_MXNA2 XI0_n1 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net105 D VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP6 pm c net105 VNW p12 l=1.3e-07 w=4.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=3e-07
MXP8 pm cn net89 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD m net89 VNW p12 l=1.3e-07 w=2.3e-07
mX_g4_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3e-07
mXI37_MXPOEN net119 cn m VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN net119 c XI4_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI0_MXPA1 s net119 VDD VNW p12 l=1.3e-07 w=3e-07
mXI0_MXPA2 s RN VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRX1MTR Q QN VDD VNW VPW VSS CK D RN
MXN2 pm cn net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net45 D net53 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net53 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 pm c net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net61 m net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net61 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE bm cn XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 net90 VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 net90 bm XI1_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI45_MXNA1 Q net90 VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP2 net68 D VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm c net68 VNW p12 l=1.3e-07 w=4.1e-07
MXP1 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MXP7 pm cn net72 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD m net72 VNW p12 l=1.3e-07 w=2.3e-07
mXI43_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI40_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI5_MXPOEN bm c XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 net90 VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA2 net90 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 net90 bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mXI45_MXPA1 Q net90 VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFRX2MTR Q QN VDD VNW VPW VSS CK D RN
MXN2 pm cn net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net45 D net53 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net53 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 pm c net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net61 m net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net61 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE bm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 net90 VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=2.7e-07
mXI1_MXNA1 net90 bm XI1_n1 VPW n12 l=1.3e-07 w=2.7e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI45_MXNA1 Q net90 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP2 net68 D VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm c net68 VNW p12 l=1.3e-07 w=4.1e-07
MXP1 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 pm cn net72 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 VDD m net72 VNW p12 l=1.3e-07 w=2.2e-07
mXI43_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI40_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI5_MXPOEN bm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 net90 VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 net90 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI1_MXPA1 net90 bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI45_MXPA1 Q net90 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFRX4MTR Q QN VDD VNW VPW VSS CK D RN
MXN2 pm cn net45 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 net45 D net53 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 net53 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI41_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI42_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN9 pm c net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 net61 m net58 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 net61 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI43_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI40_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNOE bm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 net90 VSS VPW n12 l=1.3e-07 w=1.5e-07
mXI1_MXNA2 XI1_n1 RN VSS VPW n12 l=1.3e-07 w=4.9e-07
mXI1_MXNA1 net90 bm XI1_n1 VPW n12 l=1.3e-07 w=4.9e-07
mXI46_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI46_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI45_MXNA1 Q net90 VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI45_MXNA1_2 Q net90 VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP2 net68 D VDD VNW p12 l=1.3e-07 w=4.1e-07
MXP5 pm c net68 VNW p12 l=1.3e-07 w=4.1e-07
MXP1 pm RN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI41_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mXI42_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
MXP8 pm cn net72 VNW p12 l=1.3e-07 w=2.2e-07
MXP6 VDD m net72 VNW p12 l=1.3e-07 w=2.2e-07
mXI43_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mXI40_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.6e-07
mXI5_MXPOEN bm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 net90 VDD VNW p12 l=1.3e-07 w=1.5e-07
mXI1_MXPA2 net90 RN VDD VNW p12 l=1.3e-07 w=3e-07
mXI1_MXPA1 net90 bm VDD VNW p12 l=1.3e-07 w=3e-07
mXI46_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI46_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI45_MXPA1 Q net90 VDD VNW p12 l=1.3e-07 w=8.7e-07
mXI45_MXPA1_2 Q net90 VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSHQX1MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN8 VSS SN net92 VPW n12 l=1.3e-07 w=4.5e-07
MXN7 net92 cn net89 VPW n12 l=1.3e-07 w=4.5e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=4.5e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP7 net099 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 pm nmin net091 VNW p12 l=1.3e-07 w=3.7e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=3.7e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT DFFSHQX2MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.7e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN12 VSS SN net92 VPW n12 l=1.3e-07 w=6.4e-07
MXN11 net92 cn net89 VPW n12 l=1.3e-07 w=6.4e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=6.4e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.1e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP13 net099 c cn VNW p12 l=1.3e-07 w=4.9e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7.6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP14 pm nmin net091 VNW p12 l=1.3e-07 w=5.4e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.9e-07
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSHQX4MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN14 VSS SN net92 VPW n12 l=1.3e-07 w=7.5e-07
MXN13 net92 cn net89 VPW n12 l=1.3e-07 w=7.5e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=7.5e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP15 net099 c cn VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP16 pm nmin net091 VNW p12 l=1.3e-07 w=6.9e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSHQX8MTR Q VDD VNW VPW VSS CK D SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN1 cn CK VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=4.5e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g5_MXNA1 nmset_ SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN14 VSS SN net92 VPW n12 l=1.3e-07 w=7.5e-07
MXN13 net92 cn net89 VPW n12 l=1.3e-07 w=7.5e-07
MXN3 pm nmin net89 VPW n12 l=1.3e-07 w=7.5e-07
mXI6_MXNOE pm c XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=7.8e-07
mXI53_MXNOE bm c m VPW n12 l=1.3e-07 w=8.7e-07
MXN9 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN10 VSS s net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 bm nmset_ VSS VPW n12 l=1.3e-07 w=3e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=3e-07
MXP2 net099 CK VDD VNW p12 l=1.3e-07 w=8.1e-07
MXP15 net099 c cn VNW p12 l=1.3e-07 w=8.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=9.9e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g5_MXPA1 nmset_ SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=3.8e-07
MXP16 pm nmin net091 VNW p12 l=1.3e-07 w=6.9e-07
MXP1 net091 c VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI6_MXPA1 XI6_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPOEN pm cn XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mX_g7_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
mXI53_MXPOEN bm cn m VNW p12 l=1.3e-07 w=1.15e-06
MXP12 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP11 net73 nmset_ net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP10 VDD s net76 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSQX1MTR Q VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN2 bm cn net84 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 NSN s net84 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI34_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm c net62 VNW p12 l=1.3e-07 w=2.3e-07
MXP7 VDD s net62 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSQX2MTR Q VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN2 bm cn net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 NSN s net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN1 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI34_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 bm c net53 VNW p12 l=1.3e-07 w=1.5e-07
MXP7 VDD s net53 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSQX4MTR Q VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=2.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI34_MXNOE bm c m VPW n12 l=1.3e-07 w=1.8e-07
MXN2 bm cn net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN5 NSN s net39 VPW n12 l=1.3e-07 w=1.5e-07
MXN1 NSN SN VSS VPW n12 l=1.3e-07 w=3.7e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI34_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP6 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP9 bm c net53 VNW p12 l=1.3e-07 w=1.5e-07
MXP7 VDD s net53 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRHQX1MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN13 VSS SN net62 VPW n12 l=1.3e-07 w=4.1e-07
MXN12 net62 cn net82 VPW n12 l=1.3e-07 w=4.1e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=4.1e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=4.3e-07
MXN14 VSS RN net70 VPW n12 l=1.3e-07 w=4.3e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=3.8e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net122 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP16 pm nmin net128 VNW p12 l=1.3e-07 w=3.1e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=3.1e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=4.6e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP17 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.6e-07
MXP23 bm nmset net112 VNW p12 l=1.3e-07 w=2.3e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSRHQX2MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN21 VSS SN net62 VPW n12 l=1.3e-07 w=5.8e-07
MXN20 net62 cn net82 VPW n12 l=1.3e-07 w=5.8e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=5.8e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=6.1e-07
MXN22 VSS RN net70 VPW n12 l=1.3e-07 w=6.1e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=4.2e-07
MXP15 net122 c cn VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=7e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=2.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP25 pm nmin net128 VNW p12 l=1.3e-07 w=4.5e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=4.5e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP17 m RN net144 VNW p12 l=1.3e-07 w=2.3e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP27 bm nmset net112 VNW p12 l=1.3e-07 w=2.7e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=2.7e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRHQX4MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS SN net62 VPW n12 l=1.3e-07 w=7.5e-07
MXN23 net62 cn net82 VPW n12 l=1.3e-07 w=7.5e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=7.5e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN25 VSS RN net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP28 net122 c cn VNW p12 l=1.3e-07 w=6.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.03e-06
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP29 pm nmin net128 VNW p12 l=1.3e-07 w=6.8e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP30 m RN net144 VNW p12 l=1.3e-07 w=3.1e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP31 bm nmset net112 VNW p12 l=1.3e-07 w=3.6e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRHQX8MTR Q VDD VNW VPW VSS CK D RN SN
mX_g14_MXNA1 nck CK VSS VPW n12 l=1.3e-07 w=2.6e-07
MXN10 cn CK VSS VPW n12 l=1.3e-07 w=2.6e-07
mX_g10_MXNA1 c nck VSS VPW n12 l=1.3e-07 w=3.9e-07
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g5_MXNA1 nmset SN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN24 VSS SN net62 VPW n12 l=1.3e-07 w=7.5e-07
MXN23 net62 cn net82 VPW n12 l=1.3e-07 w=7.5e-07
MXN1 pm nmin net82 VPW n12 l=1.3e-07 w=7.5e-07
mXI9_MXNOE pm c XI9_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI9_MXNA1 XI9_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 m pm net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN25 VSS RN net70 VPW n12 l=1.3e-07 w=7.2e-07
MXN5 m nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mXI62_MXNOE bm c m VPW n12 l=1.3e-07 w=5.5e-07
MXN18 bm cn net101 VPW n12 l=1.3e-07 w=1.8e-07
MXN19 net101 RN net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN17 VSS s net90 VPW n12 l=1.3e-07 w=1.8e-07
MXN16 bm nmset VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 nck CK VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP2 net122 CK VDD VNW p12 l=1.3e-07 w=6.1e-07
MXP28 net122 c cn VNW p12 l=1.3e-07 w=6.1e-07
mX_g10_MXPA1 c nck VDD VNW p12 l=1.3e-07 w=1.03e-06
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g5_MXPA1 nmset SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP4 pm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP29 pm nmin net128 VNW p12 l=1.3e-07 w=6.8e-07
MXP1 net128 c VDD VNW p12 l=1.3e-07 w=6.8e-07
mXI9_MXPOEN pm cn XI9_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI9_MXPA1 XI9_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 m pm VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP18 net144 nmset VDD VNW p12 l=1.3e-07 w=3.1e-07
MXP30 m RN net144 VNW p12 l=1.3e-07 w=3.1e-07
mXI62_MXPOEN bm cn m VNW p12 l=1.3e-07 w=6.7e-07
MXP31 bm nmset net112 VNW p12 l=1.3e-07 w=3.6e-07
MXP22 net112 RN VDD VNW p12 l=1.3e-07 w=3.6e-07
MXP19 bm c net108 VNW p12 l=1.3e-07 w=2.3e-07
MXP21 net108 nmset net136 VNW p12 l=1.3e-07 w=2.3e-07
MXP20 VDD s net136 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRX1MTR Q QN VDD VNW VPW VSS CK D RN SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm c XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MXN2 m NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MXN3 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MXN8 bm cn net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN7 NSN s net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm cn XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net_NRN NRN VDD VNW p12 l=1.3e-07 w=4.9e-07
MXP6 m pm net_NRN VNW p12 l=1.3e-07 w=3.6e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MXP7 bm c net75 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net_NRN s net75 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSRX2MTR Q QN VDD VNW VPW VSS CK D RN SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNOE pm c XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MXN2 m NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MXN3 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MXN4 bm cn net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 NSN s net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPOEN pm cn XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net_NRN NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 m pm net_NRN VNW p12 l=1.3e-07 w=4.4e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.4e-07
MXP7 bm c net75 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net_NRN s net75 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSRX4MTR Q QN VDD VNW VPW VSS CK D RN SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=2.5e-07
mXI4_MXNOE pm c XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.9e-07
mX_g5_MXNA1 NRN RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 m pm NSN VPW n12 l=1.3e-07 w=3e-07
MXN2 m NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=4.7e-07
MXN3 bm NRN NSN VPW n12 l=1.3e-07 w=1.9e-07
MXN4 bm cn net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN8 NSN s net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN6 NSN SN VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=3e-07
mXI4_MXPOEN pm cn XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.2e-07
mX_g5_MXPA1 NRN RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP2 net_NRN NRN VDD VNW p12 l=1.3e-07 w=6.9e-07
MXP6 m pm net_NRN VNW p12 l=1.3e-07 w=4.4e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=4.7e-07
MXP7 bm c net75 VNW p12 l=1.3e-07 w=2.3e-07
MXP9 net_NRN s net75 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSX1MTR Q QN VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 m pm BSN VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=1.9e-07
MXN1 bm cn net134 VPW n12 l=1.3e-07 w=1.8e-07
MXN4 BSN s net134 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 BSN SN VSS VPW n12 l=1.3e-07 w=4e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=2.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=2.4e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP7 bm c net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP6 VDD s net73 VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFSX2MTR Q QN VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
MXN0 m pm BSN VPW n12 l=1.3e-07 w=2.1e-07
MXN0_2 m pm BSN VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
MXN1 bm cn net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN4 BSN s net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN SN VSS VPW n12 l=1.3e-07 w=5.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=5.1e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=5.1e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.7e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=3.4e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=3.1e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm c net73 VNW p12 l=1.3e-07 w=1.5e-07
MXP6 VDD s net73 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFSX4MTR Q QN VDD VNW VPW VSS CK D SN
mX_g3_MXNA1 X_g3_n1 D VSS VPW n12 l=1.3e-07 w=2e-07
mX_g3_MXNOE pm cn X_g3_n1 VPW n12 l=1.3e-07 w=2e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
MXN0 m pm BSN VPW n12 l=1.3e-07 w=3.3e-07
MXN0_2 m pm BSN VPW n12 l=1.3e-07 w=3.3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=2.1e-07
mXI36_MXNOE bm c m VPW n12 l=1.3e-07 w=5.2e-07
MXN1 bm cn net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN4 BSN s net134 VPW n12 l=1.3e-07 w=1.5e-07
MXN3 BSN SN VSS VPW n12 l=1.3e-07 w=1.08e-06
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g0_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g0_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g3_MXPA1 X_g3_p1 D VDD VNW p12 l=1.3e-07 w=5.6e-07
mX_g3_MXPOEN pm c X_g3_p1 VNW p12 l=1.3e-07 w=5.6e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.4e-07
MXP0 m pm VDD VNW p12 l=1.3e-07 w=6.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5.9e-07
mXI36_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.2e-07
MXP1 m SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 bm SN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP8 bm c net73 VNW p12 l=1.3e-07 w=1.5e-07
MXP6 VDD s net73 VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g0_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g0_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFTRX1MTR Q QN VDD VNW VPW VSS CK D RN
MXN4 net129 RN VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net132 D net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 pm cn net132 VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=3.1e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=2.8e-07
mXI4_MXNOE bm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g11_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=3.6e-07
MXP4 net62 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 pm c net62 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.4e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=5.6e-07
mXI4_MXPOEN bm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g11_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFTRX2MTR Q QN VDD VNW VPW VSS CK D RN
MXN6 net129 RN VSS VPW n12 l=1.3e-07 w=2.6e-07
MXN5 net132 D net129 VPW n12 l=1.3e-07 w=2.6e-07
MXN1 pm cn net132 VPW n12 l=1.3e-07 w=2.6e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.1e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=4e-07
mXI4_MXNOE bm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g11_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 net62 RN VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=2.6e-07
MXP5 pm c net62 VNW p12 l=1.3e-07 w=2.6e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=5.7e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=8.1e-07
mXI4_MXPOEN bm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g11_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFTRX4MTR Q QN VDD VNW VPW VSS CK D RN
MXN8 net129 RN VSS VPW n12 l=1.3e-07 w=5e-07
MXN7 net132 D net129 VPW n12 l=1.3e-07 w=5e-07
MXN1 pm cn net132 VPW n12 l=1.3e-07 w=5e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNOE pm c XI3_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI3_MXNA1 XI3_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.3e-07
mX_g5_MXNA1_2 m pm VSS VPW n12 l=1.3e-07 w=4e-07
mXI47_MXNOE bm c m VPW n12 l=1.3e-07 w=8e-07
mXI4_MXNOE bm cn XI4_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI4_MXNA1 XI4_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g1_MXNA1 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 QN bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g11_MXNA1 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g11_MXNA1_2 Q s VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 net62 RN VDD VNW p12 l=1.3e-07 w=2.5e-07
MXP0 net62 D VDD VNW p12 l=1.3e-07 w=5.1e-07
MXP6 pm c net62 VNW p12 l=1.3e-07 w=5.1e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=8.6e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI3_MXPOEN pm cn XI3_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI3_MXPA1 XI3_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=3.6e-07
mX_g5_MXPA1_2 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_3 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mX_g5_MXPA1_4 m pm VDD VNW p12 l=1.3e-07 w=4e-07
mXI47_MXPOEN bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI47_MXPOEN_2 bm cn m VNW p12 l=1.3e-07 w=7.2e-07
mXI4_MXPOEN bm c XI4_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI4_MXPA1 XI4_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g1_MXPA1 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 QN bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g11_MXPA1 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g11_MXPA1_2 Q s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFX1MTR Q QN VDD VNW VPW VSS CK D
mXI14_MXNA1 XI14_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNOE pm cn XI14_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI12_MXNOE nm c XI12_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI11_MXNOE nm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mXI14_MXPA1 XI14_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI14_MXPOEN pm c XI14_p1 VNW p12 l=1.3e-07 w=3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI12_MXPOEN nm cn XI12_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI11_MXPOEN nm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT DFFX2MTR Q QN VDD VNW VPW VSS CK D
mXI14_MXNA1 XI14_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNOE pm cn XI14_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=4e-07
mXI12_MXNOE nm c XI12_n1 VPW n12 l=1.3e-07 w=4e-07
mXI11_MXNOE nm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1 XI14_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI14_MXPOEN pm c XI14_p1 VNW p12 l=1.3e-07 w=3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=4.9e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=4.9e-07
mXI12_MXPOEN nm cn XI12_p1 VNW p12 l=1.3e-07 w=4.9e-07
mXI11_MXPOEN nm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT DFFX4MTR Q QN VDD VNW VPW VSS CK D
mXI14_MXNA1 XI14_n1 D VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI14_MXNOE pm cn XI14_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 m VSS VPW n12 l=1.3e-07 w=5.8e-07
mXI12_MXNOE nm c XI12_n1 VPW n12 l=1.3e-07 w=5.8e-07
mXI11_MXNOE nm cn XI11_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI11_MXNA1 XI11_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=3.5e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mXI14_MXPA1 XI14_p1 D VDD VNW p12 l=1.3e-07 w=3e-07
mXI14_MXPOEN pm c XI14_p1 VNW p12 l=1.3e-07 w=3e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g14_MXPA1_2 cn CK VDD VNW p12 l=1.3e-07 w=3.1e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.7e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI12_MXPA1 XI12_p1 m VDD VNW p12 l=1.3e-07 w=6.6e-07
mXI12_MXPOEN nm cn XI12_p1 VNW p12 l=1.3e-07 w=6.6e-07
mXI11_MXPOEN nm c XI11_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI11_MXPA1 XI11_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=4.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends



.SUBCKT EDFFHQX1MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 VSS s net104 VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=2.3e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=3.6e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=3.6e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.5e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=4e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=3e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 nmsi E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=4.5e-07
MXP0 cn c net053 VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=6.3e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=4.4e-07
MXP2 pm nmsi net047 VNW p12 l=1.3e-07 w=4.4e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=7.9e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT EDFFHQX2MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=3.2e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 VSS s net104 VPW n12 l=1.3e-07 w=1.8e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=2e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=2.8e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=5.1e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.2e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.6e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=3.9e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=3.9e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 nmsi E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=4.5e-07
MXP0 cn c net053 VNW p12 l=1.3e-07 w=4.5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=8e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 pm nmsi net047 VNW p12 l=1.3e-07 w=6.2e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFHQX4MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=2.3e-07
MXN3 VSS s net104 VPW n12 l=1.3e-07 w=2.3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=5.1e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmsi E net73 VNW p12 l=1.3e-07 w=2.8e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=5e-07
MXP4 cn c net053 VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 pm nmsi net047 VNW p12 l=1.3e-07 w=6.2e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFHQX8MTR Q VDD VNW VPW VSS CK D E
mX_g13_MXNA1 nmin D VSS VPW n12 l=1.3e-07 w=5.7e-07
MX_t8 nmsi E nmin VPW n12 l=1.3e-07 w=3.2e-07
mX_g6_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t45 nmsi nmen net104 VPW n12 l=1.3e-07 w=2.3e-07
MXN3 VSS s net104 VPW n12 l=1.3e-07 w=2.3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3.3e-07
mX_g14_MXNA1 net132 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net132 VSS VPW n12 l=1.3e-07 w=4.6e-07
MXN2 VSS cn net98 VPW n12 l=1.3e-07 w=1.8e-07
MX_t2 pm nmsi net98 VPW n12 l=1.3e-07 w=5.1e-07
mXI5_MXNOE pm c XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=6.9e-07
mXI6_MXNOE bm cn XI6_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI6_MXNA1 XI6_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g13_MXPA1 nmin D VDD VNW p12 l=1.3e-07 w=7e-07
MX_t9 nmin nmen nmsi VNW p12 l=1.3e-07 w=7e-07
mX_g6_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP5 nmsi E net73 VNW p12 l=1.3e-07 w=2.8e-07
MX_t47 VDD s net73 VNW p12 l=1.3e-07 w=2.8e-07
mX_g14_MXPA1 net132 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net053 VNW p12 l=1.3e-07 w=5e-07
MXP4 cn c net053 VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c net132 VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t3i2 net047 c VDD VNW p12 l=1.3e-07 w=6.2e-07
MXP3 pm nmsi net047 VNW p12 l=1.3e-07 w=6.2e-07
mXI5_MXPOEN pm cn XI5_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI5_MXPA1 XI5_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI6_MXPOEN bm c XI6_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI6_MXPA1 XI6_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFTRX1MTR Q QN VDD VNW VPW VSS CK D E RN
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net122 s net140 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net122 nmen net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net107 E net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net140 D net107 VPW n12 l=1.3e-07 w=1.8e-07
MX_t3 net106 RN VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t19 pm cn net140 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI11_MXNOE bnm c XI11_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI5_MXNOE bnm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bnm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 net77 s net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 VDD nmen net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net76 D net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 VDD RN net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net77 c pm VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI11_MXPA1 XI11_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI11_MXPOEN bnm cn XI11_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI5_MXPOEN bnm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bnm VDD VNW p12 l=1.3e-07 w=6.4e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.4e-07
.ends


.SUBCKT EDFFTRX2MTR Q QN VDD VNW VPW VSS CK D E RN
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net122 s net140 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net122 nmen net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net107 E net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net140 D net107 VPW n12 l=1.3e-07 w=1.8e-07
MX_t3 net106 RN VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t19 pm cn net140 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 m VSS VPW n12 l=1.3e-07 w=3.9e-07
mXI11_MXNOE bnm c XI11_n1 VPW n12 l=1.3e-07 w=3.9e-07
mXI5_MXNOE bnm cn XI5_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI5_MXNA1 XI5_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g1_MXNA1 Q bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 net77 s net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 VDD nmen net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net76 D net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 VDD RN net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net77 c pm VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI11_MXPA1 XI11_p1 m VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI11_MXPOEN bnm cn XI11_p1 VNW p12 l=1.3e-07 w=5.2e-07
mXI5_MXPOEN bnm c XI5_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI5_MXPA1 XI5_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=2.8e-07
mX_g1_MXPA1 Q bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFTRX4MTR Q QN VDD VNW VPW VSS CK D E RN
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.4e-07
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net122 s net140 VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net122 nmen net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net107 E net106 VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net140 D net107 VPW n12 l=1.3e-07 w=1.8e-07
MX_t3 net106 RN VSS VPW n12 l=1.3e-07 w=1.7e-07
MX_t19 pm cn net140 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNOE pm c XI15_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI15_MXNA1 XI15_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI11_MXNA1 XI11_n1 m VSS VPW n12 l=1.3e-07 w=6.3e-07
mXI11_MXNOE bnm c XI11_n1 VPW n12 l=1.3e-07 w=6.3e-07
mXI5_MXNOE bnm cn XI5_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI5_MXNA1 XI5_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bnm VSS VPW n12 l=1.3e-07 w=5.3e-07
mX_g1_MXNA1 Q bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bnm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5.7e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP3 net77 s net73 VNW p12 l=1.3e-07 w=2.3e-07
MXP2 VDD E net73 VNW p12 l=1.3e-07 w=2.3e-07
MX_t5 VDD nmen net76 VNW p12 l=1.3e-07 w=2.3e-07
MXP0 net76 D net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP1 VDD RN net77 VNW p12 l=1.3e-07 w=2.3e-07
MXP4 net77 c pm VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPOEN pm cn XI15_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI15_MXPA1 XI15_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.9e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI11_MXPA1 XI11_p1 m VDD VNW p12 l=1.3e-07 w=8.2e-07
mXI11_MXPOEN bnm cn XI11_p1 VNW p12 l=1.3e-07 w=8.2e-07
mXI5_MXPOEN bnm c XI5_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI5_MXPA1 XI5_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bnm VDD VNW p12 l=1.3e-07 w=6.5e-07
mX_g1_MXPA1 Q bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bnm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFX1MTR Q QN VDD VNW VPW VSS CK D E
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net120 s net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net120 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net123 E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net129 D net123 VPW n12 l=1.3e-07 w=1.8e-07
MX_t19 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=2.8e-07
mXI1_MXNOE nm c XI1_n1 VPW n12 l=1.3e-07 w=2.8e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=3.6e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net38 s net36 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 VDD E net36 VNW p12 l=1.3e-07 w=3.8e-07
MX_t5 VDD nmen net39 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net39 D net38 VNW p12 l=1.3e-07 w=3.8e-07
MXP2 net38 c pm VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=3.4e-07
mXI1_MXPOEN nm cn XI1_p1 VNW p12 l=1.3e-07 w=3.4e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT EDFFX2MTR Q QN VDD VNW VPW VSS CK D E
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net120 s net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net120 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net123 E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net129 D net123 VPW n12 l=1.3e-07 w=1.8e-07
MX_t19 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=4.3e-07
mXI1_MXNOE nm c XI1_n1 VPW n12 l=1.3e-07 w=4.3e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=2.5e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net38 s net36 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 VDD E net36 VNW p12 l=1.3e-07 w=3.8e-07
MX_t5 VDD nmen net39 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net39 D net38 VNW p12 l=1.3e-07 w=3.8e-07
MXP2 net38 c pm VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=5e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=5.2e-07
mXI1_MXPOEN nm cn XI1_p1 VNW p12 l=1.3e-07 w=5.2e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=3e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT EDFFX4MTR Q QN VDD VNW VPW VSS CK D E
mX_g8_MXNA1 nmen E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN3 net120 s net129 VPW n12 l=1.3e-07 w=1.8e-07
MXN0 net120 nmen VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN1 net123 E VSS VPW n12 l=1.3e-07 w=1.8e-07
MXN2 net129 D net123 VPW n12 l=1.3e-07 w=1.8e-07
MX_t19 pm cn net129 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNOE pm c XI0_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI0_MXNA1 XI0_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g5_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g14_MXNA1 cn CK VSS VPW n12 l=1.3e-07 w=2.2e-07
mX_g10_MXNA1 c cn VSS VPW n12 l=1.3e-07 w=1.8e-07
mXI1_MXNA1 XI1_n1 m VSS VPW n12 l=1.3e-07 w=6.4e-07
mXI1_MXNOE nm c XI1_n1 VPW n12 l=1.3e-07 w=6.4e-07
mXI2_MXNOE nm cn XI2_n1 VPW n12 l=1.3e-07 w=1.5e-07
mXI2_MXNA1 XI2_n1 s VSS VPW n12 l=1.3e-07 w=1.5e-07
mX_g2_MXNA1 s nm VSS VPW n12 l=1.3e-07 w=4.1e-07
mX_g1_MXNA1 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q nm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g9_MXNA1_2 QN s VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g8_MXPA1 nmen E VDD VNW p12 l=1.3e-07 w=2.3e-07
MXP1 net38 s net36 VNW p12 l=1.3e-07 w=3.8e-07
MXP0 VDD E net36 VNW p12 l=1.3e-07 w=3.8e-07
MX_t5 VDD nmen net39 VNW p12 l=1.3e-07 w=3.8e-07
MXP3 net39 D net38 VNW p12 l=1.3e-07 w=3.8e-07
MXP2 net38 c pm VNW p12 l=1.3e-07 w=3.8e-07
mXI0_MXPOEN pm cn XI0_p1 VNW p12 l=1.3e-07 w=2.2e-07
mXI0_MXPA1 XI0_p1 m VDD VNW p12 l=1.3e-07 w=2.2e-07
mX_g5_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=2.7e-07
mX_g14_MXPA1 cn CK VDD VNW p12 l=1.3e-07 w=6.2e-07
mX_g10_MXPA1 c cn VDD VNW p12 l=1.3e-07 w=5e-07
mXI1_MXPA1 XI1_p1 m VDD VNW p12 l=1.3e-07 w=7.3e-07
mXI1_MXPOEN nm cn XI1_p1 VNW p12 l=1.3e-07 w=7.3e-07
mXI2_MXPOEN nm c XI2_p1 VNW p12 l=1.3e-07 w=1.5e-07
mXI2_MXPA1 XI2_p1 s VDD VNW p12 l=1.3e-07 w=1.5e-07
mX_g2_MXPA1 s nm VDD VNW p12 l=1.3e-07 w=5e-07
mX_g1_MXPA1 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q nm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g9_MXPA1_2 QN s VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MDFFHQX1MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=2.1e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=2.1e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=2.1e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=2.1e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=2.2e-07
MXN0 net135 cn VSS VPW n12 l=1.3e-07 w=3.3e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=3.3e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=4.2e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=3.7e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t9 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=2.6e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=2.6e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=3e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=3e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=4.2e-07
MXP0 cn c net50 VNW p12 l=1.3e-07 w=4.2e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=6.1e-07
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=4e-07
MXP1 pm nmsi net61 VNW p12 l=1.3e-07 w=4e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=7.3e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=7.3e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=6.2e-07
.ends


.SUBCKT MDFFHQX2MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=3.1e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=3.1e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=3e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=3e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=1.9e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=2.3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=2.7e-07
MXN1 net135 cn VSS VPW n12 l=1.3e-07 w=4.8e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=4.8e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=5.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=3.7e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=3.7e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=4.4e-07
MXP2 cn c net50 VNW p12 l=1.3e-07 w=4.4e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=7.6e-07
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=5.9e-07
MXP5 pm nmsi net61 VNW p12 l=1.3e-07 w=5.9e-07
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=9.8e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=9.8e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MDFFHQX4MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=5e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN2 net135 cn VSS VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=5.6e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.4e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net50 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net61 VNW p12 l=1.3e-07 w=1.01e-06
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends


.SUBCKT MDFFHQX8MTR Q VDD VNW VPW VSS CK D0 D1 S0
MX_t8 nmsi S0 nmin1 VPW n12 l=1.3e-07 w=5.5e-07
mX_g13_MXNA1 nmin1 D1 VSS VPW n12 l=1.3e-07 w=5.5e-07
mX_g6_MXNA1 nms0 S0 VSS VPW n12 l=1.3e-07 w=1.8e-07
MX_t11 nmsi nms0 nmin0 VPW n12 l=1.3e-07 w=4.9e-07
mX_g16_MXNA1 nmin0 D0 VSS VPW n12 l=1.3e-07 w=3.6e-07
MX_t13 cn CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g14_MXNA1 net109 CK VSS VPW n12 l=1.3e-07 w=3e-07
mX_g10_MXNA1 c net109 VSS VPW n12 l=1.3e-07 w=4.5e-07
MXN2 net135 cn VSS VPW n12 l=1.3e-07 w=5.6e-07
MX_t2 pm nmsi net135 VPW n12 l=1.3e-07 w=5.6e-07
mXI13_MXNOE pm c XI13_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI13_MXNA1 XI13_n1 m VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g7_MXNA1 m pm VSS VPW n12 l=1.3e-07 w=6.9e-07
MX_t0 bm c m VPW n12 l=1.3e-07 w=5.3e-07
mXI12_MXNOE bm cn XI12_n1 VPW n12 l=1.3e-07 w=1.8e-07
mXI12_MXNA1 XI12_n1 s VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g2_MXNA1 s bm VSS VPW n12 l=1.3e-07 w=1.8e-07
mX_g1_MXNA1 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_2 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_3 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
mX_g1_MXNA1_4 Q bm VSS VPW n12 l=1.3e-07 w=7.1e-07
MXP4 nmin1 nms0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g13_MXPA1 nmin1 D1 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g6_MXPA1 nms0 S0 VDD VNW p12 l=1.3e-07 w=2.3e-07
MX_t10 nmin0 S0 nmsi VNW p12 l=1.3e-07 w=6.8e-07
mX_g16_MXPA1 nmin0 D0 VDD VNW p12 l=1.3e-07 w=6.8e-07
mX_g14_MXPA1 net109 CK VDD VNW p12 l=1.3e-07 w=3e-07
MX_t22 VDD CK net50 VNW p12 l=1.3e-07 w=6.5e-07
MXP6 cn c net50 VNW p12 l=1.3e-07 w=6.5e-07
mX_g10_MXPA1 c net109 VDD VNW p12 l=1.3e-07 w=1.02e-06
MX_t3i2 net61 c VDD VNW p12 l=1.3e-07 w=1.01e-06
MXP7 pm nmsi net61 VNW p12 l=1.3e-07 w=1.01e-06
mXI13_MXPOEN pm cn XI13_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI13_MXPA1 XI13_p1 m VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g7_MXPA1 m pm VDD VNW p12 l=1.3e-07 w=8.9e-07
MX_t1 m cn bm VNW p12 l=1.3e-07 w=8.8e-07
mXI12_MXPOEN bm c XI12_p1 VNW p12 l=1.3e-07 w=2.3e-07
mXI12_MXPA1 XI12_p1 s VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g2_MXPA1 s bm VDD VNW p12 l=1.3e-07 w=2.3e-07
mX_g1_MXPA1 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_2 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_3 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
mX_g1_MXPA1_4 Q bm VDD VNW p12 l=1.3e-07 w=8.7e-07
.ends
