* 
* No part of this file can be released without the consent of SMIC.
*
* Note: SMIC recommends that users set VNTOL=1E-9 at .option for more smooth convergence, and please use Star-HSPICE version 2008.09.sp1 or more advance version to run gate current.
******************************************************************************************
* 0.11um Mixed Signal 1P8M with MIM Salicide 1.2V/3.3V RF SPICE Model (for HSPICE only)  *
******************************************************************************************
*
* Release version    : 1.14
*
* Release date       : 03/30/2016
*
* Simulation tool    : Synopsys Star-HSPICE version 2008.09.sp1
*
* Model type         :
*   MOSFET           : HSPICE Level 49(BSIM3V3.2)
*   Junction Diode   : HSPICE Level 3
* 
* Model and subcircuit name         :
*   MOSFET           :
*        *--------------------------------------------------*
*        |     MOSFET model   |     1.2V     |     3.3V     |
*        |==================================================|
*        |        NMOS        |  n12_ckt_rf  |  n33_ckt_rf  |
*        *--------------------------------------------------*
*        |      DNW MOS       | dnw12_ckt_rf | dnw33_ckt_rf |
*        *--------------------------------------------------*
*        |        PMOS        |  p12_ckt_rf  |  p33_ckt_rf  |
*        *--------------------------------------------------*
*
*************************
* 1.2V RF NMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt n12_ckt_rf 1 2 3 4 lr=l wr=w nf=finger sar=sa sbr=sb mr=m mismod=0 
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+atox_n12_rf=1.7e-11
+axl_n12_rf=3e-9
+lef=lr
+wef='wr*nf'
+dtox_n12_mis_rf     = 'atox_n12_rf*1/sqrt(lef*wef*1e12*mr)*sigma_mis_a_rf*mismod'
+dxl_n12_mis_rf     = 'axl_n12_rf*1/sqrt(wef*1e6*mr)*sigma_mis_b_rf*mismod'
+Rg_rf        = 'max((((-60.55*pwr((wr*0.9*1e+6),2.021)+1614)*(lr*0.9*1e+6)+(914.8*pwr((wr*0.9*1e+6),-1.604)+263.4))*pwr((nf+4),-1.5)+0.5),1e-6)'
+Cgd_rf	= 'max(((7.357e-15*pwr((wr*1e+6),0.7853)-2.388e-15)*(lr*1e+6)+(1.602e-18*exp(wr*1e+6*1.2)+0.2191e-15))*nf,1e-18)'
+Cgs_rf	= 1e-16
+Cds_rf       = 'max((((0.2441e-15*pwr((wr*1e+6),1.33)+27.75e-18)*pwr((10*lr*1e+6),-1)+(4.609e-18*exp(wr*1e+6*0.895)-0.05129e-15))*pwr(nf,1.2))*0.75,1e-18)'
+Rds_rf       = 220
+Rsub1_rf     = 10
+Rsub2_rf     = '((12.15e+3*pwr((wr*1e+6),-2.0)+1.997e+3)*pwr((10*lr*1e+6),-1)+(-10.78*pwr((wr*1e+6),3.38)+2.857e+3))*pwr((nf+2),-1)'
+Rsub3_rf     = '((12.15e+3*pwr((wr*1e+6),-2.0)+1.997e+3)*pwr((10*lr*1e+6),-1)+(-10.78*pwr((wr*1e+6),3.38)+2.857e+3))*pwr((nf+2),-1)'
+Djdb_AREA_rf = 'int(0.5*(nf+1))*(wr*(0.42e-6-2*0.065e-6))'
+Djdb_PJ_rf   = 'int(0.5*(nf+1))*(2*(0.42e-6-2*0.065e-6)+2*wr*4.6827)'
+Djsb_AREA_rf = 'int(0.5*nf+1)*(wr*(0.42e-6-2*0.065e-6))'
+Djsb_PJ_rf   = 'int(0.5*nf+1)*(2*(0.42e-6-2*0.065e-6)+2*wr*4.6827)'
*****************************************
Lgate       2 20 1p m=mr
Rgate       20 21 Rg_rf m=mr
Cgd_ext     20 11 'Cgd_rf*pwr((((-14.20*pwr((wr*1e+6),-0.302)+20.85)*pwr((lr*1e+6),0.8)+(0.9846*pwr((wr*1e+6),-0.6706)-0.7046))+pwr((((-0.02295*pwr((wr*1e+6),0.3188)+0.05779)*pwr((lr*1e+6),-2)+(0.5343*pwr((wr*1e+6),-1.7)+0.9511))+2*exp(((V(2,3)*-2.004+V(1,3))*2.31)*-1)),-1)),-1)' m=mr
Cgs_ext     20 31 'Cgs_rf+(1e-16+(0.26e-15*nf*(wr*1e+6))*pwr((1+exp((V(2,3)-0.542)*11.74)),-1))' m=mr
Rds         11 15 Rds_rf m=mr
Cds_ext     15 31 Cds_rf m=mr
Ldrain       1 11 1p m=mr
Lsource      3 31 1p m=mr
*****************************************
Djdb  12 11
+ ndio12_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
+ m     = mr
***
Djsb  32 31
+ ndio12_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
+ m     = mr
*****************************************
Rsub1      41  4  Rsub1_rf m=mr
Rsub2      41  12 Rsub2_rf m=mr
Rsub3      41  32 Rsub3_rf m=mr
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 n12_rf L=lr W='wr*nf' m=mr AD = 0 AS = 0 PD = 0 PS = 0 sa=sar sb=sbr 
* MOS Model
.MODEL  N12_RF  NMOS  
+level = 49
**************************************************************
*               MODEL FLAG PARAMETERS 
**************************************************************
+version = 3.24            lmin    = 1.3e-007        lmax    = 1e-005        
+wmin    = 1.5e-007        wmax    = 0.0001          binunit = 2             
+mobmod  = 1               capmod  = 3               nqsmod  = 0             
+stimod  = 1             
**************************************************************
*               GENERAL MODEL PARAMETERS 
**************************************************************
+tnom    = 25              tox     = '2.58e-009+dtox_n12_rf+dtox_n12_mis_rf'      toxm    = 2.58e-009     
+wint    = 0               lint    = 2.25e-008       dlc     = 2.33e-009   
+dwc     = -2.8e-008       hdif    = 1.25e-007       ldif    = 6.5e-008      
+xl      = '1.26e-8+dxl_n12_rf+dxl_n12_mis_rf'             xw      = '0+dxw_n12_rf'  xj      = 1.78e-007     
+ngate   = 1.176e+021      ll      = -8.5937e-016    wl      = -6.509098e-015
+lln     = 1.0204          wln     = 0.835           lw      = 9.069495e-017 
+ww      = -1e-014         lwn     = 0.989           wwn     = 0.892         
+lwl     = -4.8223e-022    wwl     = -6.2e-020       llc     = 0             
+wlc     = 0               lwc     = 0               wwc     = 0             
+lwlc    = 0               wwlc    = 0               xpart   = 0             
+igcmod  = 1               igbmod  = 1             
**************************************************************
*               EXPERT PARAMETERS 
**************************************************************
+vth0    = '0.275+dvth_n12_rf'  lvth0   = 3e-009          wvth0   = -1.6183e-008  
+pvth0   = '2.848e-015+dpvth0_n12_rf'  k1      = 0.51477         lk1     = -7.6162e-009  
+k2      = -0.0065         k3      = '6+dk3_n12_rf'  k3b     = 0             
+nlx     = '7.4e-008+dnlx_n12_rf'  w0      = 2e-006          dvt0    = 0.43          
+ldvt0   = 1.2e-007        dvt1    = 1.0528          dvt2    = -0.05         
+dvt0w   = 0.71578         dvt1w   = 975990          dvt2w   = -0.196        
+nch     = 2.416e+017      voff    = -0.11342        nfactor = 2             
+cdsc    = 0.001           cdscb   = 0         cdscd   = 0.001         
+cit     = 0.00065674      alpha0  = 2.1e-008        alpha1  = 0.28          
+beta0   = 11.25           eta0    = 0.04872         leta0   = 2.0135e-009   
+peta0   = 1.08e-015       etab    = -0.075924       dsub    = 0.56          
+u0      = '0.02355+du0_n12_rf'  lu0     = '0+dlu0_n12_rf'  wu0     = 2e-011        
+pu0     = '-5.1e-017+dpu0_n12_rf'  ua      = -1.2885e-009    lua     = -5.6e-018     
+wua     = 1.3e-016        ub      = 1.6248e-018     uc      = 1.4694e-010   
+wuc     = 5e-018          prwg    = 0               prwb    = 0             
+wr      = 0.95            rdsw    = 60.027          a0      = 1.25          
+ags     = 0.42302         a1      = 0               a2      = 0.99          
+b0      = -4.4e-008       lb0     = 3e-014          b1      = 0             
+vsat    = 77186           lvsat   = '0+dlvsat_n12_rf'  pvsat   = -2e-010       
+keta    = 0.006           lketa   = 2.6e-009        wketa   = -1.3e-008     
+pketa   = 6.6e-016        delta   = 0.0032          dwg     = 4.6e-010      
+dwb     = 4.3383e-009     pclm    = 1.16            pdiblc1 = 0             
+pdiblc2 = 0.003956        pdiblcb = -0.001          drout   = 0.56          
+pvag    = -1e-010         pscbe1  = 8e+008          pscbe2  = 3.9002e-005   
+elm     = 5               agidl   = '0+dagidl_n12_rf'  wagidl  = -8.4985e-006  
+bgidl   = 2.3e+009        cgidl   = 0.5             egidl   = 0.8           
+aigbacc = 0.0136          bigbacc = 0.00171         cigbacc = 0.075         
+nigbacc = 1               aigbinv = 0.0111          bigbinv = 0.000949      
+cigbinv = 0.006           eigbinv = 1.1             nigbinv = 3             
+aigc    = 0.010962        bigc    = 0.00171         cigc    = 0.075         
+nigc    = 1               pigcd   = 1               aigsd   = 0.011015      
+bigsd   = 0.0011799       cigsd   = 0.075           poxedge = 1             
+ntox    = 1             
**************************************************************
*               CAPACITANCE PARAMETERS 
**************************************************************
+acde    = 0.50083         moin    = 24.39           noff    = 1.9644        
+voffcv  = 0.062777        cgbo    = 0               cgso    = 1e-24
+cgdo    = 1e-24  cgsl    = 1e-24       cf      = 0             
+ckappa  = 0.6           
+clc = 1e-18
**************************************************************
*               TEMPERATURE PARAMETERS 
**************************************************************
+kt1     = -0.25           wkt1    = 3e-009          pkt1    = 1e-015        
+kt1l    = 1e-010          kt2     = 0               ute     = -1.5          
+lute    = 2.5557e-008     wute    = 3e-008          pute    = 1e-015        
+ua1     = 1.386e-009      lua1    = 5.001e-019      pua1    = -1.0762e-023  
+ub1     = -1.285e-018     uc1     = -9.3847e-011    luc1    = 1.5e-017      
+puc1    = 1.6646e-026     prt     = 0               at      = 40000         
+pat     = -1.15e-009    
**************************************************************
*               NOISE PARAMETERS 
**************************************************************
+noia    = 9.3101e+019     noib    = 46000           noic    = -1.2e-013     
+em      = 13865000        ef      = 0.88            noimod  = 2             
**************************************************************
*               DIODE PARAMETERS 
**************************************************************
+rsh     = 6.45            js      = 1.06e-006       jsw     = 1.5e-010   
+cj      = 0  mj      = 0.458           cjsw    = 0
+mjsw    = 0.593           cjswg   = 0  mjswg   = 0.472        
+pb      = 0.791           pbsw    = 0.955           pbswg   = 0.915          
+rd      = 0               rdc     = 1.35            rs      = 0             
+rsc     = 1.35            xti     = 3               tpb     = 0.00112       
+tpbsw   = 0.000924        tpbswg  = 0.00159         tcj     = 0.000759      
+tcjsw   = 0.000585        tcjswg  = 0.000668        acm     = 12            
+calcacm = 1               nj      = 1.083         
**************************************************************
*               STRESS PARAMETERS 
**************************************************************
+saref   = 2.25e-006       sbref   = 2.25e-006       wlod    = 0             
+kvth0   = 1.2e-008        lkvth0  = 1.7e-007        wkvth0  = 3.4e-007      
+pkvth0  = 0               llodvth = 1               wlodvth = 1             
+stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = -1.1e-007       lku0    = 1.16e-006       wku0    = 0             
+pku0    = 0               llodku0 = 1               wlodku0 = 1             
+kvsat   = -0.42           steta0  = -2.4e-008       tku0    = 0         
*
***********************************************************************************
*                            1.2V N+/PWELL DIODE MODEL                            *
***********************************************************************************
*
.MODEL NDIO12_RF D
+LEVEL    = 3                   JS       = 1.06E-06 JSW      = 1.00E-15            
+N        = 1.083   RS       = 1.0E-010              IK       = 1.0E+21           
+IKR      = 2.78E+05            BV       = 10.25                 IBV      = 277.8             
+TRS      = 1.00E-05            EG       = 1.16                  TREF     = 25.0                
+XTI      = 3.0                 TLEV     = 1                     TLEVC    = 1
+CJ       = '1.315E-03+DCJ_N12_rf'
+CJSW     = '1.04E-10+DCJSW_N12_rf'
+MJ       = 0.458               PB       = 0.791               
+MJSW     = 0.593               PHP      = 0.955                   
+CTA      = 7.59E-04            CTP      = 5.85E-04              TPB      = 1.12E-03             
+TPHP     = 9.24E-04            FC       = 0                     FCS      = 0   
+AREA     = 3.60E-09            PJ       = 2.4E-04            
*
.ends n12_ckt_rf

***************************
* 1.2V RF DNWMOS Subcircuit
***************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt dnw12_ckt_rf 1 2 3 4 lr=l wr=w nf=finger sar=sa sbr=sb mr=m mismod=0 
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+atox_n12_rf=1.7e-11
+axl_n12_rf=3e-9
+lef=lr
+wef='wr*nf'
+dtox_n12_mis_rf     = 'atox_n12_rf*1/sqrt(lef*wef*1e12*mr)*sigma_mis_a_rf*mismod'
+dxl_n12_mis_rf     = 'axl_n12_rf*1/sqrt(wef*1e6*mr)*sigma_mis_b_rf*mismod'
+Rg_rf        = 'max((((-60.55*pwr((wr*0.9*1e+6),2.021)+1614)*(lr*0.9*1e+6)+(914.8*pwr((wr*0.9*1e+6),-1.604)+263.4))*pwr((nf+4),-1.5)+0.5),1e-6)'
+Cgd_rf	= 'max(((7.357e-15*pwr((wr*1e+6),0.7853)-2.388e-15)*(lr*1e+6)+(1.602e-18*exp(wr*1e+6*1.2)+0.2191e-15))*nf,1e-18)'
+Cgs_rf	= 1e-16
+Cds_rf       = 'max((((0.2441e-15*pwr((wr*1e+6),1.33)+27.75e-18)*pwr((10*lr*1e+6),-1)+(4.609e-18*exp(wr*1e+6*0.895)-0.05129e-15))*pwr(nf,1.2))*0.75,1e-18)'
+Rds_rf       = 220
+Rsub1_rf     = 10
+Rsub2_rf     = '((12.15e+3*pwr((wr*1e+6),-2.0)+1.997e+3)*pwr((10*lr*1e+6),-1)+(-10.78*pwr((wr*1e+6),3.38)+2.857e+3))*pwr((nf+2),-1)'
+Rsub3_rf     = '((12.15e+3*pwr((wr*1e+6),-2.0)+1.997e+3)*pwr((10*lr*1e+6),-1)+(-10.78*pwr((wr*1e+6),3.38)+2.857e+3))*pwr((nf+2),-1)'
+Djdb_AREA_rf = 'int(0.5*(nf+1))*(wr*(0.42e-6-2*0.065e-6))'
+Djdb_PJ_rf   = 'int(0.5*(nf+1))*(2*(0.42e-6-2*0.065e-6)+2*wr*4.6827)'
+Djsb_AREA_rf = 'int(0.5*nf+1)*(wr*(0.42e-6-2*0.065e-6))'
+Djsb_PJ_rf   = 'int(0.5*nf+1)*(2*(0.42e-6-2*0.065e-6)+2*wr*4.6827)'
*****************************************
Lgate       2 20 1p m=mr
Rgate       20 21 Rg_rf m=mr
Cgd_ext     20 11 'Cgd_rf*pwr((((-14.20*pwr((wr*1e+6),-0.302)+20.85)*pwr((lr*1e+6),0.8)+(0.9846*pwr((wr*1e+6),-0.6706)-0.7046))+pwr((((-0.02295*pwr((wr*1e+6),0.3188)+0.05779)*pwr((lr*1e+6),-2)+(0.5343*pwr((wr*1e+6),-1.7)+0.9511))+2*exp(((V(2,3)*-2.004+V(1,3))*2.31)*-1)),-1)),-1)' m=mr
Cgs_ext     20 31 'Cgs_rf+(1e-16+(0.26e-15*nf*(wr*1e+6))*pwr((1+exp((V(2,3)-0.542)*11.74)),-1))' m=mr
Rds         11 15 Rds_rf m=mr
Cds_ext     15 31 Cds_rf m=mr
Ldrain       1 11 1p m=mr
Lsource      3 31 1p m=mr
*****************************************
Djdb  12 11
+ ndio12_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
+ m     = mr
***
Djsb  32 31
+ ndio12_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
+ m     = mr
*****************************************
Rsub1      41  4  Rsub1_rf m=mr
Rsub2      41  12 Rsub2_rf m=mr
Rsub3      41  32 Rsub3_rf m=mr
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 dnw12_rf L=lr W='wr*nf' m=mr AD = 0 AS = 0 PD = 0 PS = 0 sa=sar sb=sbr  
* MOS Model
.MODEL  dnw12_rf  NMOS  
+level = 49
**************************************************************
*               MODEL FLAG PARAMETERS 
**************************************************************
+version = 3.24            lmin    = 1.3e-007        lmax    = 1e-005        
+wmin    = 1.5e-007        wmax    = 0.0001          binunit = 2             
+mobmod  = 1               capmod  = 3               nqsmod  = 0             
+stimod  = 1             
**************************************************************
*               GENERAL MODEL PARAMETERS 
**************************************************************
+tnom    = 25              tox     = '2.58e-009+dtox_n12_rf+dtox_n12_mis_rf'      toxm    = 2.58e-009     
+wint    = 0               lint    = 2.25e-008       dlc     = 2.33e-009   
+dwc     = -2.8e-008       hdif    = 1.25e-007       ldif    = 6.5e-008      
+xl      = '1.26e-8+dxl_n12_rf+dxl_n12_mis_rf'             xw      = '0+dxw_n12_rf'  xj      = 1.78e-007     
+ngate   = 1.176e+021      ll      = -8.5937e-016    wl      = -6.509098e-015
+lln     = 1.0204          wln     = 0.835           lw      = 9.069495e-017 
+ww      = -1e-014         lwn     = 0.989           wwn     = 0.892         
+lwl     = -4.8223e-022    wwl     = -6.2e-020       llc     = 0             
+wlc     = 0               lwc     = 0               wwc     = 0             
+lwlc    = 0               wwlc    = 0               xpart   = 0             
+igcmod  = 1               igbmod  = 1             
**************************************************************
*               EXPERT PARAMETERS 
**************************************************************
+vth0    = '0.275+dvth_n12_rf'  lvth0   = 3e-009          wvth0   = -1.6183e-008  
+pvth0   = '2.848e-015+dpvth0_n12_rf'  k1      = 0.51477         lk1     = -7.6162e-009  
+k2      = -0.0065         k3      = '6+dk3_n12_rf'  k3b     = 0             
+nlx     = '7.4e-008+dnlx_n12_rf'  w0      = 2e-006          dvt0    = 0.43          
+ldvt0   = 1.2e-007        dvt1    = 1.0528          dvt2    = -0.05         
+dvt0w   = 0.71578         dvt1w   = 975990          dvt2w   = -0.196        
+nch     = 2.416e+017      voff    = -0.11342        nfactor = 2             
+cdsc    = 0.001           cdscb   = 0         cdscd   = 0.001         
+cit     = 0.00065674      alpha0  = 2.1e-008        alpha1  = 0.28          
+beta0   = 11.25           eta0    = 0.04872         leta0   = 2.0135e-009   
+peta0   = 1.08e-015       etab    = -0.075924       dsub    = 0.56          
+u0      = '0.02355+du0_n12_rf'  lu0     = '0+dlu0_n12_rf'  wu0     = 2e-011        
+pu0     = '-5.1e-017+dpu0_n12_rf'  ua      = -1.2885e-009    lua     = -5.6e-018     
+wua     = 1.3e-016        ub      = 1.6248e-018     uc      = 1.4694e-010   
+wuc     = 5e-018          prwg    = 0               prwb    = 0             
+wr      = 0.95            rdsw    = 60.027          a0      = 1.25          
+ags     = 0.42302         a1      = 0               a2      = 0.99          
+b0      = -4.4e-008       lb0     = 3e-014          b1      = 0             
+vsat    = 77186           lvsat   = '0+dlvsat_n12_rf'  pvsat   = -2e-010       
+keta    = 0.006           lketa   = 2.6e-009        wketa   = -1.3e-008     
+pketa   = 6.6e-016        delta   = 0.0032          dwg     = 4.6e-010      
+dwb     = 4.3383e-009     pclm    = 1.16            pdiblc1 = 0             
+pdiblc2 = 0.003956        pdiblcb = -0.001          drout   = 0.56          
+pvag    = -1e-010         pscbe1  = 8e+008          pscbe2  = 3.9002e-005   
+elm     = 5               agidl   = '0+dagidl_n12_rf'  wagidl  = -8.4985e-006  
+bgidl   = 2.3e+009        cgidl   = 0.5             egidl   = 0.8           
+aigbacc = 0.0136          bigbacc = 0.00171         cigbacc = 0.075         
+nigbacc = 1               aigbinv = 0.0111          bigbinv = 0.000949      
+cigbinv = 0.006           eigbinv = 1.1             nigbinv = 3             
+aigc    = 0.010962        bigc    = 0.00171         cigc    = 0.075         
+nigc    = 1               pigcd   = 1               aigsd   = 0.011015      
+bigsd   = 0.0011799       cigsd   = 0.075           poxedge = 1             
+ntox    = 1             
**************************************************************
*               CAPACITANCE PARAMETERS 
**************************************************************
+acde    = 0.50083         moin    = 24.39           noff    = 1.9644        
+voffcv  = 0.062777        cgbo    = 0               cgso    = 1e-24
+cgdo    = 1e-24  cgsl    = 1e-24       cf      = 0             
+ckappa  = 0.6           
+clc = 1e-18
**************************************************************
*               TEMPERATURE PARAMETERS 
**************************************************************
+kt1     = -0.25           wkt1    = 3e-009          pkt1    = 1e-015        
+kt1l    = 1e-010          kt2     = 0               ute     = -1.5          
+lute    = 2.5557e-008     wute    = 3e-008          pute    = 1e-015        
+ua1     = 1.386e-009      lua1    = 5.001e-019      pua1    = -1.0762e-023  
+ub1     = -1.285e-018     uc1     = -9.3847e-011    luc1    = 1.5e-017      
+puc1    = 1.6646e-026     prt     = 0               at      = 40000         
+pat     = -1.15e-009    
**************************************************************
*               NOISE PARAMETERS 
**************************************************************
+noia    = 9.3101e+019     noib    = 46000           noic    = -1.2e-013     
+em      = 13865000        ef      = 0.88            noimod  = 2             
**************************************************************
*               DIODE PARAMETERS 
**************************************************************
+rsh     = 6.45            js      = 1.06e-006       jsw     = 1.5e-010   
+cj      = 0  mj      = 0.458           cjsw    = 0
+mjsw    = 0.593           cjswg   = 0  mjswg   = 0.472        
+pb      = 0.791           pbsw    = 0.955           pbswg   = 0.915          
+rd      = 0               rdc     = 1.35            rs      = 0             
+rsc     = 1.35            xti     = 3               tpb     = 0.00112       
+tpbsw   = 0.000924        tpbswg  = 0.00159         tcj     = 0.000759      
+tcjsw   = 0.000585        tcjswg  = 0.000668        acm     = 12            
+calcacm = 1               nj      = 1.083         
**************************************************************
*               STRESS PARAMETERS 
**************************************************************
+saref   = 2.25e-006       sbref   = 2.25e-006       wlod    = 0             
+kvth0   = 1.2e-008        lkvth0  = 1.7e-007        wkvth0  = 3.4e-007      
+pkvth0  = 0               llodvth = 1               wlodvth = 1             
+stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = -1.1e-007       lku0    = 1.16e-006       wku0    = 0             
+pku0    = 0               llodku0 = 1               wlodku0 = 1             
+kvsat   = -0.42           steta0  = -2.4e-008       tku0    = 0         
*
***********************************************************************************
*                            1.2V N+/PWELL DIODE MODEL                            *
***********************************************************************************
*
.MODEL NDIO12_RF D
+LEVEL    = 3                   JS       = 1.06E-06 JSW      = 1.00E-15            
+N        = 1.083   RS       = 1.0E-010              IK       = 1.0E+21           
+IKR      = 2.78E+05            BV       = 10.25                 IBV      = 277.8             
+TRS      = 1.00E-05            EG       = 1.16                  TREF     = 25.0                
+XTI      = 3.0                 TLEV     = 1                     TLEVC    = 1
+CJ       = '1.315E-03+DCJ_N12_rf'
+CJSW     = '1.04E-10+DCJSW_N12_rf'
+MJ       = 0.458               PB       = 0.791               
+MJSW     = 0.593               PHP      = 0.955                   
+CTA      = 7.59E-04            CTP      = 5.85E-04              TPB      = 1.12E-03             
+TPHP     = 9.24E-04            FC       = 0                     FCS      = 0   
+AREA     = 3.60E-09            PJ       = 2.4E-04            
*
.ends dnw12_ckt_rf
*************************
* 1.2V RF PMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt p12_ckt_rf 1 2 3 4 lr=l wr=w nf=finger sar=sa sbr=sb mr=1 mismod=0 
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+atox_p12_rf=2.85e-11
+axl_p12_rf=8e-10
+lef=lr 
+wef=wr
+dtox_p12_rf_mis='atox_p12_rf*1/sqrt(lef*wef*1e12*mr*nf)*sigma_mis_a_rf*mismod'
+dxl_p12_rf_mis='axl_p12_rf*1/sqrt(wef*1e6*mr*nf)*sigma_mis_b_rf*mismod'
+dtox_p12_rf_mismatch         = 'dtox_p12_rf+dtox_p12_rf_mis' 
+dxl_p12_rf_mismatch         = 'dxl_p12_rf+dxl_p12_rf_mis'              
+Rg_rf		= 'max((((-5341*pwr((wr*0.9*1e+6),0.2654)+9321)*(lr*0.9*1e+6)+(1160*pwr((wr*0.9*1e+6),-2.877)+231.1))*pwr((nf+4),-1.5)+1), 1e-6)'
+Cgd_rf	= 'max(((2.64850076E-16*wr*1e6+1.84365144E-16)*lr*1e6+(4.19497690E-16*wr*1e6+1.40715320E-16))*nf,1e-18)'
+Cgs_rf	= 'max(((-2.86095151E-18*wr*wr*1e12+1.03812351E-17*wr*1e6-1.87094266E-17)*lr*lr*1e12+(1.28779805E-17*wr*wr*1e12-7.55186057E-17*wr*1e6+6.57478360E-17)*lr*1e6+(-1.84418296E-18*wr*wr*1e12+1.01606428E-17*wr*1e6-8.75192944E-18))*nf*nf+((4.47990652E-16*wr*wr*1e12-2.66963228E-15*wr*1e6+3.98528199E-15)*lr*lr*1e12+(-3.44447750E-16*wr*wr*1e12+1.92571880E-15*wr*1e6-3.03397356E-15)*lr*1e6+(8.21218223E-17*wr*wr*1e12-5.44799464E-16*wr*1e6+7.12107807E-16))*nf+((4.92041304E-16*wr*wr*1e12-2.95963348E-15*wr*1e6+2.33018270E-15)*lr*lr*1e12+(3.61458691E-15*wr*wr*1e12-2.21771252E-14*wr*1e6+1.83442198E-14)*lr*1e6+(-5.44547212E-16*wr*wr*1e12+3.33982238E-15*wr*1e6-2.09516516E-15)),1e-18)'
+Cds_rf	= 'max((((2.933e-17*pwr((wr*0.9*1e+6),1.155)-2.83e-18)*pwr((lr*0.9*1e+6),-1)+(4.396e-16*(wr*0.9*1e+6)-7.3e-17))*nf-(7.654e-16*pwr((wr*0.9*1e+6),0.5752)-6.208e-16)), 1e-18)'
+Rds_rf	= 'max((((8805*pwr((wr*0.9*1e+6),-2.69)+3416)*(lr*0.9*1e+6)+(-126.3*pwr((wr*0.9*1e+6),1.417)+1574))*pwr((nf+3),-1)+5),1e-6)'
+Rsub1_rf	= 10
+Rsub2_rf	= 100
+Rsub3_rf	= 100
+Djdb_AREA_rf	= '(int((nf+1)/2)*(wr*0.9*(0.42e-6*0.9-2*6.5e-8)))/0.81'
+Djdb_PJ_rf	= '(int((nf+1)/2)*(2*(0.42e-6*0.9-2*6.5e-8)+2*wr*0.9*4.670E-10/7.53E-11))/0.9'
+Djsb_AREA_rf	= '((int(nf/2)+1)*(wr*0.9*(0.42e-6*0.9-2*6.5e-8)))/0.81'
+Djsb_PJ_rf	= '((int(nf/2)+1)*(2*(0.42e-6*0.9-2*6.5e-8)+2*wr*0.9*4.670E-10/7.53E-11))/0.9'
+Rdc_p12	= 'max((307.9*pwr((wr*0.9*1e+6),-1.333)-4.347),1e-6)'
+Rsc_p12	= 'max((307.9*pwr((wr*0.9*1e+6),-1.333)-4.347),1e-6)'
*****************************************
Lgate       2 20 1p m=mr
Rgate       20 21 'Rg_rf*2' m=mr
Cgd_ext     20 11 'Cgd_rf' m=mr
Cgs_ext     20 31 'max(Cgs_rf+(1e-17+(0.26e-15*nf*(wr*1e+6))*pwr((1+exp((-v(2,3)-0.3)*5)),-1)),1e-18)' m=mr
Rds         11 15 Rds_rf m=mr
Cds_ext     15 31 'max(Cds_rf*(((7.17048693E-04*wr*wr*1e12-5.11775620E-03*wr*1e6+6.49302354E-03)*nf*nf+(-8.91828728E-02*wr*wr*1e12+6.29713310E-01*wr*1e6-8.20559008E-01)*nf+(1.85468115E+00*wr*wr*1e12- 1.26959133E+01*wr*1e6+1.84411904E+01))*lr*lr*1e12+((-3.24470143E-04*wr*wr*1e12+2.55743062E-03*wr*1e6-3.79808399E-03)*nf*nf+(4.30812000E-02*wr*wr*1e12- 3.29474125E-01*wr*1e6+4.80432895E-01)*nf+(-9.74937677E-01*wr*wr*1e12+6.96001900E+00*wr*1e6- 1.14824242E+01))*lr*1e6+((3.72103444E-05*wr*wr*1e12- 3.54043277E-04*wr*1e6+6.28262588E-04)*nf*nf+(-5.05023994E-03*wr*wr*1e12+4.49903867E-02*wr*1e6- 7.32290732E-02)*nf+( 1.10339667E-01*wr*wr*1e12- 8.44616443E-01*wr*1e6+2.01143061E+00))),1e-18)' m=mr
Ldrain       1 11 1p m=mr
Lsource      3 31 1p m=mr
*****************************************
Djdb  11 12
+ pdio12_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
+ m     = mr
***
Djsb  31 32
+ pdio12_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
+ m     = mr
*****************************************
Rsub1      41  4  Rsub1_rf m=mr
Rsub2      41  12 Rsub2_rf m=mr
Rsub3      41  32 Rsub3_rf m=mr
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 p12_rf L=lr W='wr*nf' m=mr AD = 0 AS = 0 PD = 0 PS = 0 sa=sar sb=sbr rdc='Rdc_p12/nf' rsc='Rsc_p12/nf'
* MOS Model
.MODEL  P12_RF  PMOS
+level = 49
**************************************************************
*               MODEL FLAG PARAMETERS 
**************************************************************
+version = 3.24            lmin    = 1.3e-007        lmax    = 2e-005        
+wmin    = 1.5e-007        wmax    = 0.0001          binunit = 2             
+mobmod  = 1               capmod  = 3               nqsmod  = 0             
+stimod  = 1             
**************************************************************
*               GENERAL MODEL PARAMETERS 
**************************************************************
+tnom    = 25              tox     = '2.52e-009+dtox_p12_rf_mismatch'       toxm    = 2.52e-009     
+wint    = 1.2989999e-008  lint    = 0               dlc     = 1.3e-009      
+dwc     = -2.8e-008       hdif    = 1.25e-007       ldif    = 6.5e-008      
+xl      = '1.26e-8+dxl_p12_rf_mismatch'               xw      = '0+dxw_p12_rf'               xj      = 1.6e-007      
+ngate   = 2.6e+020    dlcig   = 3.6e-009      ll      = 3.5e-013        wl      = -2.5270001e-012
+lln     = 0.39            wln     = 0.36            lw      = -3.182e-012   
+ww      = -5.77e-016      lwn     = 0.73            wwn     = 1.1           
+lwl     = 4.5e-015        wwl     = -2.355e-018     llc     = 0             
+wlc     = 0               lwc     = 0               wwc     = 0             
+lwlc    = 0               wwlc    = 0               xpart   = 0             
+igcmod  = 1               igbmod  = 1             
**************************************************************
*               EXPERT PARAMETERS 
**************************************************************
+vth0    = '-0.273+dvth_p12_rf'          lvth0   = -1.3e-008     wvth0   = -7e-009       
+pvth0   = '-7.6e-015+dpvth0_p12_rf'       k1      = 0.37086         wk1     = -5.412e-010   
+pk1     = 3.493e-015      k2      = 0.011828        k3      = -9.37         
+k3b     = 3.4704          nlx     = '1.63e-008+dnlx_p12_rf'       w0      = 6.85e-008     
+dvt0    = 33              ldvt0   = 7.207e-009      dvt1    = 1.65          
+dvt2    = 1.5             ldvt2   = -1.6830001e-007  dvt0w   = 1.2           
+dvt1w   = 1380000         dvt2w   = 0.005831        nch     = 3.5e+017      
+voff    = -0.10809        lvoff   = -3.6e-009       nfactor = 1.2232        
+cdsc    = 0               cdscb   = 0               cdscd   = 0             
+cit     = 0.00036965      lcit    = 4.5e-010        alpha0  = 2.561e-008    
+lalpha0 = 2.655e-016      alpha1  = 0.1669          beta0   = 14.81         
+eta0    = 0.215           etab    = -0.082          dsub    = 0.56          
+pdsub   = -1.4e-014       u0      = '0.0078+du0_p12_rf'          lu0     = '1.095e-010+dlu0_p12_rf'    
+wu0     = '-9.35e-013+dwu0_p12_rf'      pu0     = '3.3e-016+dpu0_p12_rf'        ua      = -4.55e-010    
+wua     = -3.6064e-017    ub      = 1.9e-018        lub     = -1.67e-025    
+pub     = -3.368e-032     uc      = -1.1372e-011    luc     = -2.0000001e-018
+puc     = -4.708e-024     prwg    = 1.3             prwb    = 0.3           
+wr      = 1.0586609       pwr     = 3.401076e-016   rdsw    = 0           
+a0      = 1.58            ags     = 0.36            lags    = 1.556e-007    
+wags    = 5e-008          a1      = 0               a2      = 0.9252        
+pa2     = 1.5e-014        b0      = 6e-008          b1      = 0             
+vsat    = 250000          lvsat   = '-0.021199999+dlvsat_p12_rf'    pvsat   = '-1e-009+dpvsat_p12_rf'       
+keta    = 0.063704        lketa   = 1e-009          wketa   = -6e-009       
+pketa   = -1.5e-015       delta   = 0.018           dwg     = -6.1e-009     
+dwb     = -1.576e-009     pclm    = 0.4512          lpclm   = 1e-007        
+ppclm   = 3.5e-013        pdiblc1 = 0.0001          pdiblc2 = 0.0086        
+pdiblcb = 0               drout   = 0.56            pvag    = 0             
+pscbe1  = 4.2e+008        pscbe2  = 5e-007          elm     = 5             
+agidl   = '9.1278e-012+dagidl_p12_rf'     bgidl   = 86254000        cgidl   = 122           
+egidl   = 0.25            aigbacc = 0.0136          bigbacc = 0.00171          
+cigbacc = 0.075           nigbacc = 1               aigbinv = 0.0111        
+bigbinv = 0.000949        cigbinv = 0.006           eigbinv = 1.1           
+nigbinv = 3               aigc    = 0.007548          bigc    = 0.00075075      
+cigc    = 0.03            nigc    = 3              pigcd   = 2             
+aigsd   = 0.0062          bigsd   = 0.0003          cigsd   = 0.04          
+poxedge = 1               ntox    = 1             
**************************************************************
*               CAPACITANCE PARAMETERS 
**************************************************************
+acde    = 0.49772         moin    = 10              noff    = 1.65          
+voffcv  = 0.00043808      cgbo    = 0               cgso    = 0      
+cgdo    = 0        cf      = 0             
+clc     = 1e-18 
**************************************************************
*               TEMPERATURE PARAMETERS 
**************************************************************
+kt1     = -0.2519         kt1l    = -3.792e-009     kt2     = 0             
+pkt2    = -2.3e-015       ute     = -1.18           lute    = 5.2e-008      
+wute    = -2e-008         pute    = 2.2e-014        ua1     = 8e-010        
+lua1    = 3.388e-018      wua1    = 4.1e-017        ub1     = -1.5e-018     
+lub1    = 1.2e-025        wub1    = -5e-026         pub1    = -5e-033       
+uc1     = -5e-011         prt     = 0               at      = 33000         
+pat     = 1e-009        
**************************************************************
*               NOISE PARAMETERS 
**************************************************************
+noia    = 6.7163E+18      noib    = 6.8409E+06      noic    = -1.6028E-11  
+em      = 7.4377E+07      ef      = 1.16005         noimod  = 2               
**************************************************************
*               DIODE PARAMETERS 
**************************************************************
+rsh     = 6.98            js      = 2.3e-007        jsw     = 5e-012        
+cj      = 0         mj      = 0.431           cjsw    = 0    
+mjsw    = 0.346           cjswg   = 0         mjswg   = 0.499         
+pb      = 0.785           pbsw    = 0.472           pbswg   = 0.93          
+rd      = 0               rdc     = 'Rdc_p12/nf'             rs      = 0             
+rsc     = 'Rsc_p12/nf'             xti     = 3               tpb     = 0.0012231       
+tpbsw   = 0.00036         tpbswg  = 0.00277         tcj     = 0.000872      
+tcjsw   = 0.000755        tcjswg  = 0.000787        acm     = 12            
+calcacm = 1               nj      = 1.0188        
**************************************************************
*               STRESS PARAMETERS 
**************************************************************
+saref   = 2.25e-006       sbref   = 2.25e-006       wlod    = 0             
+kvth0   = 1.5e-008        lkvth0  = 1e-005          wkvth0  = 1e-006        
+pkvth0  = 0               llodvth = 1               wlodvth = 1             
+stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 2e-007          lku0    = 4e-007          wku0    = 5e-007        
+pku0    = 0               llodku0 = 1               wlodku0 = 1             
+kvsat   = -1              steta0  = 0               tku0    = 0             
*
***********************************************************************************
*                            1.2V P+/NWELL DIODE MODEL                            *
***********************************************************************************
*
.MODEL PDIO12_RF D
+LEVEL    = 3                   JS       = 2.30E-07  JSW      = 1.31E-13
+N        = 1.0188  RS       = 1.0E-010              IK       = 1.0E+21 
+IKR      = 2.78E+05            BV       = 10.1                  IBV      = 277.8
+TRS      = 1.09E-03            EG       = 1.16                  TREF     = 25.0
+XTI      = 3.0                 TLEV     = 1                     TLEVC    = 1
+CJ       = '1.22E-03+DCJ_P12_RF'
+CJSW     = '7.53E-11+DCJSW_P12_RF'
+MJ       = 0.431               PB       = 0.785
+MJSW     = 0.346               PHP      = 0.472
+CTA      = 8.72E-04            CTP      = 7.55E-04              TPB      = 0.0012231
+TPHP     = 3.60E-04            FC       = 0                     FCS      = 0
+AREA     = 3.60E-09            PJ       = 2.4E-04
.ends p12_ckt_rf
*
*************************
* 3.3V RF NMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt n33_ckt_rf 1 2 3 4 lr=l wr=w nf=finger sar=sa sbr=sb mr=m mismod=0 
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+atox_n33_rf = 4e-11
+axl_n33_rf = 3e-9
+avth_n33_rf = 9.5e-3
+au0_n33_rf = 6e-4
+lef = lr
+wef = 'wr*nf'
+dtox_n33_mis_rf = 'atox_n33_rf*1/sqrt(lef*wef*1e12*mr)*sigma_mis_a_rf*mismod'
+dxl_n33_mis_rf = 'axl_n33_rf*1/sqrt(wef*1e6*mr)*sigma_mis_b_rf*mismod'
+dvth_n33_mis_rf = 'avth_n33_rf*1/sqrt(lef*wef*1e12*mr)*sigma_mis_c_rf*mismod'
+du0_n33_mis_rf = 'au0_n33_rf*1/sqrt(lef*wef*1e12*mr)*sigma_mis_d_rf*mismod'
+Rg_rf        = 'max(((-24.56*pwr((wr*1e+6),2)+874.3)*pwr((10*lr*1e+6),-1)+(733.3*pwr((wr*1e+6),-1)+27.34))*pwr((nf+3),-1)+1, 1e-6)'
+Cgd_rf       = 'max((((2.899e-15*pwr((wr*1e+6),0.4868)-1.844e-15)*pwr((10*lr*1e+6),0.1)+(-4.973e-15*pwr((wr*1e+6),0.2754)+4.324e-15))*nf)*0.9, 1e-18)'
+Cgs_rf       = 'max((((5.533e-18*pwr((wr*1e+6),-1)-7.483e-18)*pwr((10*lr*1e+6),2)+(-0.8197e-15*pwr((wr*1e+6),-0.1142)+1.356e-15))*pwr(nf,0.9))*1.2,1e-18)'
+Rsub2_rf     = 'max((((78.26e+3*pwr((wr*1e+6),-0.220)-49.51e+3)*pwr((10*lr*1e+6),-1)+(-1.119e+3*(wr*1e+6)+7.89e+3))*pwr((nf+3),-1))*0.4,1)'
+Rsub3_rf     = 'max((((78.26e+3*pwr((wr*1e+6),-0.220)-49.51e+3)*pwr((10*lr*1e+6),-1)+(-1.119e+3*(wr*1e+6)+7.89e+3))*pwr((nf+3),-1))*0.4,1)'
+Djdb_AREA_rf = 'int(0.5*(nf+1))*(wr*(0.46e-6-2*0.0825e-6))'
+Djdb_PJ_rf   = 'int(0.5*(nf+1))*(2*(0.46e-6-2*0.0825e-6)+2*wr*2.2322)'
+Djsb_AREA_rf = 'int(0.5*nf+1)*(wr*(0.46e-6-2*0.0825e-6))'
+Djsb_PJ_rf   = 'int(0.5*nf+1)*(2*(0.46e-6-2*0.0825e-6)+2*wr*2.2322)'
*****************************************
Lgate       2 20 1p m=mr
Rgate       20 21 Rg_rf m=mr
Cgd_ext     20 11 Cgd_rf m=mr
Cgs_ext     20 31 Cgs_rf m=mr
Cds_ext     15 31 1e-18 m=mr
Rds         11 15 220 m=mr
Ldrain       1 11 1p m=mr
Lsource      3 31 1p m=mr
*****************************************
Djdb  12 11 
+ ndio33_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
+ m     = mr
***
Djsb  32 31 
+ ndio33_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
+ m      = mr
*****************************************
Rsub1      41  4  0.75 m=mr
Rsub2      41  12 Rsub2_rf m=mr
Rsub3      41  32 Rsub3_rf m=mr
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 n33_rf L=lr W='wr*nf' m=mr AD = 0 AS = 0 PD = 0 PS = 0 sa=sar sb=sbr 
* MOS Model
.model  n33_rf  nmos
+level = 49
**************************************************************
*               MODEL FLAG PARAMETERS 
**************************************************************
+version = 3.24            lmin    = 3.5e-007        lmax    = 2e-005        
+wmin    = 1.5e-007        wmax    = 0.0001          binunit = 2             
+mobmod  = 1               capmod  = 3               nqsmod  = 0             
+stimod  = 1             
**************************************************************
*               GENERAL MODEL PARAMETERS 
**************************************************************
+tnom    = 25              tox     = '6.9e-009+dtox_n33_rf+dtox_n33_mis_rf'        toxm    = 6.9e-009      
+wint    = 3.8e-008        lint    = 4.2e-008        dlc     = 2e-008        
+dwc     = -2.8e-008       hdif    = 1.275e-007      ldif    = 8.25e-008     
+xl      = '2.88e-008+dxl_n33_rf+dxl_n33_mis_rf'               xw      = '0+dxw_n33_rf'               xj      = 1.75e-007     
+ngate   = 2.8e+020        dlcig   = 4.2e-008        ll      = 0             
+wl      = 0               lln     = 1               wln     = 1             
+lw      = 0               ww      = -5.36e-015      lwn     = 1             
+wwn     = 1.016           lwl     = 0               wwl     = 0             
+llc     = 0               wlc     = 0               lwc     = 0             
+wwc     = 0               lwlc    = 0               wwlc    = 0             
+xpart   = 0             
**************************************************************
*               EXPERT PARAMETERS 
**************************************************************
+vth0    = '0.597+dvth_n33_rf'           lvth0   = '-2.115e-008+dlvth0_n33_rf'      wvth0   = '-1.68e-008+dwvth0_n33_rf'    
+pvth0   = '-5e-015+dpvth0_n33_rf'         k1      = 0.78            k2      = -0.04         
+lk2     = -4e-008         wk2     = -2e-008         pk2     = 2.2e-015      
+k3      = 10              k3b     = 0               nlx     = 1.74e-007     
+w0      = 1.992e-006      pw0     = 1e-019          dvt0    = 1.95          
+pdvt0   = 4e-014          dvt1    = 0.8             pdvt1   = 4.4e-014      
+dvt2    = -0.032          dvt0w   = 0               dvt1w   = 5300000       
+dvt2w   = -0.032          nch     = 4e+016          voff    = -0.14         
+nfactor = 1               cdsc    = 0               cdscb   = 0             
+cdscd   = 0               cit     = 0.001           lcit    = -1.2e-010     
+pcit    = -1.8e-017       alpha0  = 2.6499001e-007  alpha1  = 5.45624       
+beta0   = 22.700001       eta0    = 0.05            etab    = -0.015        
+dsub    = 0.56            u0      = '0.0356+du0_n33_rf'          wu0     = '-1.28e-009+dwu0_n33_rf'   
+lu0     = '0+dlu0_n33_rf'    pu0     = '0+dpu0_n33_rf'  
+ua      = -2.4e-010       ub      = 1.35e-018       lub     = -1.32e-025    
+wub     = -1e-026         pub     = -2.8e-032       uc      = 5.611685e-011 
+luc     = -2.85e-017      prwg    = 0               prwb    = 0.001         
+wr      = 1               rdsw    = 500             a0      = 0.765         
+la0     = 1.4e-008        pa0     = -5e-014         ags     = 0.233         
+lags    = 1.1e-007        pags    = 9e-014          a1      = 0             
+a2      = 1               b0      = 1e-008          b1      = 0             
+vsat    = 77080           lvsat   = '-0.0005+dlvsat_n33_rf'         pvsat   = 6e-010        
+keta    = -0.04           lketa   = 5e-009          pketa   = 3e-015        
+delta   = 0.01            dwg     = 0               dwb     = 0             
+pclm    = 1.2             pdiblc1 = 0.05616         pdiblc2 = 0.0008        
+pdiblcb = 0               drout   = 0.56            pvag    = 0             
+pscbe1  = 4.24e+008       pscbe2  = 1e-005          elm     = 5             
+agidl   = '4.5e-011+dagidl_n33_rf'        bgidl   = 1.5062e+009     cgidl   = 100           
+egidl   = 1             
**************************************************************
*               CAPACITANCE PARAMETERS 
**************************************************************
+clc     = 1e-18             cle     = 0.6             acde    = 0.4           
+moin    = 5               noff    = 2.5             voffcv  = -0.03         
+lvoffcv = -3e-008         cgbo    = 0               cgso    = '1e-18'        
+cgdo    = '1e-18'          cgdl    = 1.0e-018        cgsl    = 1.0e-18      
+cf      = 1e-18        
**************************************************************
*               TEMPERATURE PARAMETERS 
**************************************************************
+kt1     = -0.337001       lkt1    = 1e-009          wkt1    = 2e-009        
+pkt1    = 3e-015          kt1l    = 5.192e-009      kt2     = -0.03845153   
+lkt2    = -7.5e-009       pkt2    = 6e-016          ute     = -1.6497999    
+lute    = 1.5e-007        wute    = 8e-008          pute    = 1e-014        
+ua1     = 1.5619001e-009  lua1    = 5e-016          pua1    = -1e-023       
+ub1     = -2.1351e-018    uc1     = -1.84e-011      prt     = 0             
+at      = 30000           lat     = -0.005          pat     = 1e-010        
**************************************************************
*               NOISE PARAMETERS 
**************************************************************
+noia    = 2.4433E+20       noib    = 3.1826E+04      noic    = -4.1964E-13    
+em      = 8.0759E+07       ef      = 0.8202          noimod  = 2             
**************************************************************
*               DIODE PARAMETERS 
**************************************************************
+rsh     = 6.45            js      = 1.5e-007        jsw     = 5e-012        
+cj      = '1e-18'          mj      = 0.267           cjsw    = '1e-18'     
+mjsw    = 0.193           cjswg   = '1e-18'       mjswg   = 0.359         
+pb      = 0.653           pbsw    = 0.996           pbswg   = 0.86          
+rd      = 0               rdc     = 1.5             rs      = 0             
+rsc     = 1.5             xti     = 3               tpb     = 0.00198       
+tpbsw   = 0.00142         tpbswg  = 0.00188         tcj     = 0.00095       
+tcjsw   = 0.000617        tcjswg  = 0.000934        acm     = 12            
+calcacm = 1               nj      = 1.012         
**************************************************************
*               STRESS PARAMETERS 
**************************************************************
+saref   = 3.32e-006       sbref   = 3.32e-006       wlod    = 0             
+kvth0   = 2e-008          lkvth0  = 2.5e-007        wkvth0  = 0             
+pkvth0  = 0               llodvth = 1               wlodvth = 1             
+stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = -1.015e-007     lku0    = 1.5e-007        wku0    = 1e-007        
+pku0    = 0               llodku0 = 1               wlodku0 = 1             
+kvsat   = 0.45            steta0  = 0               tku0    = 0             
*
*
.model ndio33_rf d
+LEVEL    = 3                       JS       = 1.50E-07 JSW      = 1.00E-15             
+N        = 1.012       RS       = 1.0E-010              IK       = 1.0E+21                   
+IKR      = 2.78E+05                BV       = 11.36                 IBV      = 277.8            
+TRS      = 1.11E-03                EG       = 1.16                  TREF     = 25.0                
+XTI      = 3.0                     TLEV     = 1                     TLEVC    = 1
+CJ       = '9.00E-04+DCJ_N33_rf'   MJ       = 0.267                 PB       = 0.653               
+CJSW     = '1.016E-10+DCJSW_N33_rf' MJSW     = 0.193                 PHP      = 0.996               
+TPB      = 1.7E-03                TPHP     = 1.42E-03              FCS      = 0
+CTA      = 9.50E-04                CTP      = 6.17E-04              FC       = 0
+AREA     = 3.60E-09                PJ       = 2.4E-04  
*
.ends n33_ckt_rf
*************************
* 3.3V RF DNWMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt dnw33_ckt_rf 1 2 3 4 lr=l wr=w nf=finger sar=sa sbr=sb mr=m mismod=0 
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+atox_n33_rf = 4e-11
+axl_n33_rf = 3e-9
+avth_n33_rf = 9.5e-3
+au0_n33_rf = 6e-4
+lef = lr
+wef = 'wr*nf'
+dtox_n33_mis_rf = 'atox_n33_rf*1/sqrt(lef*wef*1e12*mr)*sigma_mis_a_rf*mismod'
+dxl_n33_mis_rf = 'axl_n33_rf*1/sqrt(wef*1e6*mr)*sigma_mis_b_rf*mismod'
+dvth_n33_mis_rf = 'avth_n33_rf*1/sqrt(lef*wef*1e12*mr)*sigma_mis_c_rf*mismod'
+du0_n33_mis_rf = 'au0_n33_rf*1/sqrt(lef*wef*1e12*mr)*sigma_mis_d_rf*mismod'
+Rg_rf        = 'max(((-24.56*pwr((wr*1e+6),2)+874.3)*pwr((10*lr*1e+6),-1)+(733.3*pwr((wr*1e+6),-1)+27.34))*pwr((nf+3),-1)+1, 1e-6)'
+Cgd_rf       = 'max((((2.899e-15*pwr((wr*1e+6),0.4868)-1.844e-15)*pwr((10*lr*1e+6),0.1)+(-4.973e-15*pwr((wr*1e+6),0.2754)+4.324e-15))*nf)*0.9, 1e-18)'
+Cgs_rf       = 'max((((5.533e-18*pwr((wr*1e+6),-1)-7.483e-18)*pwr((10*lr*1e+6),2)+(-0.8197e-15*pwr((wr*1e+6),-0.1142)+1.356e-15))*pwr(nf,0.9))*1.2,1e-18)'
+Rsub2_rf     = 'max((((78.26e+3*pwr((wr*1e+6),-0.220)-49.51e+3)*pwr((10*lr*1e+6),-1)+(-1.119e+3*(wr*1e+6)+7.89e+3))*pwr((nf+3),-1))*0.4,1)'
+Rsub3_rf     = 'max((((78.26e+3*pwr((wr*1e+6),-0.220)-49.51e+3)*pwr((10*lr*1e+6),-1)+(-1.119e+3*(wr*1e+6)+7.89e+3))*pwr((nf+3),-1))*0.4,1)'
+Djdb_AREA_rf = 'int(0.5*(nf+1))*(wr*(0.46e-6-2*0.0825e-6))'
+Djdb_PJ_rf   = 'int(0.5*(nf+1))*(2*(0.46e-6-2*0.0825e-6)+2*wr*2.2322)'
+Djsb_AREA_rf = 'int(0.5*nf+1)*(wr*(0.46e-6-2*0.0825e-6))'
+Djsb_PJ_rf   = 'int(0.5*nf+1)*(2*(0.46e-6-2*0.0825e-6)+2*wr*2.2322)'
*****************************************
Lgate       2 20 1p m=mr
Rgate       20 21 Rg_rf m=mr
Cgd_ext     20 11 Cgd_rf m=mr
Cgs_ext     20 31 Cgs_rf m=mr
Cds_ext     15 31 1e-18 m=mr
Rds         11 15 220 m=mr
Ldrain       1 11 1p m=mr
Lsource      3 31 1p m=mr
*****************************************
Djdb  12 11 
+ ndio33_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
+ m     = mr
***
Djsb  32 31 
+ ndio33_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
+ m      = mr
*****************************************
Rsub1      41  4  0.75 m=mr
Rsub2      41  12 Rsub2_rf m=mr
Rsub3      41  32 Rsub3_rf m=mr
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 dnw33_rf L=lr W='wr*nf' m=mr AD = 0 AS = 0 PD = 0 PS = 0 sa=sar sb=sbr 
* MOS Model
.model  dnw33_rf  nmos
+level = 49
**************************************************************
*               MODEL FLAG PARAMETERS 
**************************************************************
+version = 3.24            lmin    = 3.5e-007        lmax    = 2e-005        
+wmin    = 1.5e-007        wmax    = 0.0001          binunit = 2             
+mobmod  = 1               capmod  = 3               nqsmod  = 0             
+stimod  = 1             
**************************************************************
*               GENERAL MODEL PARAMETERS 
**************************************************************
+tnom    = 25              tox     = '6.9e-009+dtox_n33_rf+dtox_n33_mis_rf'        toxm    = 6.9e-009      
+wint    = 3.8e-008        lint    = 4.2e-008        dlc     = 2e-008        
+dwc     = -2.8e-008       hdif    = 1.275e-007      ldif    = 8.25e-008     
+xl      = '2.88e-008+dxl_n33_rf+dxl_n33_mis_rf'               xw      = '0+dxw_n33_rf'               xj      = 1.75e-007     
+ngate   = 2.8e+020        dlcig   = 4.2e-008        ll      = 0             
+wl      = 0               lln     = 1               wln     = 1             
+lw      = 0               ww      = -5.36e-015      lwn     = 1             
+wwn     = 1.016           lwl     = 0               wwl     = 0             
+llc     = 0               wlc     = 0               lwc     = 0             
+wwc     = 0               lwlc    = 0               wwlc    = 0             
+xpart   = 0             
**************************************************************
*               EXPERT PARAMETERS 
**************************************************************
+vth0    = '0.597+dvth_n33_rf'           lvth0   = '-2.115e-008+dlvth0_n33_rf'      wvth0   = '-1.68e-008+dwvth0_n33_rf'    
+pvth0   = '-5e-015+dpvth0_n33_rf'         k1      = 0.78            k2      = -0.04         
+lk2     = -4e-008         wk2     = -2e-008         pk2     = 2.2e-015      
+k3      = 10              k3b     = 0               nlx     = 1.74e-007     
+w0      = 1.992e-006      pw0     = 1e-019          dvt0    = 1.95          
+pdvt0   = 4e-014          dvt1    = 0.8             pdvt1   = 4.4e-014      
+dvt2    = -0.032          dvt0w   = 0               dvt1w   = 5300000       
+dvt2w   = -0.032          nch     = 4e+016          voff    = -0.14         
+nfactor = 1               cdsc    = 0               cdscb   = 0             
+cdscd   = 0               cit     = 0.001           lcit    = -1.2e-010     
+pcit    = -1.8e-017       alpha0  = 2.6499001e-007  alpha1  = 5.45624       
+beta0   = 22.700001       eta0    = 0.05            etab    = -0.015        
+dsub    = 0.56            u0      = '0.0356+du0_n33_rf'          wu0     = '-1.28e-009+dwu0_n33_rf'   
+lu0     = '0+dlu0_n33_rf'    pu0     = '0+dpu0_n33_rf'  
+ua      = -2.4e-010       ub      = 1.35e-018       lub     = -1.32e-025    
+wub     = -1e-026         pub     = -2.8e-032       uc      = 5.611685e-011 
+luc     = -2.85e-017      prwg    = 0               prwb    = 0.001         
+wr      = 1               rdsw    = 500             a0      = 0.765         
+la0     = 1.4e-008        pa0     = -5e-014         ags     = 0.233         
+lags    = 1.1e-007        pags    = 9e-014          a1      = 0             
+a2      = 1               b0      = 1e-008          b1      = 0             
+vsat    = 77080           lvsat   = '-0.0005+dlvsat_n33_rf'         pvsat   = 6e-010        
+keta    = -0.04           lketa   = 5e-009          pketa   = 3e-015        
+delta   = 0.01            dwg     = 0               dwb     = 0             
+pclm    = 1.2             pdiblc1 = 0.05616         pdiblc2 = 0.0008        
+pdiblcb = 0               drout   = 0.56            pvag    = 0             
+pscbe1  = 4.24e+008       pscbe2  = 1e-005          elm     = 5             
+agidl   = '4.5e-011+dagidl_n33_rf'        bgidl   = 1.5062e+009     cgidl   = 100           
+egidl   = 1             
**************************************************************
*               CAPACITANCE PARAMETERS 
**************************************************************
+clc     = 1e-18             cle     = 0.6             acde    = 0.4           
+moin    = 5               noff    = 2.5             voffcv  = -0.03         
+lvoffcv = -3e-008         cgbo    = 0               cgso    = '1e-18'        
+cgdo    = '1e-18'          cgdl    = 1.0e-018        cgsl    = 1.0e-18      
+cf      = 1e-18        
**************************************************************
*               TEMPERATURE PARAMETERS 
**************************************************************
+kt1     = -0.337001       lkt1    = 1e-009          wkt1    = 2e-009        
+pkt1    = 3e-015          kt1l    = 5.192e-009      kt2     = -0.03845153   
+lkt2    = -7.5e-009       pkt2    = 6e-016          ute     = -1.6497999    
+lute    = 1.5e-007        wute    = 8e-008          pute    = 1e-014        
+ua1     = 1.5619001e-009  lua1    = 5e-016          pua1    = -1e-023       
+ub1     = -2.1351e-018    uc1     = -1.84e-011      prt     = 0             
+at      = 30000           lat     = -0.005          pat     = 1e-010        
**************************************************************
*               NOISE PARAMETERS 
**************************************************************
+noia    = 2.4433E+20       noib    = 3.1826E+04      noic    = -4.1964E-13    
+em      = 8.0759E+07       ef      = 0.8202          noimod  = 2             
**************************************************************
*               DIODE PARAMETERS 
**************************************************************
+rsh     = 6.45            js      = 1.5e-007        jsw     = 5e-012        
+cj      = '1e-18'          mj      = 0.267           cjsw    = '1e-18'     
+mjsw    = 0.193           cjswg   = '1e-18'       mjswg   = 0.359         
+pb      = 0.653           pbsw    = 0.996           pbswg   = 0.86          
+rd      = 0               rdc     = 1.5             rs      = 0             
+rsc     = 1.5             xti     = 3               tpb     = 0.00198       
+tpbsw   = 0.00142         tpbswg  = 0.00188         tcj     = 0.00095       
+tcjsw   = 0.000617        tcjswg  = 0.000934        acm     = 12            
+calcacm = 1               nj      = 1.012         
**************************************************************
*               STRESS PARAMETERS 
**************************************************************
+saref   = 3.32e-006       sbref   = 3.32e-006       wlod    = 0             
+kvth0   = 2e-008          lkvth0  = 2.5e-007        wkvth0  = 0             
+pkvth0  = 0               llodvth = 1               wlodvth = 1             
+stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = -1.015e-007     lku0    = 1.5e-007        wku0    = 1e-007        
+pku0    = 0               llodku0 = 1               wlodku0 = 1             
+kvsat   = 0.45            steta0  = 0               tku0    = 0             
*
.model ndio33_rf d
+LEVEL    = 3                       JS       = 1.50E-07 JSW      = 1.00E-15             
+N        = 1.012       RS       = 1.0E-010              IK       = 1.0E+21                   
+IKR      = 2.78E+05                BV       = 11.36                 IBV      = 277.8            
+TRS      = 1.11E-03                EG       = 1.16                  TREF     = 25.0                
+XTI      = 3.0                     TLEV     = 1                     TLEVC    = 1
+CJ       = '9.00E-04+DCJ_N33_rf'   MJ       = 0.267                 PB       = 0.653               
+CJSW     = '1.016E-10+DCJSW_N33_rf' MJSW     = 0.193                 PHP      = 0.996               
+TPB      = 1.7E-03                TPHP     = 1.42E-03              FCS      = 0
+CTA      = 9.50E-04                CTP      = 6.17E-04              FC       = 0
+AREA     = 3.60E-09                PJ       = 2.4E-04  
*
.ends dnw33_ckt_rf
*************************
* 3.3V RF PMOS Subcircuit
*************************
* 11=drain, 2=gate, 31=source, 4=bulk
* lr=gate length, wr=finger width, nf=finger number
.subckt p33_ckt_rf 1 2 3 4 lr=l wr=w nf=finger sar=sa sbr=sb mr=1 mismod=0 
* scalable unit parameter
* euqivalent circuit saclable parameter
.param
+atox_p33_rf=3e-11
+axl_p33_rf=3e-10
+avth_p33_rf=3.5e-3
+au0_p33_rf=1e-4
+lef=lr
+wef=wr
+dtox_p33_rf_mis='atox_p33_rf*1/sqrt(lef*wef*1e12*mr*nf)*sigma_mis_a_rf*mismod'
+dxl_p33_rf_mis='axl_p33_rf*1/sqrt(wef*1e6*mr*nf)*sigma_mis_b_rf*mismod'
+dvth_p33_rf_mis='avth_p33_rf*1/sqrt(lef*wef*1e12*mr*nf)*sigma_mis_c_rf*mismod'
+du0_p33_rf_mis='au0_p33_rf*1/sqrt(lef*wef*1e12*mr*nf)*sigma_mis_d_rf*mismod'
+dtox_p33_rf_mismatch         = 'dtox_p33_rf+dtox_p33_rf_mis' 
+dxl_p33_rf_mismatch         = 'dxl_p33_rf+dxl_p33_rf_mis' 
+dvth_p33_rf_mismatch         = 'dvth_p33_rf+dvth_p33_rf_mis' 
+du0_p33_rf_mismatch         = 'du0_p33_rf_mis' 
*define lsh as shrunk length, wsh as shrunk width, and the unit is um
+lsh  = 'lr*1e+6*0.9+0.0288'        wsh    = 'wr*1e+6*0.9'
+Rg_rf        = 'max(((-9.3001*pwr(lsh,2)+14.937*lsh-4.1198)*pwr(wsh,2)+(67.514*pwr(lsh,2)-104.17*lsh+26.521)*wsh+(-84.985*pwr(lsh,2)+123.63*lsh-20.093))+((466.56*pwr(lsh,2)-816.42*lsh+373.94)*pwr(wsh,2)+(-3480.1*pwr(lsh,2)+5874.3*lsh-2760.5)*wsh+(7052.4*pwr(lsh,2)-10449*lsh+5055.5))/nf, 1e-6)'
+Rds_rf       = 'max(((-3.644*pwr(lsh,2)+4.7372*lsh-1.0932)*pwr(wsh,2)+(23.413*pwr(lsh,2)-26.213*lsh+5.2978)*wsh+(-34.588*pwr(lsh,2)+34.762*lsh-6.2572))*nf+((220*pwr(lsh,2)-286*lsh+66)*pwr(wsh,2)+(-1217.2*pwr(lsh,2)+1502.6*lsh-315.92)*wsh+(1439*pwr(lsh,2)-1678.9*lsh+367.41)), 1e-3)'
+Cgd_rf       = 'max(((1.85820000E-19*wr*wr*1e12+3.96236300E-17*wr*1e6-1.12700745E-15)*lr*lr*lr*1e18+(6.91922667E-18*wr*wr*1e12-1.49251960E-16*wr*1e6+1.55616373E-15)*lr*lr*1e12+(-1.43913933E-17*wr*wr*1e12+2.25474910E-16*wr*1e6-4.42827917E-16)*lr*1e6+(5.02854000E-18*wr*wr*1e12+2.09109910E-16*wr*1e6+2.85209950E-16))*nf+((-2.33573863E-16*wr*wr*1e12+3.63961563E-15*wr*1e6-2.76600356E-15)*lr*lr*lr*1e18+(2.89285395E-16*wr*wr*1e12-6.70547717E-15*wr*1e6+5.97036097E-15)*lr*lr*1e12+(-1.60514807E-17*wr*wr*1e12+3.43888741E-15*wr*1e6-3.81974003E-15)*lr*1e6+(-4.05390861E-17*wr*wr*1e12-3.75779826E-16*wr*1e6+4.46127282E-16)),1e-18)'
+Cgs_rf       = 'max(((4.70325107E-17*wr*wr*1e12-2.16946909E-16*wr*1e6+3.64865980E-16)*lr*lr*1e12+(-9.34999398E-17*wr*wr*1e12+2.42129081E-16*wr*1e6-6.87636912E-16)*lr*1e6+(3.85222690E-17*wr*wr*1e12+1.60751395E-18*wr*1e6+5.44514706E-16))*nf+((-9.44616018E-16*wr*wr*1e12+5.53137711E-15*wr*1e6-9.86636049E-15)*lr*lr*1e12+(1.40434764E-15*wr*wr*1e12-8.75908051E-15*wr*1e6+1.42587707E-14)*lr*1e6+(-3.71698937E-16*wr*wr*1e12+2.73125740E-15*wr*1e6-3.75676788E-15)),1e-18)'
+Cds_rf       = 'max(((-4.61639493E-16*wr*wr*1e12+1.42197020E-15*wr*1e6+3.83562333E-16)*lr*lr*1e12+(5.99650987E-16*wr*wr*1e12-2.12031960E-15*wr*1e6-5.13246667E-16)*lr*1e6+(-1.31118272E-16*wr*wr*1e12+6.35147746E-16*wr*1e6+1.05148738E-16))*nf+((6.76813867E-15*wr*wr*1e12-9.59323200E-15*wr*1e6-3.15398867E-14)*lr*lr*1e12+(-8.98097700E-15*wr*wr*1e12+1.37834595E-14*wr*1e6+4.60339275E-14)*lr*1e6+(2.19337400E-15*wr*wr*1e12-4.17706900E-15*wr*1e6-1.45621050E-14)),1e-18)'
+Rsub1_rf     = 0.75
+Rsub2_rf     = 100
+Rsub3_rf     = 100
+Djdb_AREA_rf = '(int((nf+1)/2)*(wr*0.9*(4.14e-7-2*8.25e-8)))/0.81'
+Djdb_PJ_rf   = '(int((nf+1)/2)*(2*(4.14e-7-2*8.25e-8)+2*wr*0.9*4.700E-10*0.8/4.56E-11))/0.9'
+Djsb_AREA_rf = '((int(nf/2)+1)*(wr*0.9*(4.14e-7-2*8.25e-8)))/0.81'
+Djsb_PJ_rf   = '((int(nf/2)+1)*(2*(4.14e-7-2*8.25e-8)+2*wr*0.9*4.700E-10*0.8/4.56E-11))/0.9'
+Rdc_p33      = 'max(18.7215/(wr*1e6*0.9)+0.0964*nf, 1e-6)'
+Rsc_p33      = 'max(18.7215/(wr*1e6*0.9)+0.0964*nf, 1e-6)'
*****************************************
Lgate       2 20 1p m=mr
Rgate       20 21 Rg_rf m=mr
Cgd_ext     20 11 Cgd_rf m=mr
Cgs_ext     20 31 Cgs_rf m=mr
Cds_ext     15 31 'Cds_rf*0.8' m=mr
Rds         11 15 Rds_rf m=mr
Ldrain       1 11 1p m=mr
Lsource      3 31 1p m=mr
*****************************************
Djdb  11 12
+ pdio33_rf
+ AREA  = Djdb_AREA_rf
+ PJ    = Djdb_PJ_rf 
+ m     = mr
***
Djsb  31 32
+ pdio33_rf
+ AREA  = Djsb_AREA_rf
+ PJ    = Djsb_PJ_rf
+ m     = mr
*****************************************
Rsub1      41  4  Rsub1_rf m=mr
Rsub2      41  12 Rsub2_rf m=mr
Rsub3      41  32 Rsub3_rf m=mr
*
* --------- ideal mos transistor ----------------------
MAIN 11 21 31 41 p33_rf L=lr W='wr*nf' m=mr AD = 0 AS = 0 PD = 0 PS = 0 sa=sar sb=sbr rdc='Rdc_p33/nf' rsc='Rsc_p33/nf' 
* MOS Model
.model p33_rf PMOS
+level = 49
**************************************************************
*               MODEL FLAG PARAMETERS 
**************************************************************
+version = 3.24            lmin    = 3e-007          lmax    = 2e-005        
+wmin    = 1.5e-007        wmax    = 0.0001          binunit = 2             
+mobmod  = 1               capmod  = 3               nqsmod  = 0             
+stimod  = 1             
**************************************************************
*               GENERAL MODEL PARAMETERS 
**************************************************************
+tnom    = 25              tox     = '6.9e-009+dtox_p33_rf_mismatch'        toxm    = 6.9e-009      
+wint    = -1.9e-008       lint    = 2.2e-008        dlc     = 3.6e-008      
+dwc     = -2.8e-008       hdif    = 1.275e-007      ldif    = 8.25e-008     
+xl      = '2.88e-8+dxl_p33_rf_mismatch'               xw      = '0+dxw_p33_rf'               xj      = 2e-007        
+ngate   = 2e+020          dlcig   = 2.1838e-008     ll      = 0             
+wl      = 0               lln     = 1               wln     = 0.972         
+lw      = 0               ww      = -4.6e-015       lwn     = 1             
+wwn     = 1.02            lwl     = 0               wwl     = 0             
+llc     = 0               wlc     = 0               lwc     = 0             
+wwc     = 0               lwlc    = 0               wwlc    = 0             
+xpart   = 0             
**************************************************************
*               EXPERT PARAMETERS 
**************************************************************
+vth0    = '-0.64554+dvth_p33_rf'        lvth0   = '6.53e-008+dlvth0_p33_rf'       wvth0   = '1.8e-008+dwvth0_p33_rf'      
+pvth0   = '-1.2e-016+dpvth0_p33_rf'       k1      = 0.92            k2      = -0.0001       
+lk2     = -1.1e-008       wk2     = -1e-008         pk2     = -2e-015       
+k3      = -4.8            k3b     = 0               nlx     = 1.74e-007     
+w0      = 2e-006          dvt0    = 1.23            dvt1    = 0.8           
+dvt2    = -0.05           dvt0w   = 0               dvt1w   = 5300000       
+dvt2w   = -0.032          nch     = 6e+016          voff    = -0.15         
+nfactor = 1               cdsc    = 0.00024         cdscb   = 0             
+cdscd   = 0               cit     = 0.0007          alpha0  = 4.19e-007     
+alpha1  = 6.746904        beta0   = 29.209999       eta0    = 0.01          
+etab    = -0.012          dsub    = 0.56            u0      = '0.0107+du0_p33_rf'        
+lu0     = '4e-010+dlu0_p33_rf'           wu0     = '-1.44e-009+dwu0_p33_rf'       pu0     = '-5e-017+dpu0_p33_rf'        
+ua      = 6.147218e-010   ub      = 1.2e-018        lub     = 4.4e-026      
+wub     = -4e-025         pub     = 8e-032          uc      = -4.30592e-011 
+wuc     = -1e-017         puc     = 3e-024          prwg    = 0             
+prwb    = 0               wr      = 1               rdsw    = 820           
+a0      = 1.1             ags     = 0.17            a1      = 0             
+a2      = 0.99            b0      = 0               b1      = 0             
+vsat    = 77000           lvsat   = '0.0072+dlvsat_p33_rf'            pvsat   = '-1.2e-009+dpvsat_p33_rf'                 
+keta    = 0               delta   = 0.01            ldelta  = 8.4e-009      
+pdelta  = 2e-015          dwg     = 0               dwb     = 0             
+pclm    = 0.9             pdiblc1 = 0.078           pdiblc2 = 0.0001        
+ppdiblc2= 3e-015          pdiblcb = 0               drout   = 0.56          
+pvag    = 0               pscbe1  = 6e+008          pscbe2  = 5e-006        
+elm     = 5               agidl   = '6e-012+dagidl_p33_rf'          bgidl   = 7.5255e+008   
+cgidl   = 150             egidl   = 0.5             lagidl  = '0+dlagidl_p33_rf'              
**************************************************************
*               CAPACITANCE PARAMETERS 
**************************************************************
+acde    = 0.5             moin    = 5               noff    = 2             
+voffcv  = 0.01            lvoffcv = -3e-008         cgbo    = 0             
+cgso    = '1e-18'          cgdo    = '1e-18'          cgdl    = 1e-018        
+cgsl    = 1e-18          cf      = 1e-018        clc = 1e-18
**************************************************************
*               TEMPERATURE PARAMETERS 
**************************************************************
+kt1     = -0.33176        pkt1    = 2.9999999e-015  kt1l    = -6.5317e-009  
+kt2     = -0.040277       ute     = -1.2391         wute    = 1.6e-007      
+ua1     = 1.1414e-009     lua1    = -3.0000001e-017  wua1    = 3.9e-016      
+pua1    = -8e-024         ub1     = -3.098e-018     uc1     = 5.8e-012      
+prt     = 0               at      = 3930            lat     = -0.02         
+wat     = 0.055           pat     = -1.9e-008     
**************************************************************
*               NOISE PARAMETERS 
**************************************************************
+noia    = 8.8903E+18      noib    = 1.143E+06      noic    = -2.4438E-13  
+em      = 5.2557E+06         ef      = 1.16281         noimod  = 2             
**************************************************************
*               DIODE PARAMETERS 
**************************************************************
+rsh     = 6.98            js      = 1.82e-007       jsw     = 4e-012        
+cj      = '1e-18'         mj      = 0.378           cjsw    = '1e-18'     
+mjsw    = 0.304           cjswg   = '1e-18'        mjswg   = 0.319         
+pb      = 0.814           pbsw    = 0.923           pbswg   = 0.741         
+rd      = 0               rdc     = 'Rdc_p33/nf'               rs      = 0             
+rsc     = 'Rsc_p33/nf'               xti     = 3.2             tpb     = 0.0015        
+tpbsw   = 0.00073         tpbswg  = 0.0015          tcj     = 0.00078       
+tcjsw   = 0.000911        tcjswg  = 0.000764        acm     = 12            
+calcacm = 1               nj      = 1.0187        
**************************************************************
*               STRESS PARAMETERS 
**************************************************************
+saref   = 3.32e-006       sbref   = 3.32e-006       wlod    = 0             
+kvth0   = 1e-008          lkvth0  = 2.5e-007        wkvth0  = 9e-007        
+pkvth0  = 0               llodvth = 1               wlodvth = 1             
+stk2    = 0               lodk2   = 1               lodeta0 = 1             
+ku0     = 1.915e-007      lku0    = 9.2e-007        wku0    = 2.5e-007      
+pku0    = 0               llodku0 = 1               wlodku0 = 1             
+kvsat   = 0.45            steta0  = 0               tku0    = 0              
*
*
.MODEL pdio33_rf D
+LEVEL    = 3                       JS       = 1.82E-07            JSW      = 1.00E-15  
+N        = 1.0187      RS       = 1.0E-010             IK       = 1.0E+21              
+IKR      = 2.78E+05                BV       = 9.24                  IBV      = 277.8                   
+TRS      = 9.86E-04                EG       = 1.16                  TREF     = 25.0                
+XTI      = 3.0                     TLEV     = 1                     TLEVC    = 1
+CJ       = '1.22E-03+DCJ_P33_RF'   MJ       = 0.378                 PB       = 0.814                
+CJSW     = '4.56E-11+DCJSW_P33_RF' MJSW     = 0.304                 PHP      = 0.923               
+TPB      = 1.50E-03                TPHP     = 7.30E-04              FCS      = 0    
+CTA      = 7.80E-04                CTP      = 9.11E-04              FC       = 0
+AREA     = 3.60E-09                PJ       = 2.40E-04
.ends p33_ckt_rf

