.model nch nmos4 l=1 w=1 n=1
.model pch pmos4 l=1 w=1 n=1