//* No part of this file can be released without the consent of SMIC.
//*
//******************************************************************************************
//* 0.11um Mixed Signal 1P8M with MIM Salicide 1.2V/3.3V RF SPICE Model (for SPECTRE only) *
//******************************************************************************************
//*
//* Release version    : 1.14
//*
//* Release date       : 03/30/2016
//*
//* Simulation tool    : Cadence spectre V6.0
//*
//*
//*  Inductor   :
//*
//*        *---------------------------------------------------------------------------------------------* 
//*        | Inductor subckt |  diff_ind_rf  | diff_ind_rf_pgs | diff_ind_rf_psub | diff_ind_rf_pgs_psub |  
//*        *---------------------------------------------------------------------------------------------*
simulator lang=spectre  insensitive=yes
//*********************************
//* 0.11um differential Inductor
//*********************************
//* 1=port1(M8), 2=port2(M8)
//* R means inner redius; N means turns
//* Spacing is fixed at 1.5um and width is fixed at 8um
subckt diff_ind_rf (1 2) 
parameters r=120e-6 n=3 
+L00    = max((88.81e-12*pwr((r*1e+4),1.29)+12.90e-12)*pwr(n,2)+(128.0e-12*(r*1e+4)-59.23e-12),1e-12)
+R00    = max((0.3257*pwr((r*1e+4),0.9274)+0.1961)*n+(0.09286*(r*1e+4)-0.3465),1e-3)
+L01    = max((61.08e-12*pwr((r*1e+4),2.257)+58.39e-12)*n+(-12.82e-12*pwr((r*1e+4),-0.4249)-83.58e-12),1e-12)
+COXM   = max((31.31e-15*pwr((r*1e+4),0.707)+1.520e-15)*pwr(n,1.2)+(27.95e-15*(r*1e+4)-12.55e-15),1e-18)
+RSM    = max((58.77e+3*pwr((r*1e+6),-1)+13.65)*pwr(n,-1)+(1.091e+3*pwr((r*1e+6),-0.5028)+39.07),1e-3)
+CSM    = 1e-15
+CPASS  = max((15.97e-15*pwr((r*1e+4),1.171)+7.596e-15)*pwr(n,1.2)+(-13.35e-15*pwr((r*1e+4),2.0)-18.82e-15),1e-18)
+COXI   = max((0.2715e-15*pwr((r*1e+4),1.341)+0.5962e-15)*pwr(n,2)+(23.74e-15*pwr((r*1e+4),1.5)+4.7e-15),1e-18)
+RSI    = 300  
+CSI    = max(2.0e-15*pwr(n,1.2)+(77.23e-15*pwr((r*1e+4),0.7531)),1e-18)
+COXO   = COXI
+RSO    = (RSI-5.0)
+CSO    = CSI
+kk     = max((-0.1962*pwr((r*1e+6),0.1493)+0.4354),1e-3)
//* equivalent circuit
l00_rf (1 n1)      inductor     l=(L00*(1+dl00_rf))
r00_rf (n1 nm)     resistor     r=(R00*(1+dr00_rf)) tc1=3.69e-03
l01_rf (n1 n11)    inductor     l=L01
r01_rf (n11 nm)    resistor     r=(R00*2*(1+dr00_rf)) tc1=3.69e-03
l10_rf (nm n2)     inductor     l=(L00*(1+dl00_rf))
r10_rf (n2 2)      resistor     r=(R00*(1+dr00_rf)) tc1=3.69e-03
l11_rf (n2 n21)    inductor     l=L01
r11_rf (n21 2)     resistor     r=(R00*2*(1+dr00_rf)) tc1=3.69e-03
coxm_rf (nm nsm)   capacitor    c=COXM
rsm_rf (nsm 0)     resistor     r=RSM
csm_rf (nsm 0)     capacitor    c=CSM
cpass_rf (1 2)     capacitor    c=CPASS
cci_rf (1 nm)      capacitor    c=0.1e-15
cco_rf (nm 2)      capacitor    c=0.1e-15
rci_rf (nsi nsm)   resistor     r=1e+6
rco_rf (nsm nso)   resistor     r=1e+6
coxi_rf (1 nsi)    capacitor    c=COXI
rsi_rf (nsi 0)     resistor     r=RSI
csi_rf (nsi 0)     capacitor    c=CSI
coxo_rf (2 nso)    capacitor    c=COXO
rso_rf (nso 0)     resistor     r=RSO
cso_rf (nso 0)     capacitor    c=CSO      
k01_rf mutual_inductor coupling=kk ind1=l10_rf ind2=l01_rf
k11_rf mutual_inductor coupling=kk ind1=l00_rf ind2=l11_rf
k12_rf mutual_inductor coupling=0.85 ind1=l00_rf ind2=l10_rf
ka1 mutual_inductor coupling=(kk*0.85) ind1=l01_rf ind2=l00_rf
ka2 mutual_inductor coupling=(kk*0.85) ind1=l11_rf ind2=l10_rf
ends diff_ind_rf
//*
**********************************
* 0.11um differential Inductor with PGS *
**********************************
* 1=port1(M8), 2=port2(M8)
* R means inner redius; N means turns
* Spacing is fixed at 1.5um and width is fixed at 8um
subckt diff_ind_rf_pgs (1 2) 
* inductor scalable model parameters
parameters R=radius N=turns 
+L00  = max((88.81e-12*pwr((R*1e+4),1.29)+12.90e-12)*pwr(N,2)+(128.0e-12*(R*1e+4)-59.23e-12),1e-12)
+R00 = max((0.3257*pwr((R*1e+4),0.9274)+0.1961)*N+(0.09286*(R*1e+4)-0.3465),1e-3)
+L01  = max((61.08e-12*pwr((R*1e+4),2.257)+58.39e-12)*N+(-12.82e-12*pwr((R*1e+4),-0.4249)-83.58e-12),1e-12)
+COXM = max(((31.31e-15*pwr((R*1e+4),0.707)+1.520e-15)*pwr(N,1.2)+(27.95e-15*(R*1e+4)-12.55e-15))*1.16,1e-18)
+RSM = 10
+CSM    = 1e-15
+CPASS = max((15.97e-15*pwr((R*1e+4),1.171)+7.596e-15)*pwr(N,1.2)+(-13.35e-15*pwr((R*1e+4),2.0)-18.82e-15),1e-18)
+COXI  = max(((0.2715e-15*pwr((R*1e+4),1.341)+0.5962e-15)*pwr(N,2)+(23.74e-15*pwr((R*1e+4),1.5)+4.7e-15))*0.95,1e-18)
+RSI = 150  
+CSI    = max(2.0e-15*pwr(N,1.2)+(77.23e-15*pwr((R*1e+4),0.7531)),1e-18)
+COXO  = COXI
+RSO    = RSI-1.0
+CSO    = CSI
+kk = max((-0.1962*pwr((R*1e+6),0.1493)+0.4354),1e-3)
* equivalent circuit
L00_rf  (1 N1)    inductor  l=(L00*(1+dl00_rf)) 
R00_rf  (N1 NM)   resistor  r=(R00*(1+dr00_rf)) tc1=3.69e-03
L01_rf  (N1 N11)  inductor  l=L01 
R01_rf  (N11 NM)  resistor  r=(2.0*R00*(1+dr00_rf)) tc1=3.69e-03
L10_rf  (NM N2)   inductor  l=(L00*(1+dl00_rf))  
R10_rf  (N2 2)    resistor  r=(R00*(1+dr00_rf)) tc1=3.69e-03
L11_rf  (N2 N21)  inductor  l=L01
R11_rf  (N21 2)   resistor  r=(2.0*R00*(1+dr00_rf)) tc1=3.69e-03
COXM_rf  (NM NSM) capacitor c=COXM
RSM_rf  (NSM 0)   resistor  r=RSM  
CSM_rf  (NSM 0)   capacitor c=CSM
CPASS_rf  (1 2)   capacitor c=CPASS 
CCI_rf  (1 NM)    capacitor c=0.1e-15 
CCO_rf  (NM 2)    capacitor c=0.1e-15  
RCI_rf  (NSI NSM) resistor  r=1e+6  
RCO_rf  (NSM NSO) resistor  r=1e+6  
COXI_rf (1 NSI)   capacitor c=COXI
RSI_rf  (NSI 0)   resistor  r=RSI  
CSI_rf  (NSI 0)   capacitor c=CSI 
COXO_rf (2 NSO)   capacitor c=COXO
RSO_rf  (NSO 0)   resistor  r=RSO  
CSO_rf  (NSO 0)   capacitor c=CSO
K01 mutual_inductor coupling=kk ind1=L10_rf ind2=L01_rf 
K11 mutual_inductor coupling=kk ind1=L00_rf ind2=L11_rf
K12 mutual_inductor coupling=0.85 ind1=L00_rf ind2=L10_rf 
ka1 mutual_inductor coupling=(kk*0.85) ind1=L01_rf ind2=L00_rf
ka2 mutual_inductor coupling=(kk*0.85) ind1=L11_rf ind2=L10_rf
ends diff_ind_rf_pgs
//****************************************************
//* 0.11um differential Inductor with psub terminals *
//****************************************************
//* 1=port1(M8), 2=port2(M8)
//* R means inner redius; N means turns
//* Spacing is fixed at 1.5um and width is fixed at 8um
subckt diff_ind_rf_psub (1 2 psub) 
parameters r=120e-6 n=3 
+L00    = max((88.81e-12*pwr((r*1e+4),1.29)+12.90e-12)*pwr(n,2)+(128.0e-12*(r*1e+4)-59.23e-12),1e-12)
+R00    = max((0.3257*pwr((r*1e+4),0.9274)+0.1961)*n+(0.09286*(r*1e+4)-0.3465),1e-3)
+L01    = max((61.08e-12*pwr((r*1e+4),2.257)+58.39e-12)*n+(-12.82e-12*pwr((r*1e+4),-0.4249)-83.58e-12),1e-12)
+COXM   = max((31.31e-15*pwr((r*1e+4),0.707)+1.520e-15)*pwr(n,1.2)+(27.95e-15*(r*1e+4)-12.55e-15),1e-18)
+RSM    = max((58.77e+3*pwr((r*1e+6),-1)+13.65)*pwr(n,-1)+(1.091e+3*pwr((r*1e+6),-0.5028)+39.07),1e-3)
+CSM    = 1e-15
+CPASS  = max((15.97e-15*pwr((r*1e+4),1.171)+7.596e-15)*pwr(n,1.2)+(-13.35e-15*pwr((r*1e+4),2.0)-18.82e-15),1e-18)
+COXI   = max((0.2715e-15*pwr((r*1e+4),1.341)+0.5962e-15)*pwr(n,2)+(23.74e-15*pwr((r*1e+4),1.5)+4.7e-15),1e-18)
+RSI    = 300  
+CSI    = max(2.0e-15*pwr(n,1.2)+(77.23e-15*pwr((r*1e+4),0.7531)),1e-18)
+COXO   = COXI
+RSO    = (RSI-5.0)
+CSO    = CSI
+kk     = max((-0.1962*pwr((r*1e+6),0.1493)+0.4354),1e-3)
//* equivalent circuit
l00_rf (1 n1)      inductor     l=(L00*(1+dl00_rf))
r00_rf (n1 nm)     resistor     r=(R00*(1+dr00_rf)) tc1=3.69e-03
l01_rf (n1 n11)    inductor     l=L01
r01_rf (n11 nm)    resistor     r=(R00*2*(1+dr00_rf)) tc1=3.69e-03
l10_rf (nm n2)     inductor     l=(L00*(1+dl00_rf))
r10_rf (n2 2)      resistor     r=(R00*(1+dr00_rf)) tc1=3.69e-03
l11_rf (n2 n21)    inductor     l=L01
r11_rf (n21 2)     resistor     r=(R00*2*(1+dr00_rf)) tc1=3.69e-03
coxm_rf (nm nsm)   capacitor    c=COXM
rsm_rf (nsm psub)     resistor     r=RSM
csm_rf (nsm psub)     capacitor    c=CSM
cpass_rf (1 2)     capacitor    c=CPASS
cci_rf (1 nm)      capacitor    c=0.1e-15
cco_rf (nm 2)      capacitor    c=0.1e-15
rci_rf (nsi nsm)   resistor     r=1e+6
rco_rf (nsm nso)   resistor     r=1e+6
coxi_rf (1 nsi)    capacitor    c=COXI
rsi_rf (nsi psub)     resistor     r=RSI
csi_rf (nsi psub)     capacitor    c=CSI
coxo_rf (2 nso)    capacitor    c=COXO
rso_rf (nso psub)     resistor     r=RSO
cso_rf (nso psub)     capacitor    c=CSO      
k01_rf mutual_inductor coupling=kk ind1=l10_rf ind2=l01_rf
k11_rf mutual_inductor coupling=kk ind1=l00_rf ind2=l11_rf
k12_rf mutual_inductor coupling=0.85 ind1=l00_rf ind2=l10_rf
ka1 mutual_inductor coupling=(kk*0.85) ind1=l01_rf ind2=l00_rf
ka2 mutual_inductor coupling=(kk*0.85) ind1=l11_rf ind2=l10_rf
ends diff_ind_rf_psub
//*
************************************************************
* 0.11um differential Inductor with PGS and psub terminals *
************************************************************
* 1=port1(M8), 2=port2(M8)
* R means inner redius; N means turns
* Spacing is fixed at 1.5um and width is fixed at 8um
subckt diff_ind_rf_pgs_psub (1 2 psub) 
* inductor scalable model parameters
parameters R=radius N=turns 
+L00  = max((88.81e-12*pwr((R*1e+4),1.29)+12.90e-12)*pwr(N,2)+(128.0e-12*(R*1e+4)-59.23e-12),1e-12)
+R00 = max((0.3257*pwr((R*1e+4),0.9274)+0.1961)*N+(0.09286*(R*1e+4)-0.3465),1e-3)
+L01  = max((61.08e-12*pwr((R*1e+4),2.257)+58.39e-12)*N+(-12.82e-12*pwr((R*1e+4),-0.4249)-83.58e-12),1e-12)
+COXM = max(((31.31e-15*pwr((R*1e+4),0.707)+1.520e-15)*pwr(N,1.2)+(27.95e-15*(R*1e+4)-12.55e-15))*1.16,1e-18)
+RSM = 10
+CSM    = 1e-15
+CPASS = max((15.97e-15*pwr((R*1e+4),1.171)+7.596e-15)*pwr(N,1.2)+(-13.35e-15*pwr((R*1e+4),2.0)-18.82e-15),1e-18)
+COXI  = max(((0.2715e-15*pwr((R*1e+4),1.341)+0.5962e-15)*pwr(N,2)+(23.74e-15*pwr((R*1e+4),1.5)+4.7e-15))*0.95,1e-18)
+RSI = 150  
+CSI    = max(2.0e-15*pwr(N,1.2)+(77.23e-15*pwr((R*1e+4),0.7531)),1e-18)
+COXO  = COXI
+RSO    = RSI-1.0
+CSO    = CSI
+kk = max((-0.1962*pwr((R*1e+6),0.1493)+0.4354),1e-3)
* equivalent circuit
L00_rf  (1 N1)    inductor  l=(L00*(1+dl00_rf)) 
R00_rf  (N1 NM)   resistor  r=(R00*(1+dr00_rf)) tc1=3.69e-03
L01_rf  (N1 N11)  inductor  l=L01 
R01_rf  (N11 NM)  resistor  r=(2.0*R00*(1+dr00_rf)) tc1=3.69e-03
L10_rf  (NM N2)   inductor  l=(L00*(1+dl00_rf))  
R10_rf  (N2 2)    resistor  r=(R00*(1+dr00_rf)) tc1=3.69e-03
L11_rf  (N2 N21)  inductor  l=L01
R11_rf  (N21 2)   resistor  r=(2.0*R00*(1+dr00_rf)) tc1=3.69e-03
COXM_rf  (NM NSM) capacitor c=COXM
RSM_rf  (NSM psub)   resistor  r=RSM  
CSM_rf  (NSM psub)   capacitor c=CSM
CPASS_rf  (1 2)   capacitor c=CPASS 
CCI_rf  (1 NM)    capacitor c=0.1e-15 
CCO_rf  (NM 2)    capacitor c=0.1e-15  
RCI_rf  (NSI NSM) resistor  r=1e+6  
RCO_rf  (NSM NSO) resistor  r=1e+6  
COXI_rf (1 NSI)   capacitor c=COXI
RSI_rf  (NSI psub)   resistor  r=RSI  
CSI_rf  (NSI psub)   capacitor c=CSI 
COXO_rf (2 NSO)   capacitor c=COXO
RSO_rf  (NSO psub)   resistor  r=RSO  
CSO_rf  (NSO psub)   capacitor c=CSO
K01 mutual_inductor coupling=kk ind1=L10_rf ind2=L01_rf 
K11 mutual_inductor coupling=kk ind1=L00_rf ind2=L11_rf
K12 mutual_inductor coupling=0.85 ind1=L00_rf ind2=L10_rf 
ka1 mutual_inductor coupling=(kk*0.85) ind1=L01_rf ind2=L00_rf
ka2 mutual_inductor coupling=(kk*0.85) ind1=L11_rf ind2=L10_rf
ends diff_ind_rf_pgs_psub

