
.subckt diff_opamp dd gnd inp inn net7 out

M1 net1 inn  net3 net3 n33 W={w1} L={l1}
M2 net2 inp  net3 net3 n33 W={w1} L={l1}
M3 net1 net1 dd   dd   p33 W={w2} L={l2} 
M4 net2 net1 dd   dd   p33 W={w2} L={l2}  
M5 net3 net7 gnd  gnd  n33 W={w3} L={l3} 
M6 out  net2 dd   dd   p33 W={w4} L={l4} 
M7 out  net7 gnd  gnd  n33 W={w5} L={l5}
M8 net7 net7 gnd  gnd  n33 W={w3} L={l3}
cc net8 out  {cc}
r1 net2 net8  {cr}

.ends