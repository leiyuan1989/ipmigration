//*Spectre Model Format
simulator lang=spectre  insensitive=yes
ahdl_include "res_rf.va"
// *
// * no part of this file can be released without the consent of smic.
// *****************************************************************************************************
// * SMIC 0.11um Radio Frequency 1P8M(1P7M, 1P6M, 1P5M) Top Metal SPICE Resistor model (for spectre only) *
// *****************************************************************************************************
// *
// * release version    : 1.14
// *
// * release date       : 03/30/2016
// *
// * simulation tool    : Cadence spectre V6.0
// *
// *   resistor         :
// *        *------------------------------------------*
// *        |       resistor type       |      	       |
// *        |==========================================|
// *        |          metal 8(TM2)     |    rtm2_rf   |
// *        |------------------------------------------|
// *        |            ALPA           |    ralpa_rf  |
// *        *------------------------------------------*
// *
// *   the valid temperature range is from -40c to 125c
// *
// ******************************************************************
// *                         resistor model                         *
// ******************************************************************

// ******************************************************************
// *                      metal 8(TM2) resistance                   *
// ******************************************************************
subckt rtm2_rf (n2 n1 sub)  
parameters l=0 w=0 devt=temp    rtc1 = 3.69E-03     rtc2 = -1.8E-08
+ dw = 3.2167E-08+ddw_rtm2_rf         tref = 25           rsh = 7E-03+drsh_rtm2_rf
+ rjc1a = -5.7371E-03             rjc1b = 5.7922E-05
+ rjc2a = 5.785E-05              rjc2b = 9.0221E-07
+ cj = 5.53E-06+dcox_tm2_rf                cjsw = 1.1540E-10+dcapsw_tm2_rf
+ dl = 3.2167E-08+ddw_rtm2_rf  
+ cap = cj*(w*0.9-2.0*dw)*(l*0.9-2.0*dl)/2+cjsw*(w*0.9-2.0*dw+l*0.9-2.0*dl)
C1 (n2 sub) capacitor c = cap
R1 (n2 n1 n2 n1) metalres_rf_hdl lr=l wr=w rtemp=devt etch=dw etchl=dl tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rmaxvcoef=1.10 
C2 (n1 sub) capacitor c = cap
ends rtm2_rf
// ******************************************************************
// *                         ALPA resistance                        *
// ******************************************************************
subckt ralpa_rf (n2 n1 sub)  
parameters l=0 w=0 devt=temp    rtc1 = 3.8865E-03   rtc2 = 5.5735E-08
+ dw = -5.79E-08+ddw_ralpa_rf         tref = 25           rsh = 0.0231+drsh_ralpa_rf
+ rjc1a = 1.9362E-05              rjc1b = -9.0694E-08
+ rjc2a = 1.6459E-05              rjc2b = 2.523E-07
+ cj = 3.53E-06+dcox_alpa_rf                cjsw = 4.649E-11+dcapsw_alpa_rf
+ dl = -5.79E-08+ddw_ralpa_rf  
+ cap = cj*(w*0.9-2.0*dw)*(l*0.9-2.0*dl)/2+cjsw*(w*0.9-2.0*dw+l*0.9-2.0*dl)

C1 (n2 sub) capacitor c = cap
R1 (n2 n1 n2 n1) metalres_rf_hdl lr=l wr=w rtemp=devt etch=dw etchl=dl tc1=rtc1 tc2=rtc2 jc1a=rjc1a jc1b=rjc1b jc2a=rjc2a jc2b=rjc2b rsh0=rsh tnom=tref rmaxvcoef=1.10 
C2 (n1 sub) capacitor c = cap
ends ralpa_rf
