****Sub-Circuit for CLKLAHAQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHAQHSV1 CK E ECK BC VDD VSS
MM51 s c VSS VPW N12LL W=200.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=200.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=260.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=200.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM0 ten BC VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=220.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=320.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=260.00n L=60.00n
MM45 s c nt21 VNW P12LL W=540.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=540.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=500.00n L=60.00n
MM1 ten BC VDD VNW P12LL W=300.00n L=60.00n
MM54 nt21 pm VDD VNW P12LL W=540.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=330.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=460.00n L=60.00n
MM39 pm cn nt11 VNW P12LL W=500.00n L=60.00n
.ENDS CLKLAHAQHSV1
****Sub-Circuit for CLKLAHAQHSV2, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHAQHSV2 CK E ECK BC VDD VSS
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM39 pm cn nt11 VNW P12LL W=440.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=250.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=540.00n L=60.00n
MM45 s c nt21 VNW P12LL W=440.00n L=60.00n
MM54 nt21 pm VDD VNW P12LL W=540.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=540.00n L=60.00n
MM1 ten BC VDD VNW P12LL W=340.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=440.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=350.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=350.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=350.00n L=60.00n
MM51 s c VSS VPW N12LL W=350.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=430.00n L=60.00n
MM0 ten BC VSS VPW N12LL W=270.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=350.00n L=60.00n
.ENDS CLKLAHAQHSV2
****Sub-Circuit for CLKLAHAQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHAQHSV4 CK E ECK BC VDD VSS
MM51 s c VSS VPW N12LL W=300.00n L=60.00n
MM49 m pm VSS VPW N12LL W=300.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=300.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=260.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=300.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM0 ten BC VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=220.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=860.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=260.00n L=60.00n
MM45 s c nt21 VNW P12LL W=600.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=600.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=600.00n L=60.00n
MM1 ten BC VDD VNW P12LL W=300.00n L=60.00n
MM54 nt21 pm VDD VNW P12LL W=590.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=330.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.2u L=60.00n
MM39 pm cn nt11 VNW P12LL W=600.00n L=60.00n
.ENDS CLKLAHAQHSV4
****Sub-Circuit for CLKLAHAQHSV8, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHAQHSV8 CK E ECK BC VDD VSS
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM39 pm cn nt11 VNW P12LL W=540.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=250.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=1.3u L=60.00n
MM45 s c nt21 VNW P12LL W=1.08u L=60.00n
MM54 nt21 pm VDD VNW P12LL W=1.3u L=60.00n
MM21 ECK s VDD VNW P12LL W=2.16u L=60.00n
MM1 ten BC VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=540.00n L=60.00n
MM51 s c VSS VPW N12LL W=860.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=430.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=860.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=860.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=1.72u L=60.00n
MM0 ten BC VSS VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=430.00n L=60.00n
.ENDS CLKLAHAQHSV8
****Sub-Circuit for CLKLAHQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHQHSV1 CK E ECK FC VDD VSS
MM51 hnet12 FC VSS VPW N12LL W=300.00n L=60.00n
MM49 m pm VSS VPW N12LL W=300.00n L=60.00n
MM43 s pm VSS VPW N12LL W=230.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=300.00n L=60.00n
MM44 s c VSS VPW N12LL W=230.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=270n L=60.00n
MM27 cn CK VSS VPW N12LL W=220n L=60.00n
MM22 ECK s VSS VPW N12LL W=340.00n L=60.00n
MM36 pm c hnet12 VPW N12LL W=300.00n L=60.00n
MM45 s c hnet31 VNW P12LL W=550.00n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=550.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=590.0n L=60.00n
MM54 hnet13 FC VDD VNW P12LL W=590.0n L=60.00n
MM14 hnet21 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400n L=60.00n
MM28 cn CK VDD VNW P12LL W=330n L=60.00n
MM21 ECK s VDD VNW P12LL W=440.00n L=60.00n
MM39 pm cn hnet11 VNW P12LL W=590.0n L=60.00n
.ENDS CLKLAHQHSV1
****Sub-Circuit for CLKLAHQHSV2, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHQHSV2 CK E ECK FC VDD VSS
MM22 ECK s VSS VPW N12LL W=430.00n L=60.00n
MM44 s c VSS VPW N12LL W=270.00n L=60.00n
MM43 s pm VSS VPW N12LL W=270.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM51 hnet12 FC VSS VPW N12LL W=350.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=350.00n L=60.00n
MM36 pm c hnet12 VPW N12LL W=350.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270n L=60.00n
MM30 c cn VSS VPW N12LL W=350n L=60.00n
MM21 ECK s VDD VNW P12LL W=540.00n L=60.00n
MM45 s c hnet31 VNW P12LL W=500.00n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=500.00n L=60.00n
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM14 hnet21 c pm VNW P12LL W=250.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=250.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=440.0n L=60.00n
MM39 pm cn hnet11 VNW P12LL W=440.0n L=60.00n
MM54 hnet13 FC VDD VNW P12LL W=440.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=340n L=60.00n
MM29 c cn VDD VNW P12LL W=440n L=60.00n
.ENDS CLKLAHQHSV2
****Sub-Circuit for CLKLAHQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHQHSV4 CK E ECK FC VDD VSS
MM51 hnet12 FC VSS VPW N12LL W=340.00n L=60.00n
MM49 m pm VSS VPW N12LL W=400.00n L=60.00n
MM43 s pm VSS VPW N12LL W=280.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=340.00n L=60.00n
MM44 s c VSS VPW N12LL W=280.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=270n L=60.00n
MM27 cn CK VSS VPW N12LL W=220n L=60.00n
MM22 ECK s VSS VPW N12LL W=860n L=60.00n
MM36 pm c hnet12 VPW N12LL W=340.00n L=60.00n
MM45 s c hnet31 VNW P12LL W=640.00n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=640.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=650.0n L=60.00n
MM54 hnet13 FC VDD VNW P12LL W=650.0n L=60.00n
MM14 hnet21 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400n L=60.00n
MM28 cn CK VDD VNW P12LL W=330n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.2u L=60.00n
MM39 pm cn hnet11 VNW P12LL W=650.0n L=60.00n
.ENDS CLKLAHQHSV4
****Sub-Circuit for CLKLAHQHSV8, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHQHSV8 CK E ECK FC VDD VSS
MM22 ECK s VSS VPW N12LL W=1.72u L=60.00n
MM44 s c VSS VPW N12LL W=580.00n L=60.00n
MM43 s pm VSS VPW N12LL W=580.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM51 hnet12 FC VSS VPW N12LL W=430.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=430.00n L=60.00n
MM36 pm c hnet12 VPW N12LL W=430.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270n L=60.00n
MM30 c cn VSS VPW N12LL W=430n L=60.00n
MM21 ECK s VDD VNW P12LL W=2.16u L=60.00n
MM45 s c hnet31 VNW P12LL W=1080n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=1080n L=60.00n
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM14 hnet21 c pm VNW P12LL W=250.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=250.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=540.00n L=60.00n
MM39 pm cn hnet11 VNW P12LL W=540.00n L=60.00n
MM54 hnet13 FC VDD VNW P12LL W=540.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340n L=60.00n
MM29 c cn VDD VNW P12LL W=540n L=60.00n
.ENDS CLKLAHQHSV8
****Sub-Circuit for CLKLANAQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANAQHSV1 CK E ECK BC VDD VSS
MM51 nt22 BC VSS VPW N12LL W=300.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c nt22 VPW N12LL W=300.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=260.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=300.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=290.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=260.00n L=60.00n
MM45 s m nt21 VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=400.00n L=60.00n
MM54 nt21 BC VDD VNW P12LL W=300.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=360.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=460.00n L=60.00n
MM39 pm c nt11 VNW P12LL W=400.00n L=60.00n
.ENDS CLKLANAQHSV1
****Sub-Circuit for CLKLANAQHSV2, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT CLKLANAQHSV2 CK E ECK BC VDD VSS
MM39 pm c nt11 VNW P12LL W=440.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=440.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=250.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM50 m pm VDD VNW P12LL W=350.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM29 c cn VDD VNW P12LL W=430.00n L=60.00n
MM54 nt21 BC VDD VNW P12LL W=350.00n L=60.00n
MM45 s m nt21 VNW P12LL W=350.00n L=60.00n
MM46 s c VDD VNW P12LL W=350.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=540.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=350.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=350.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM49 m pm VSS VPW N12LL W=280.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=350.00n L=60.00n
MM51 nt22 BC VSS VPW N12LL W=350.00n L=60.00n
MM43 s c nt22 VPW N12LL W=350.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=430.00n L=60.00n
.ENDS CLKLANAQHSV2
****Sub-Circuit for CLKLANAQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANAQHSV4 CK E ECK BC VDD VSS
MM51 nt22 BC VSS VPW N12LL W=430.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c nt22 VPW N12LL W=430.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=320.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=270.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=800.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=320.00n L=60.00n
MM45 s m nt21 VNW P12LL W=430.00n L=60.00n
MM46 s c VDD VNW P12LL W=430.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=450.00n L=60.00n
MM54 nt21 BC VDD VNW P12LL W=430.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=360.00n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.3u L=60.00n
MM39 pm c nt11 VNW P12LL W=450.00n L=60.00n
.ENDS CLKLANAQHSV4
****Sub-Circuit for CLKLANAQHSV8, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT CLKLANAQHSV8 CK E ECK BC VDD VSS
MM21 ECK s VDD VNW P12LL W=2.16u L=60.00n
MM46 s c VDD VNW P12LL W=860.00n L=60.00n
MM45 s m nt21 VNW P12LL W=860.00n L=60.00n
MM54 nt21 BC VDD VNW P12LL W=860.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM50 m pm VDD VNW P12LL W=540.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=250.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=540.00n L=60.00n
MM39 pm c nt11 VNW P12LL W=540.00n L=60.00n
MM43 s c nt22 VPW N12LL W=860.00n L=60.00n
MM22 ECK s VSS VPW N12LL W=1.72u L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM51 nt22 BC VSS VPW N12LL W=860.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=860.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM49 m pm VSS VPW N12LL W=430.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=430.00n L=60.00n
.ENDS CLKLANAQHSV8
****Sub-Circuit for CLKLANQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV1 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK s VSS VPW N12LL W=290.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK s VDD VNW P12LL W=460.00n L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV1
****Sub-Circuit for CLKLANQHSV12, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV12 CK E ECK FC VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=860.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK pq VSS VPW N12LL W=2.46u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.2u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK pq VDD VNW P12LL W=3.9u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV12
****Sub-Circuit for CLKLANQHSV16, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV16 CK E ECK FC VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=860.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK pq VSS VPW N12LL W=3.42u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.2u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK pq VDD VNW P12LL W=5.2u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV16
****Sub-Circuit for CLKLANQHSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV2 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK s VSS VPW N12LL W=420.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK s VDD VNW P12LL W=650.00n L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV2
****Sub-Circuit for CLKLANQHSV20, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV20 CK E ECK FC VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=1.29u L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK pq VSS VPW N12LL W=4.2u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.74u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK pq VDD VNW P12LL W=6.5u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV20
****Sub-Circuit for CLKLANQHSV24, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV24 CK E ECK FC VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=1.29u L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK pq VSS VPW N12LL W=5.16u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.74u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK pq VDD VNW P12LL W=7.8u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV24
****Sub-Circuit for CLKLANQHSV3, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV3 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=360.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=360.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK s VSS VPW N12LL W=620.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=400.00n L=60.00n
MM46 s c VDD VNW P12LL W=400.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK s VDD VNW P12LL W=960.00n L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV3
****Sub-Circuit for CLKLANQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV4 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=430.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=260n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 ECK s VSS VPW N12LL W=800.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=500.00n L=60.00n
MM46 s c VDD VNW P12LL W=500.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.3u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV4
****Sub-Circuit for CLKLANQHSV6, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV6 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=340.00n L=60.00n
MM49 m pm VSS VPW N12LL W=380.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=430.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=340.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=360n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM22 ECK s VSS VPW N12LL W=1.14u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=340.00n L=60.00n
MM45 s m VDD VNW P12LL W=440.00n L=60.00n
MM46 s c VDD VNW P12LL W=440.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=600.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=600.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540n L=60.00n
MM28 cn CK VDD VNW P12LL W=450n L=60.00n
MM21 ECK s VDD VNW P12LL W=1.95u L=60.00n
MM39 pm c hnet24 VNW P12LL W=600.0n L=60.00n
.ENDS CLKLANQHSV6
****Sub-Circuit for CLKLANQHSV8, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV8 CK E ECK FC VDD VSS
MM51 hnet22 FC VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=360.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=740.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=740.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=360n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM22 ECK s VSS VPW N12LL W=1.6u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=800.0n L=60.00n
MM46 s c VDD VNW P12LL W=800.0n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 FC VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540n L=60.00n
MM28 cn CK VDD VNW P12LL W=450n L=60.00n
MM21 ECK s VDD VNW P12LL W=2.6u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV8

****Sub-Circuit for LAHHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHHSV1 D G Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 c pm VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=400.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHHSV1
****Sub-Circuit for LAHHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHHSV2 D G Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 c pm VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=570.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=570.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LAHHSV2
****Sub-Circuit for LAHHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHHSV4 D G Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 c pm VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=650.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LAHHSV4
****Sub-Circuit for LAHRNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRNHSV1 D G Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=340.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=340.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=600.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=560.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=560.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHRNHSV1
****Sub-Circuit for LAHRNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRNHSV2 D G Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=410.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=390.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=410.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=560.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=560.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHRNHSV2
****Sub-Circuit for LAHRNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRNHSV4 D G Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net117 cn pm VNW P12LL W=350.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=350.00n L=60.00n
MM10 pm c net128 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LAHRNHSV4
****Sub-Circuit for LAHRSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRSNHSV1 D G Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=330.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=330.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=330.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHRSNHSV1
****Sub-Circuit for LAHRSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRSNHSV2 D G Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LAHRSNHSV2
****Sub-Circuit for LAHRSNHSV4, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT LAHRSNHSV4 D G Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM51 pm s VSS VPW N12LL W=240.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=360.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=650.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=640.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=640.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=510.00n L=60.00n
.ENDS LAHRSNHSV4
****Sub-Circuit for LAHSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHSNHSV1 D G Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=290.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c G VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 c net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c G VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=430.00n L=60.00n
MM47 Q net0127 VDD VNW P12LL W=430.00n L=60.00n
MM14 net0285 cn net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 c net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHSNHSV1
****Sub-Circuit for LAHSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHSNHSV2 D G Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=430.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 c net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 cn net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q net0127 VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 cn net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 c net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=440.00n L=60.00n
.ENDS LAHSNHSV2
****Sub-Circuit for LAHSNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHSNHSV4 D G Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=860.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=405.00n L=60.00n
MM27 c G VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 c net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=320.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=650.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c G VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q net0127 VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 cn net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 c net0292 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=510.00n L=60.00n
.ENDS LAHSNHSV4
****Sub-Circuit for LALHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALHSV1 D GN Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=400.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALHSV1
****Sub-Circuit for LALHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALHSV2 D GN Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=570.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=570.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LALHSV2
****Sub-Circuit for LALHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALHSV4 D GN Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=650.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LALHSV4
****Sub-Circuit for LALRNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRNHSV1 D GN Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=230.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=230.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=230.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=200.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS LALRNHSV1
****Sub-Circuit for LALRNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRNHSV2 D GN Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=310.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=390.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=310.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net117 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net128 VNW P12LL W=560.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=560.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALRNHSV2
****Sub-Circuit for LALRNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRNHSV4 D GN Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=380.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net117 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net128 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LALRNHSV4
****Sub-Circuit for LALRSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRSNHSV1 D GN Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=330.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=330.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=330.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALRSNHSV1
****Sub-Circuit for LALRSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRSNHSV2 D GN Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM51 pm s VSS VPW N12LL W=200.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=550.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=250.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LALRSNHSV2
****Sub-Circuit for LALRSNHSV4, Mon May 30 19:34:53 CST 2011****
.SUBCKT LALRSNHSV4 D GN Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0145 VSS VPW N12LL W=860.00n L=60.00n
MM51 net0145 s VSS VPW N12LL W=200.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=360.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 cn net0145 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 net0145 c net69 VPW N12LL W=420.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=420.00n L=60.00n
MM0 net_0154 net0145 VSS VPW N12LL W=360.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM52 net0145 s net0252 VNW P12LL W=290.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=290.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=640.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q net0145 VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 c net0145 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0145 cn net0292 VNW P12LL W=605.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=550.00n L=60.00n
MM1 net_0154 net0145 VDD VNW P12LL W=510.00n L=60.00n
.ENDS LALRSNHSV4
****Sub-Circuit for LALSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALSNHSV1 D GN Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c GN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c GN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALSNHSV1
****Sub-Circuit for LALSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALSNHSV2 D GN Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=430.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 cn net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 c net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q net0127 VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 c net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 cn net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=440.00n L=60.00n
.ENDS LALSNHSV2
****Sub-Circuit for LALSNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALSNHSV4 D GN Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=860.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c GN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 cn net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 c net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=320.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=650.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c GN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q net0127 VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 c net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 cn net0292 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=510.00n L=60.00n
.ENDS LALSNHSV4

***********************************************************

****Sub-Circuit for DGRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNHSV1 CK D Q QN RN VDD VSS
MM39 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM3 m c net43 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=250.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=250.00n L=60.00n
MM0 m pm VSS VPW N12LL W=340.00n L=60.00n
MM40 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM4 m cn net43 VNW P12LL W=500.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=330.00n L=60.00n
MM1 m pm VDD VNW P12LL W=500.00n L=60.00n
.ENDS DGRNHSV1
****Sub-Circuit for DGRNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNHSV2 CK D Q QN RN VDD VSS
MM39 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM3 m c net43 VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM40 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM4 m cn net43 VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=450.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS DGRNHSV2
****Sub-Circuit for DGRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNHSV4 CK D Q QN RN VDD VSS
MM39 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM3 m c net43 VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=360.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 m pm VSS VPW N12LL W=390.00n L=60.00n
MM40 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM4 m cn net43 VNW P12LL W=580.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=540.0n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=580.00n L=60.00n
.ENDS DGRNHSV4
****Sub-Circuit for DGRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNQHSV1 CK D Q RN VDD VSS
MM3 m c net43 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=250.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=250.00n L=60.00n
MM0 m pm VSS VPW N12LL W=340.00n L=60.00n
MM4 m cn net43 VNW P12LL W=500.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=330.00n L=60.00n
MM1 m pm VDD VNW P12LL W=500.00n L=60.00n
.ENDS DGRNQHSV1
****Sub-Circuit for DGRNQHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT DGRNQHSV2 CK D Q RN VDD VSS
MM3 m c net43 VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=270.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=270.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM4 m cn net43 VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=450.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=350.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS DGRNQHSV2
****Sub-Circuit for DGRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNQHSV4 CK D Q RN VDD VSS
MM3 m c net43 VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=340.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=270.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=270.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM4 m cn net43 VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.0n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=350.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS DGRNQHSV4
****Sub-Circuit for DGRSNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRSNHSV1 CK D Q QN RN SN VDD VSS
MM43 snn SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN net073 VSS VPW N12LL W=290.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=340.00n L=60.00n
MM42 net69 snn net_0162 VPW N12LL W=250.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=250.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=290.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=250.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=340.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=450.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=380.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=440.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=500.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=440.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=380.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=380.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=500.00n L=60.00n
.ENDS DGRSNHSV1
****Sub-Circuit for DGRSNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRSNHSV2 CK D Q QN RN SN VDD VSS
MM43 snn SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN net073 VSS VPW N12LL W=430.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=360.00n L=60.00n
MM42 net69 snn net_0162 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=430.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=360.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=450.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=650.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=650.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGRSNHSV2
****Sub-Circuit for DGRSNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRSNHSV4 CK D Q QN RN SN VDD VSS
MM43 snn SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN net073 VSS VPW N12LL W=860.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=360.00n L=60.00n
MM42 net69 snn net_0162 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=860.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=360.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=450.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=1.3u L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=1.3u L=60.00n
MM18 net063 net073 VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGRSNHSV4
****Sub-Circuit for DGSNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGSNHSV1 CK D Q QN SN VDD VSS
MM39 QN net073 VSS VPW N12LL W=290.00n L=60.00n
MM43 snn SN VSS VPW N12LL W=200.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=270.00n L=60.00n
MM42 net69 snn VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=290.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=250.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=270.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=440.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=440.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=300.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=440.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=440.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=400.00n L=60.00n
.ENDS DGSNHSV1
****Sub-Circuit for DGSNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGSNHSV2 CK D Q QN SN VDD VSS
MM39 QN net073 VSS VPW N12LL W=430.00n L=60.00n
MM43 snn SN VSS VPW N12LL W=200.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=350.00n L=60.00n
MM42 net69 snn VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=380.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=430.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=260.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=260.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=350.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=650.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=300.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=570.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=650.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGSNHSV2
****Sub-Circuit for DGSNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGSNHSV4 CK D Q QN SN VDD VSS
MM39 QN net073 VSS VPW N12LL W=860.00n L=60.00n
MM43 snn SN VSS VPW N12LL W=200.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=340.00n L=60.00n
MM42 net69 snn VSS VPW N12LL W=250.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=860.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=270.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=270.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=340.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=1.3u L=60.00n
MM44 snn SN VDD VNW P12LL W=300.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=1.3u L=60.00n
MM18 net063 net073 VDD VNW P12LL W=490.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGSNHSV4
****Sub-Circuit for DHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DHSV1 CK D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=290.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM43 QN s VDD VNW P12LL W=440.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DHSV1
****Sub-Circuit for DHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DHSV2 CK D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=430.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=640.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=640.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DHSV2
****Sub-Circuit for DHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DHSV4 CK D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 net43 c net_099 VPW N12LL W=300.00n L=60.00n m=2
MM40 net_099 m VSS VPW N12LL W=300.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM17 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 net43 cn net_0158 VNW P12LL W=450.00n L=60.00n m=2
MM41 net_0158 m VDD VNW P12LL W=450.00n L=60.00n m=2
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM18 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DHSV4
****Sub-Circuit for DQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DQHSV1 CK D Q VDD VSS
MM39 net43 c net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS DQHSV1
****Sub-Circuit for DQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DQHSV2 CK D Q VDD VSS
MM39 net43 c net_099 VPW N12LL W=430.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=290.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=290.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=440.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=440.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DQHSV2
****Sub-Circuit for DQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DQHSV4 CK D Q VDD VSS
MM39 net43 c net_099 VPW N12LL W=600.0n L=60.00n
MM40 net_099 m VSS VPW N12LL W=600.0n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=290.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=290.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=910.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=910.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=440.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=440.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DQHSV4
****Sub-Circuit for DRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNHSV1 CK D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DRNHSV1
****Sub-Circuit for DRNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNHSV2 CK D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNHSV2
****Sub-Circuit for DRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNHSV4 CK D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=330.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=330.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNHSV4
****Sub-Circuit for DRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNQHSV1 CK D Q RDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DRNQHSV1
****Sub-Circuit for DRNQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNQHSV2 CK D Q RDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNQHSV2
****Sub-Circuit for DRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNQHSV4 CK D Q RDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=330.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=330.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNQHSV4
****Sub-Circuit for DRSNHSV1, Mon May 30 16:01:10 CST 2011****
.SUBCKT DRSNHSV1 CK D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=290.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=220.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=220.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=360.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=440.00n L=60.00n
.ENDS DRSNHSV1
****Sub-Circuit for DRSNHSV2, Mon May 30 19:07:49 CST 2011****
.SUBCKT DRSNHSV2 CK D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=360.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=380.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=400.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=390.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=220.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=220.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=400.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=600.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=600.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=600.00n L=60.00n
.ENDS DRSNHSV2
****Sub-Circuit for DRSNHSV4, Mon May 30 19:07:49 CST 2011****
.SUBCKT DRSNHSV4 CK D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=360.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=410.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n m=2
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=320.00n L=60.00n m=2
MM40 net43 R net_0132 VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=220.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=220.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 s net43 VDD VNW P12LL W=600.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=650.00n L=60.00n m=2
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=290.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=290.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=630.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=650.00n L=60.00n
.ENDS DRSNHSV4
****Sub-Circuit for DSNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DSNHSV1 CK D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=400.00n L=60.00n
.ENDS DSNHSV1
****Sub-Circuit for DSNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DSNHSV2 CK D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=300.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=390.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS DSNHSV2
****Sub-Circuit for DSNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DSNHSV4 CK D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=780.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=780.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM38 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=570.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=910.00n L=60.00n
.ENDS DSNHSV4
****Sub-Circuit for DXHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DXHSV1 CK DA DB Q QN SA VDD VSS
MM33 m c net43 VPW N12LL W=350.00n L=60.00n
MM16 net_0144 DB VSS VPW N12LL W=350.00n L=60.00n
MM31 san SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=350.00n L=60.00n
MM19 QN s VSS VPW N12LL W=350.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=310.00n L=60.00n
MM3 net_0148 SA n43 VPW N12LL W=240.00n L=60.00n
MM7 net69 n43 VSS VPW N12LL W=310.00n L=60.00n
MM5 net_0144 san n43 VPW N12LL W=240.00n L=60.00n
MM2 net_0148 DA VSS VPW N12LL W=350.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM38 m cn net43 VNW P12LL W=440.00n L=60.00n
MM37 net_0144 DB VDD VNW P12LL W=440.00n L=60.00n
MM15 net_0148 DA VDD VNW P12LL W=440.00n L=60.00n
MM32 san SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM20 QN s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 n43 VDD VNW P12LL W=390.00n L=60.00n
MM4 net_0148 san n43 VNW P12LL W=300.00n L=60.00n
MM6 net_0144 SA n43 VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DXHSV1
****Sub-Circuit for DXHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DXHSV2 CK DA DB Q QN SA VDD VSS
MM5 net_0150 san n43 VPW N12LL W=240.00n L=60.00n
MM2 net_0138 DA VSS VPW N12LL W=350.00n L=60.00n
MM31 san SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM19 QN s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM33 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=310.00n L=60.00n
MM16 net_0150 DB VSS VPW N12LL W=350.00n L=60.00n
MM7 net69 n43 VSS VPW N12LL W=430.00n L=60.00n
MM3 net_0138 SA n43 VPW N12LL W=240.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM15 net_0138 DA VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0150 DB VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0138 san n43 VNW P12LL W=300.00n L=60.00n
MM6 net_0150 SA n43 VNW P12LL W=300.00n L=60.00n
MM32 san SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=550.00n L=60.00n
MM20 QN s VDD VNW P12LL W=550.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 m cn net43 VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 n43 VDD VNW P12LL W=550.00n L=60.00n
MM1 m pm VDD VNW P12LL W=550.00n L=60.00n
.ENDS DXHSV2
****Sub-Circuit for DXHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DXHSV4 CK DA DB Q QN SA VDD VSS
MM2 net_0156 DA VSS VPW N12LL W=350.00n L=60.00n
MM5 net_0144 san n43 VPW N12LL W=240.00n L=60.00n
MM3 net_0156 SA n43 VPW N12LL W=240.00n L=60.00n
MM16 net_0144 DB VSS VPW N12LL W=350.00n L=60.00n
MM31 san SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM19 QN s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM33 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=260.00n L=60.00n
MM7 net69 n43 VSS VPW N12LL W=260.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM6 net_0144 SA n43 VNW P12LL W=300.00n L=60.00n
MM4 net_0156 san n43 VNW P12LL W=300.00n L=60.00n
MM15 net_0156 DA VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0144 DB VDD VNW P12LL W=440.00n L=60.00n
MM32 san SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.1u L=60.00n
MM20 QN s VDD VNW P12LL W=1.1u L=60.00n
MM18 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM38 m cn net43 VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 n43 VDD VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=550.00n L=60.00n
.ENDS DXHSV4
****Sub-Circuit for EDGRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNHSV1 CK D E Q QN RN VDD VSS
MM43 QN s VSS VPW N12LL W=290.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=280.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=280.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM44 QN s VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNHSV1
****Sub-Circuit for EDGRNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNHSV2 CK D E Q QN RN VDD VSS
MM43 QN s VSS VPW N12LL W=390.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=390.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM44 QN s VDD VNW P12LL W=610.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=610.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=440.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNHSV2
****Sub-Circuit for EDGRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNHSV4 CK D E Q QN RN VDD VSS
MM43 QN s VSS VPW N12LL W=860.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=260.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=260.00n L=60.00n
MM44 QN s VDD VNW P12LL W=1.3u L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=500.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=400.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=400.00n L=60.00n
.ENDS EDGRNHSV4
****Sub-Circuit for EDGRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNQHSV1 CK D E Q RN VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=300.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=280.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=280.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=415.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNQHSV1
****Sub-Circuit for EDGRNQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNQHSV2 CK D E Q RN VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=420.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=420.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=440.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNQHSV2
****Sub-Circuit for EDGRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNQHSV4 CK D E Q RN VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=300.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.0n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=450.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=440.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNQHSV4
****Sub-Circuit for EDHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDHSV1 CK D E Q QN VDD VSS
MM43 QN s VSS VPW N12LL W=290.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=395.00n L=60.00n
MM42 QN s VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=495.00n L=60.00n
.ENDS EDHSV1
****Sub-Circuit for EDHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT EDHSV2 CK D E Q QN VDD VSS
MM43 QN s VSS VPW N12LL W=430.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=340.00n L=60.00n
MM42 QN s VDD VNW P12LL W=650.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=400.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=400.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=550.00n L=60.00n
.ENDS EDHSV2
****Sub-Circuit for EDHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDHSV4 CK D E Q QN VDD VSS
MM43 QN s VSS VPW N12LL W=860.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 QN s VDD VNW P12LL W=1.3u L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDHSV4
****Sub-Circuit for EDQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDQHSV1 CK D E Q VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=395.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=495.00n L=60.00n
.ENDS EDQHSV1
****Sub-Circuit for EDQHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT EDQHSV2 CK D E Q VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=340.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=400.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=400.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=550.00n L=60.00n
.ENDS EDQHSV2
****Sub-Circuit for EDQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDQHSV4 CK D E Q VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDQHSV4
****Sub-Circuit for EDRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNHSV1 CK D E Q QN RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM47 QN s VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM48 QN s VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=320.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=320.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNHSV1
****Sub-Circuit for EDRNHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT EDRNHSV2 CK D E Q QN RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM47 QN s VSS VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM48 QN s VDD VNW P12LL W=650.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=430.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=430.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNHSV2
****Sub-Circuit for EDRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNHSV4 CK D E Q QN RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM47 QN s VSS VPW N12LL W=860.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM48 QN s VDD VNW P12LL W=1.3u L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNHSV4
****Sub-Circuit for EDRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNQHSV1 CK D E Q RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=320.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=320.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNQHSV1
****Sub-Circuit for EDRNQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNQHSV2 CK D E Q RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=430.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=430.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNQHSV2
****Sub-Circuit for EDRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNQHSV4 CK D E Q RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNQHSV4



****Sub-Circuit for NDHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDHSV1 CKN D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=290.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM43 QN s VDD VNW P12LL W=440.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDHSV1
****Sub-Circuit for NDHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDHSV2 CKN D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=230.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=230.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=480.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDHSV2
****Sub-Circuit for NDHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDHSV4 CKN D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 net43 c net_099 VPW N12LL W=400.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=400.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM17 s net43 VSS VPW N12LL W=400.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 net43 cn net_0158 VNW P12LL W=450.00n L=60.00n m=2
MM41 net_0158 m VDD VNW P12LL W=450.00n L=60.00n m=2
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM18 s net43 VDD VNW P12LL W=600.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDHSV4
****Sub-Circuit for NDRNHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRNHSV1 CKN D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=200.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=200.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS NDRNHSV1
****Sub-Circuit for NDRNHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRNHSV2 CKN D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=200.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=300.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=200.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS NDRNHSV2
****Sub-Circuit for NDRNHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRNHSV4 CKN D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM3 net_0154 c net43 VPW N12LL W=360.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=200.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=190.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=280.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=280.00n L=60.00n m=2
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=190.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=190.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=260.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=560n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=650.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=610.00n L=60.00n
.ENDS NDRNHSV4
****Sub-Circuit for NDRSNHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRSNHSV1 CKN D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=200.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=200.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=380.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=440.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=350.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=440.00n L=60.00n
.ENDS NDRSNHSV1
****Sub-Circuit for NDRSNHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRSNHSV2 CKN D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=250.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=260.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=240.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=250.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=250.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=240.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=320.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=460.00n L=60.00n m=1
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=650.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=580.00n L=60.00n
.ENDS NDRSNHSV2
****Sub-Circuit for NDRSNHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRSNHSV4 CKN D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=260.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=240.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=420.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=240.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 s net43 VDD VNW P12LL W=470.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=460n L=60.00n
MM29 cn c VDD VNW P12LL W=640.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=650.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=430.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=620.00n L=60.00n
.ENDS NDRSNHSV4
****Sub-Circuit for NDSNHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDSNHSV1 CKN D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=290.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=270.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=290.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDSNHSV1
****Sub-Circuit for NDSNHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDSNHSV2 CKN D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=260.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=390.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=390.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=395.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=395.00n L=60.00n
.ENDS NDSNHSV2
****Sub-Circuit for NDSNHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDSNHSV4 CKN D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=390.00n L=60.00n
MM30 cn c VSS VPW N12LL W=400.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=400.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 s net43 VDD VNW P12LL W=580.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=600.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=600.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=620.00n L=60.00n
.ENDS NDSNHSV4


***********************************************************


****Sub-Circuit for SDGRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNHSV1 CK D Q QN RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM52 QN ps VSS VPW N12LL W=290.00n L=60.00n
MM3 m c ps VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=410.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=270.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=410.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM53 QN ps VDD VNW P12LL W=440.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=530.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=410.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=530.00n L=60.00n
MM1 m pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS SDGRNHSV1
****Sub-Circuit for SDGRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNHSV2 CK D Q QN RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM52 QN ps VSS VPW N12LL W=430.00n L=60.00n
MM3 m c ps VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=410.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=340.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=270.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=410.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM53 QN ps VDD VNW P12LL W=650.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=530.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=410.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=530.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRNHSV2
****Sub-Circuit for SDGRNHSV4, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT SDGRNHSV4 CK D Q QN RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM52 QN ps VSS VPW N12LL W=860.00n L=60.00n
MM3 m c ps VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=360.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=410.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=270.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=410.00n L=60.00n
MM0 m pm VSS VPW N12LL W=390.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM53 QN ps VDD VNW P12LL W=1.3u L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=540.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=530.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=410.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=530.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRNHSV4
****Sub-Circuit for SDGRNQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNQHSV1 CK D Q RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM3 m c ps VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=380.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=250.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=380.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=530.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=500.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=380.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS SDGRNQHSV1
****Sub-Circuit for SDGRNQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNQHSV2 CK D Q RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM3 m c ps VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=330.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=330.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=380.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=340.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=250.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=380.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=500.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=380.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRNQHSV2
****Sub-Circuit for SDGRNQHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SDGRNQHSV4 CK D Q RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM3 m c ps VPW N12LL W=370.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=360.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=380.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=250.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=380.00n L=60.00n
MM0 m pm VSS VPW N12LL W=390.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=540.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=500.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=360.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=580.00n L=60.00n
.ENDS SDGRNQHSV4
****Sub-Circuit for SDGRSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRSNHSV1 CK D Q QN RN SE SI SN VDD VSS
MM45 net0370 SE net201 VPW N12LL W=300.00n L=60.00n
MM46 net201 SI VSS VPW N12LL W=300.00n L=60.00n
MM47 net0172 RN VSS VPW N12LL W=390.00n L=60.00n
MM48 net0370 SEN net213 VPW N12LL W=340.00n L=60.00n
MM49 net213 D net205 VPW N12LL W=390.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN OS VSS VPW N12LL W=290.00n L=60.00n
MM62 OS c net181 VPW N12LL W=260.00n L=60.00n
MM63 net181 S VSS VPW N12LL W=260.00n L=60.00n
MM61 M cn net193 VPW N12LL W=300.00n L=60.00n
MM58 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM70 net205 SN net0172 VPW N12LL W=390.00n L=60.00n
MM60 net193 net0370 VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=230.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=230.00n L=60.00n
MM24 net172 cn OS VPW N12LL W=200.00n L=60.00n
MM23 VSS NET64 net172 VPW N12LL W=200.00n L=60.00n
MM69 net213 SNN net0172 VPW N12LL W=300.00n L=60.00n
MM19 Q NET64 VSS VPW N12LL W=290.00n L=60.00n
MM17 NET64 OS VSS VPW N12LL W=260.00n L=60.00n
MM12 net240 c M VPW N12LL W=200.00n L=60.00n
MM11 VSS S net240 VPW N12LL W=200.00n L=60.00n
MM0 S M VSS VPW N12LL W=300.00n L=60.00n
MM66 net0418 SNN net296 VNW P12LL W=590.00n L=60.00n
MM50 net288 SI VDD VNW P12LL W=420.00n L=60.00n
MM51 net0370 SEN net288 VNW P12LL W=420.00n L=60.00n
MM52 net296 D VDD VNW P12LL W=590.00n L=60.00n
MM53 net0370 SE net0418 VNW P12LL W=590.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=450.00n L=60.00n
MM40 QN OS VDD VNW P12LL W=440.00n L=60.00n
MM64 net268 S VDD VNW P12LL W=390.00n L=60.00n
MM65 OS cn net268 VNW P12LL W=390.00n L=60.00n
MM67 net0418 RN VDD VNW P12LL W=450.00n L=60.00n
MM59 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=360.00n L=60.00n
MM26 VDD NET64 net253 VNW P12LL W=300.00n L=60.00n
MM25 net253 c OS VNW P12LL W=300.00n L=60.00n
MM20 Q NET64 VDD VNW P12LL W=440.00n L=60.00n
MM18 NET64 OS VDD VNW P12LL W=390.00n L=60.00n
MM14 net313 cn M VNW P12LL W=300.00n L=60.00n
MM13 VDD S net313 VNW P12LL W=300.00n L=60.00n
MM55 net280 net0370 VDD VNW P12LL W=450.00n L=60.00n
MM56 M c net280 VNW P12LL W=450.00n L=60.00n
MM1 S M VDD VNW P12LL W=450.00n L=60.00n
.ENDS SDGRSNHSV1
****Sub-Circuit for SDGRSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRSNHSV2 CK D Q QN RN SE SI SN VDD VSS
MM45 net0370 SE net201 VPW N12LL W=270.00n L=60.00n
MM46 net201 SI VSS VPW N12LL W=270.00n L=60.00n
MM47 net0172 RN VSS VPW N12LL W=350.00n L=60.00n
MM48 net0370 SEN net213 VPW N12LL W=350.00n L=60.00n
MM49 net213 D net205 VPW N12LL W=350.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=290.00n L=60.00n
MM39 QN OS VSS VPW N12LL W=430.00n L=60.00n
MM62 OS c net181 VPW N12LL W=400.00n L=60.00n
MM63 net181 S VSS VPW N12LL W=400.00n L=60.00n
MM61 M cn net193 VPW N12LL W=260.00n L=60.00n
MM58 SEN SE VSS VPW N12LL W=290.00n L=60.00n
MM70 net205 SN net0172 VPW N12LL W=350.00n L=60.00n
MM60 net193 net0370 VSS VPW N12LL W=260.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net172 cn OS VPW N12LL W=200.00n L=60.00n
MM23 VSS NET64 net172 VPW N12LL W=200.00n L=60.00n
MM69 net213 SNN net0172 VPW N12LL W=300.00n L=60.00n
MM19 Q NET64 VSS VPW N12LL W=430.00n L=60.00n
MM17 NET64 OS VSS VPW N12LL W=300.00n L=60.00n
MM12 net240 c M VPW N12LL W=200.00n L=60.00n
MM11 VSS S net240 VPW N12LL W=200.00n L=60.00n
MM0 S M VSS VPW N12LL W=360.00n L=60.00n
MM66 net0418 SNN net296 VNW P12LL W=590.00n L=60.00n
MM50 net288 SI VDD VNW P12LL W=410.00n L=60.00n
MM51 net0370 SEN net288 VNW P12LL W=410.00n L=60.00n
MM52 net296 D VDD VNW P12LL W=590.00n L=60.00n
MM53 net0370 SE net0418 VNW P12LL W=590.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=440.00n L=60.00n
MM40 QN OS VDD VNW P12LL W=650.00n L=60.00n
MM64 net268 S VDD VNW P12LL W=480.00n L=60.00n
MM65 OS cn net268 VNW P12LL W=480.00n L=60.00n
MM67 net0418 RN VDD VNW P12LL W=400.00n L=60.00n
MM59 SEN SE VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD NET64 net253 VNW P12LL W=300.00n L=60.00n
MM25 net253 c OS VNW P12LL W=300.00n L=60.00n
MM20 Q NET64 VDD VNW P12LL W=650.00n L=60.00n
MM18 NET64 OS VDD VNW P12LL W=450.00n L=60.00n
MM14 net313 cn M VNW P12LL W=300.00n L=60.00n
MM13 VDD S net313 VNW P12LL W=300.00n L=60.00n
MM55 net280 net0370 VDD VNW P12LL W=390.00n L=60.00n
MM56 M c net280 VNW P12LL W=390.00n L=60.00n
MM1 S M VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRSNHSV2
****Sub-Circuit for SDGRSNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRSNHSV4 CK D Q QN RN SE SI SN VDD VSS
MM45 net0370 SE net201 VPW N12LL W=300.00n L=60.00n
MM46 net201 SI VSS VPW N12LL W=300.00n L=60.00n
MM47 net0172 RN VSS VPW N12LL W=350.00n L=60.00n
MM48 net0370 SEN net213 VPW N12LL W=350.00n L=60.00n
MM49 net213 D net205 VPW N12LL W=350.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=290.00n L=60.00n
MM39 QN OS VSS VPW N12LL W=860.00n L=60.00n
MM62 OS c net181 VPW N12LL W=450.00n L=60.00n
MM63 net181 S VSS VPW N12LL W=450.00n L=60.00n
MM61 M cn net193 VPW N12LL W=260.00n L=60.00n
MM58 SEN SE VSS VPW N12LL W=290.00n L=60.00n
MM70 net205 SN net0172 VPW N12LL W=350.00n L=60.00n
MM60 net193 net0370 VSS VPW N12LL W=260.00n L=60.00n
MM30 c cn VSS VPW N12LL W=260.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net172 cn OS VPW N12LL W=200.00n L=60.00n
MM23 VSS NET64 net172 VPW N12LL W=200.00n L=60.00n
MM69 net213 SNN net0172 VPW N12LL W=300.00n L=60.00n
MM19 Q NET64 VSS VPW N12LL W=860.00n L=60.00n
MM17 NET64 OS VSS VPW N12LL W=360.00n L=60.00n
MM12 net240 c M VPW N12LL W=200.00n L=60.00n
MM11 VSS S net240 VPW N12LL W=200.00n L=60.00n
MM0 S M VSS VPW N12LL W=360.00n L=60.00n
MM66 net0418 SNN net296 VNW P12LL W=590.00n L=60.00n
MM50 net288 SI VDD VNW P12LL W=450.00n L=60.00n
MM51 net0370 SEN net288 VNW P12LL W=450.00n L=60.00n
MM52 net296 D VDD VNW P12LL W=590.00n L=60.00n
MM53 net0370 SE net0418 VNW P12LL W=590.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=440.00n L=60.00n
MM40 QN OS VDD VNW P12LL W=1.3u L=60.00n
MM64 net268 S VDD VNW P12LL W=570.00n L=60.00n
MM65 OS cn net268 VNW P12LL W=570.00n L=60.00n
MM67 net0418 RN VDD VNW P12LL W=400.00n L=60.00n
MM59 SEN SE VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=390.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD NET64 net253 VNW P12LL W=300.00n L=60.00n
MM25 net253 c OS VNW P12LL W=300.00n L=60.00n
MM20 Q NET64 VDD VNW P12LL W=1.3u L=60.00n
MM18 NET64 OS VDD VNW P12LL W=540.00n L=60.00n
MM14 net313 cn M VNW P12LL W=300.00n L=60.00n
MM13 VDD S net313 VNW P12LL W=300.00n L=60.00n
MM55 net280 net0370 VDD VNW P12LL W=390.00n L=60.00n
MM56 M c net280 VNW P12LL W=390.00n L=60.00n
MM1 S M VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRSNHSV4
****Sub-Circuit for SDGSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGSNHSV1 CK D Q QN SE SI SN VDD VSS
MM39 QN PS VSS VPW N12LL W=290.00n L=60.00n
MM45 N74 SE net0128 VPW N12LL W=200.00n L=60.00n
MM46 net0128 SI VSS VPW N12LL W=200.00n L=60.00n
MM48 N74 cn PM VPW N12LL W=270.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=200.00n L=60.00n
MM52 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM3 M c PS VPW N12LL W=270.00n L=60.00n
MM42 net69 SNN VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=250.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn PS VPW N12LL W=200.00n L=60.00n
MM23 VSS S net48 VPW N12LL W=200.00n L=60.00n
MM19 Q S VSS VPW N12LL W=290.00n L=60.00n
MM17 S PS VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c PM VPW N12LL W=200.00n L=60.00n
MM11 VSS M net52 VPW N12LL W=200.00n L=60.00n
MM9 N74 SEN net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=250.00n L=60.00n
MM0 M PM VSS VPW N12LL W=270.00n L=60.00n
MM41 net_0231 SNN VDD VNW P12LL W=400.00n L=60.00n
MM40 QN PS VDD VNW P12LL W=440.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=300.00n L=60.00n
MM50 net0207 SI VDD VNW P12LL W=300.00n L=60.00n
MM51 N74 SEN net0207 VNW P12LL W=300.00n L=60.00n
MM54 N74 c PM VNW P12LL W=400.00n L=60.00n
MM4 M cn PS VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=380.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD S net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c PS VNW P12LL W=300.00n L=60.00n
MM20 Q S VDD VNW P12LL W=440.00n L=60.00n
MM18 S PS VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn PM VNW P12LL W=300.00n L=60.00n
MM13 VDD M net117 VNW P12LL W=300.00n L=60.00n
MM10 N74 SE net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=400.00n L=60.00n
MM56 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM1 M PM VDD VNW P12LL W=400.00n L=60.00n
.ENDS SDGSNHSV1
****Sub-Circuit for SDGSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGSNHSV2 CK D Q QN SE SI SN VDD VSS
MM39 QN PS VSS VPW N12LL W=430.00n L=60.00n
MM45 N74 SE net0128 VPW N12LL W=200.00n L=60.00n
MM46 net0128 SI VSS VPW N12LL W=200.00n L=60.00n
MM48 N74 cn PM VPW N12LL W=360.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=200.00n L=60.00n
MM52 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM3 M c PS VPW N12LL W=390.00n L=60.00n
MM42 net69 SNN VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=380.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn PS VPW N12LL W=200.00n L=60.00n
MM23 VSS S net48 VPW N12LL W=200.00n L=60.00n
MM19 Q S VSS VPW N12LL W=430.00n L=60.00n
MM17 S PS VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c PM VPW N12LL W=200.00n L=60.00n
MM11 VSS M net52 VPW N12LL W=200.00n L=60.00n
MM9 N74 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 M PM VSS VPW N12LL W=390.00n L=60.00n
MM41 net_0231 SNN VDD VNW P12LL W=600.0n L=60.00n
MM40 QN PS VDD VNW P12LL W=650.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=300.00n L=60.00n
MM50 net0207 SI VDD VNW P12LL W=300.00n L=60.00n
MM51 N74 SEN net0207 VNW P12LL W=300.00n L=60.00n
MM54 N74 c PM VNW P12LL W=540.00n L=60.00n
MM4 M cn PS VNW P12LL W=580.00n L=60.00n
MM29 c cn VDD VNW P12LL W=570.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD S net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c PS VNW P12LL W=300.00n L=60.00n
MM20 Q S VDD VNW P12LL W=650.00n L=60.00n
MM18 S PS VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn PM VNW P12LL W=300.00n L=60.00n
MM13 VDD M net117 VNW P12LL W=300.00n L=60.00n
MM10 N74 SE net128 VNW P12LL W=600.0n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=600.0n L=60.00n
MM56 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM1 M PM VDD VNW P12LL W=580.00n L=60.00n
.ENDS SDGSNHSV2
****Sub-Circuit for SDGSNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGSNHSV4 CK D Q QN SE SI SN VDD VSS
MM39 QN PS VSS VPW N12LL W=860.00n L=60.00n
MM45 N74 SE net0128 VPW N12LL W=200.00n L=60.00n
MM46 net0128 SI VSS VPW N12LL W=200.00n L=60.00n
MM48 N74 cn PM VPW N12LL W=400.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=200.00n L=60.00n
MM52 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM3 M c PS VPW N12LL W=430.00n L=60.00n
MM42 net69 SNN VSS VPW N12LL W=250.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn PS VPW N12LL W=200.00n L=60.00n
MM23 VSS S net48 VPW N12LL W=200.00n L=60.00n
MM19 Q S VSS VPW N12LL W=860.00n L=60.00n
MM17 S PS VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c PM VPW N12LL W=200.00n L=60.00n
MM11 VSS M net52 VPW N12LL W=200.00n L=60.00n
MM9 N74 SEN net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 M PM VSS VPW N12LL W=430.00n L=60.00n
MM41 net_0231 SNN VDD VNW P12LL W=650.00n L=60.00n
MM40 QN PS VDD VNW P12LL W=1.3u L=60.00n
MM44 SNN SN VDD VNW P12LL W=300.00n L=60.00n
MM50 net0207 SI VDD VNW P12LL W=300.00n L=60.00n
MM51 N74 SEN net0207 VNW P12LL W=300.00n L=60.00n
MM54 N74 c PM VNW P12LL W=600.0n L=60.00n
MM4 M cn PS VNW P12LL W=650.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD S net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c PS VNW P12LL W=300.00n L=60.00n
MM20 Q S VDD VNW P12LL W=1.3u L=60.00n
MM18 S PS VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn PM VNW P12LL W=300.00n L=60.00n
MM13 VDD M net117 VNW P12LL W=300.00n L=60.00n
MM10 N74 SE net128 VNW P12LL W=650.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=650.00n L=60.00n
MM56 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM1 M PM VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDGSNHSV4
****Sub-Circuit for SDHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDHSV1 CK D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=290.00n L=60.00n
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=280.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=280.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=290.00n L=60.00n
MM53 QN s VDD VNW P12LL W=440.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=300.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=300.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDHSV1
****Sub-Circuit for SDHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDHSV2 CK D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=430.00n L=60.00n
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=400.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=400.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM53 QN s VDD VNW P12LL W=650.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDHSV2
****Sub-Circuit for SDHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDHSV4 CK D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=860.00n L=60.00n
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=420.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=300.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=300.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM53 QN s VDD VNW P12LL W=1.3u L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=520.0n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=520.0n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.0n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDHSV4
****Sub-Circuit for SDQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDQHSV1 CK D Q SE SI VDD VSS
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=280.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=280.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=290.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=300.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=300.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDQHSV1
****Sub-Circuit for SDQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDQHSV2 CK D Q SE SI VDD VSS
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=400.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=400.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDQHSV2
****Sub-Circuit for SDQHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SDQHSV4 CK D Q SE SI VDD VSS
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=430.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=300.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=300.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=490.0n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=490.0n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.0n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDQHSV4
****Sub-Circuit for SDRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNHSV1 CK D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=290.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=290.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=290.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=290.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=440.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=330.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=330.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=330.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDRNHSV1
****Sub-Circuit for SDRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNHSV2 CK D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=430.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=320.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=320.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=650.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=350.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=350.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=350.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNHSV2
****Sub-Circuit for SDRNHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SDRNHSV4 CK D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=430.00n L=60.00n m=2
MM45 net_0137 sen net_0133 VPW N12LL W=430.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=400.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=300.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=300.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=650.00n L=60.00n m=2
MM47 net_0137 SE net_0212 VNW P12LL W=500n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=450.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=500n L=60.00n
MM8 net128 SI VDD VNW P12LL W=500n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNHSV4
****Sub-Circuit for SDRNQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNQHSV1 CK D Q RDN SE SI VDD VSS
MM45 net_0137 sen net_0133 VPW N12LL W=290.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=290.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=290.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=330.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=330.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=330.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDRNQHSV1
****Sub-Circuit for SDRNQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNQHSV2 CK D Q RDN SE SI VDD VSS
MM45 net_0137 sen net_0133 VPW N12LL W=320.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=320.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=350.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=350.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=350.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNQHSV2
****Sub-Circuit for SDRNQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNQHSV4 CK D Q RDN SE SI VDD VSS
MM45 net_0137 sen net_0133 VPW N12LL W=430.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=400.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=300.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=300.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=500n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=450.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=500n L=60.00n
MM8 net128 SI VDD VNW P12LL W=500n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNQHSV4
****Sub-Circuit for SDRSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRSNHSV1 CK D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=250.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=290.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=200.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=260.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=260.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=260.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=260.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=280.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=330.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=420.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=380.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=330.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=330.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=330.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=440.00n L=60.00n
.ENDS SDRSNHSV1
****Sub-Circuit for SDRSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRSNHSV2 CK D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=280.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=250.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=360.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=390.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=200.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=220.00n L=60.00n
MM40 net43 R L VPW N12LL W=280.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=220.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=220.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=220.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=380.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=300.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=300.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=600.00n L=60.00n
.ENDS SDRSNHSV2
****Sub-Circuit for SDRSNHSV4, Mon May 30 16:10:14 CST 2011****
.SUBCKT SDRSNHSV4 CK D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=280.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=250.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=320.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=430.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=400.00n L=60.00n
MM40 net43 R L VPW N12LL W=280.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=400.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=400.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=500.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM57 net_0140 c net_0139 VNW P12LL W=580.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=600.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=520.00n L=60.00n
MM29 c cn VDD VNW P12LL W=620.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=380.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=500.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=500.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=500.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=650.00n L=60.00n
.ENDS SDRSNHSV4
****Sub-Circuit for SDSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDSNHSV1 CK D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=300.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=300.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=200.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=400.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=400.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=300.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=450.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=450.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=400.00n L=60.00n
.ENDS SDSNHSV1
****Sub-Circuit for SDSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDSNHSV2 CK D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=300.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=300.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=200.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=420.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=420.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=300.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=450.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=450.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=390.00n L=60.00n
.ENDS SDSNHSV2
****Sub-Circuit for SDSNHSV4, Mon May 30 17:13:17 CST 2011****
.SUBCKT SDSNHSV4 CK D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=300.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=300.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=200.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=360.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=300.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=450.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=450.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM38 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=625.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=480.00n L=60.00n
.ENDS SDSNHSV4
****Sub-Circuit for SDXHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDXHSV1 CK DA DB Q QN SA SE SI VDD VSS
MM5 net41 SB net_0171 VPW N12LL W=240.00n L=60.00n
MM49 net39 DA VSS VPW N12LL W=350.00n L=60.00n
MM48 net39 SA net_0171 VPW N12LL W=240.00n L=60.00n
MM37 SEN SE VSS VPW N12LL W=240.00n L=60.00n
MM41 net41 DB VSS VPW N12LL W=350.00n L=60.00n
MM31 SB SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=350.00n L=60.00n
MM19 QN s VSS VPW N12LL W=350.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM7 m c net43 VPW N12LL W=350.00n L=60.00n
MM12 net52 c net_0157 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM46 net_0169 SE VSS VPW N12LL W=240.00n L=60.00n
MM45 net_0153 sin net_0169 VPW N12LL W=240.00n L=60.00n
MM43 net_0161 SEN VSS VPW N12LL W=300.00n L=60.00n
MM9 net_0157 cn net_0153 VPW N12LL W=300.00n L=60.00n
MM42 net_0153 net_0171 net_0161 VPW N12LL W=300.00n L=60.00n
MM6 sin SI VSS VPW N12LL W=350.00n L=60.00n
MM0 m net_0157 VSS VPW N12LL W=350.00n L=60.00n
MM52 net39 DA VDD VNW P12LL W=440.0n L=60.00n
MM53 sin SI VDD VNW P12LL W=440.0n L=60.00n
MM54 net41 SA net_0171 VNW P12LL W=300.0n L=60.00n
MM55 net41 DB VDD VNW P12LL W=440.0n L=60.00n
MM56 net39 SB net_0171 VNW P12LL W=300.0n L=60.00n
MM38 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM4 m cn net43 VNW P12LL W=440.0n L=60.00n
MM44 net_0236 SE VDD VNW P12LL W=450.00n L=60.00n
MM32 SB SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM20 QN s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM47 net_0233 net_0171 net_0236 VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0157 VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM51 net_0233 sin net_0252 VNW P12LL W=300.00n L=60.00n
MM50 net_0252 SEN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0157 c net_0233 VNW P12LL W=450.00n L=60.00n
MM1 m net_0157 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDXHSV1
****Sub-Circuit for SDXHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDXHSV2 CK DA DB Q QN SA SE SI VDD VSS
MM8 sin SI VSS VPW N12LL W=350.00n L=60.00n
MM41 net41 DB VSS VPW N12LL W=430.00n L=60.00n
MM37 SEN SE VSS VPW N12LL W=240.00n L=60.00n
MM31 SB SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM19 QN s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM2 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0157 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM46 net_0169 SE VSS VPW N12LL W=240.00n L=60.00n
MM45 net_0153 sin net_0169 VPW N12LL W=240.00n L=60.00n
MM43 net_0161 SEN VSS VPW N12LL W=350.00n L=60.00n
MM9 net_0157 cn net_0153 VPW N12LL W=350.00n L=60.00n
MM42 net_0153 net_0152 net_0161 VPW N12LL W=350.00n L=60.00n
MM48 net39 SA net_0152 VPW N12LL W=240.00n L=60.00n
MM5 net41 SB net_0152 VPW N12LL W=240.00n L=60.00n
MM49 net39 DA VSS VPW N12LL W=430.00n L=60.00n
MM0 m net_0157 VSS VPW N12LL W=430.00n L=60.00n
MM38 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM53 sin SI VDD VNW P12LL W=440.0n L=60.00n
MM44 net_0236 SE VDD VNW P12LL W=440.00n L=60.00n
MM32 SB SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=550.00n L=60.00n
MM20 QN s VDD VNW P12LL W=550.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM7 m cn net43 VNW P12LL W=540.00n L=60.00n
MM47 net_0233 net_0152 net_0236 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0157 VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM51 net_0233 sin net_0252 VNW P12LL W=300.00n L=60.00n
MM50 net_0252 SEN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0157 c net_0233 VNW P12LL W=440.00n L=60.00n
MM56 net39 SB net_0152 VNW P12LL W=300.0n L=60.00n
MM54 net41 SA net_0152 VNW P12LL W=300.0n L=60.00n
MM55 net41 DB VDD VNW P12LL W=550.0n L=60.00n
MM52 net39 DA VDD VNW P12LL W=550.0n L=60.00n
MM1 m net_0157 VDD VNW P12LL W=550.00n L=60.00n
.ENDS SDXHSV2
****Sub-Circuit for SDXHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDXHSV4 CK DA DB Q QN SA SE SI VDD VSS
MM8 sin SI VSS VPW N12LL W=350.00n L=60.00n
MM41 net41 DB VSS VPW N12LL W=430.00n L=60.00n
MM37 SEN SE VSS VPW N12LL W=240.00n L=60.00n
MM31 SB SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM19 QN s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM2 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0157 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM46 net_0169 SE VSS VPW N12LL W=240.00n L=60.00n
MM45 net_0153 sin net_0169 VPW N12LL W=240.00n L=60.00n
MM43 net_0161 SEN VSS VPW N12LL W=350.00n L=60.00n
MM9 net_0157 cn net_0153 VPW N12LL W=350.00n L=60.00n
MM42 net_0153 net_0152 net_0161 VPW N12LL W=350.00n L=60.00n
MM49 net39 DA VSS VPW N12LL W=430.00n L=60.00n
MM5 net41 SB net_0152 VPW N12LL W=240.00n L=60.00n
MM48 net39 SA net_0152 VPW N12LL W=240.00n L=60.00n
MM0 m net_0157 VSS VPW N12LL W=430.00n L=60.00n
MM38 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0236 SE VDD VNW P12LL W=440.00n L=60.00n
MM56 net39 SB net_0152 VNW P12LL W=300.0n L=60.00n
MM54 net41 SA net_0152 VNW P12LL W=300.0n L=60.00n
MM52 net39 DA VDD VNW P12LL W=550.0n L=60.00n
MM55 net41 DB VDD VNW P12LL W=550.0n L=60.00n
MM32 SB SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.1u L=60.00n
MM20 QN s VDD VNW P12LL W=1.1u L=60.00n
MM18 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM53 sin SI VDD VNW P12LL W=440.0n L=60.00n
MM7 m cn net43 VNW P12LL W=540.00n L=60.00n
MM47 net_0233 net_0152 net_0236 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0157 VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM51 net_0233 sin net_0252 VNW P12LL W=300.00n L=60.00n
MM50 net_0252 SEN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0157 c net_0233 VNW P12LL W=440.00n L=60.00n
MM1 m net_0157 VDD VNW P12LL W=550.00n L=60.00n
.ENDS SDXHSV4
****Sub-Circuit for SEDGRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNHSV1 CK D E Q QN RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM64 QN s VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=290.00n L=60.00n
MM17 sp s VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM65 QN s VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=440.00n L=60.00n
MM18 sp s VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNHSV1
****Sub-Circuit for SEDGRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNHSV2 CK D E Q QN RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM64 QN s VSS VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=430.00n L=60.00n
MM17 sp s VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM65 QN s VDD VNW P12LL W=650.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=650.00n L=60.00n
MM18 sp s VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNHSV2
****Sub-Circuit for SEDGRNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNHSV4 CK D E Q QN RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM64 QN s VSS VPW N12LL W=860.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=860.00n L=60.00n
MM17 sp s VSS VPW N12LL W=400.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM65 QN s VDD VNW P12LL W=1.3u L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=1.3u L=60.00n
MM18 sp s VDD VNW P12LL W=480.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNHSV4
****Sub-Circuit for SEDGRNQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNQHSV1 CK D E Q RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=290.00n L=60.00n
MM17 sp s VSS VPW N12LL W=220.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=440.00n L=60.00n
MM18 sp s VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNQHSV1
****Sub-Circuit for SEDGRNQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNQHSV2 CK D E Q RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=430.00n L=60.00n
MM17 sp s VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=650.00n L=60.00n
MM18 sp s VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNQHSV2
****Sub-Circuit for SEDGRNQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNQHSV4 CK D E Q RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=860.00n L=60.00n
MM17 sp s VSS VPW N12LL W=310.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=1.3u L=60.00n
MM18 sp s VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNQHSV4
****Sub-Circuit for SEDHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDHSV1 CK D E Q QN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=300.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=300.00n L=60.00n
MM68 QN s VSS VPW N12LL W=290.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=420.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=420.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=420.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=420.00n L=60.00n
MM0 m pm VSS VPW N12LL W=400.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=300.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=300.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM69 QN s VDD VNW P12LL W=440.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=600.00n L=60.00n
.ENDS SEDHSV1
****Sub-Circuit for SEDHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDHSV2 CK D E Q QN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 QN s VSS VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=400.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=400.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM69 QN s VDD VNW P12LL W=650.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDHSV2
****Sub-Circuit for SEDHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDHSV4 CK D E Q QN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 QN s VSS VPW N12LL W=860.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=390.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=440.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=440.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM69 QN s VDD VNW P12LL W=1.3u L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDHSV4
****Sub-Circuit for SEDQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDQHSV1 CK D E Q SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=300.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=300.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=300.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=300.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDQHSV1
****Sub-Circuit for SEDQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDQHSV2 CK D E Q SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=400.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=400.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDQHSV2
****Sub-Circuit for SEDQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDQHSV4 CK D E Q SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=420.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=420.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDQHSV4
****Sub-Circuit for SEDRNHSV1, Fri May 27 10:36:55 CST 2011****
.SUBCKT SEDRNHSV1 CK D E Q QN RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=390.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM73 QN s VSS VPW N12LL W=290.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=250.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=250.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=275.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=250.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=270.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM74 QN s VDD VNW P12LL W=440.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=355.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=390.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=390.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=380.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=400.00n L=60.00n
.ENDS SEDRNHSV1
****Sub-Circuit for SEDRNHSV2, Thu May 26 17:37:04 CST 2011****
.SUBCKT SEDRNHSV2 CK D E Q QN RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=390.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM73 QN s VSS VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=250.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=250.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=275.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM74 QN s VDD VNW P12LL W=650.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=355.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=390.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=390.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SEDRNHSV2
****Sub-Circuit for SEDRNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDRNHSV4 CK D E Q QN RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=360.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=360.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM73 QN s VSS VPW N12LL W=860.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=250.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=250.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=275.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=400.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=400.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=470.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=470.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM74 QN s VDD VNW P12LL W=1.3u L=60.00n
MM53 net0267 SE VDD VNW P12LL W=355.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=390.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=390.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=600.00n L=60.00n
.ENDS SEDRNHSV4
****Sub-Circuit for SEDRNQHSV1, Thu May 26 14:31:08 CST 2011****
.SUBCKT SEDRNQHSV1 CK D E Q RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=390.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=240.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=240.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=300.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=385.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=385.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=370.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=380.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=380.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDRNQHSV1
****Sub-Circuit for SEDRNQHSV2, Thu May 26 13:48:52 CST 2011****
.SUBCKT SEDRNQHSV2 CK D E Q RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=240.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=240.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=290.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=380.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=380.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=380.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDRNQHSV2
****Sub-Circuit for SEDRNQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDRNQHSV4 CK D E Q RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=240.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=240.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=300.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=390.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=380.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=380.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDRNQHSV4
****Sub-Circuit for SNDHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDHSV1 CKN D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=290.00n L=60.00n
MM46 net_0107 SE VSS VPW N12LL W=250.00n L=60.00n
MM45 net_0163 SI net_0107 VPW N12LL W=250.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=230.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=230.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=250.00n L=60.00n
MM30 cn c VSS VPW N12LL W=250.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=250.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=250.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=270.00n L=60.00n
MM53 QN s VDD VNW P12LL W=440.00n L=60.00n
MM51 net128 SI net_0174 VNW P12LL W=650.00n L=60.00n
MM50 net_0174 SEN VDD VNW P12LL W=650.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=380.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=650.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=650.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=650.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=400.00n L=60.00n
.ENDS SNDHSV1
****Sub-Circuit for SNDHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDHSV2 CKN D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=430.00n L=60.00n
MM46 net_0107 SE VSS VPW N12LL W=250.00n L=60.00n
MM45 net_0163 SI net_0107 VPW N12LL W=250.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=230.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=230.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=250.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=250.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=250.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=390.00n L=60.00n
MM53 QN s VDD VNW P12LL W=650.00n L=60.00n
MM51 net128 SI net_0174 VNW P12LL W=650.00n L=60.00n
MM50 net_0174 SEN VDD VNW P12LL W=650.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=650.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=650.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=650.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=580.00n L=60.00n
.ENDS SNDHSV2
****Sub-Circuit for SNDHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDHSV4 CKN D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=860.00n L=60.00n
MM46 net_0107 SE VSS VPW N12LL W=260.00n L=60.00n
MM45 net_0163 SI net_0107 VPW N12LL W=260.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=250.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=250.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=260.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=260.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=260.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM53 QN s VDD VNW P12LL W=1.3u L=60.00n
MM51 net128 SI net_0174 VNW P12LL W=650.00n L=60.00n
MM50 net_0174 SEN VDD VNW P12LL W=650.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=650.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=650.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=650.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SNDHSV4
****Sub-Circuit for SNDRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRNHSV1 CKN D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=290.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=300.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=300.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=300.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=300.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=300.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM39 s ps net_099 VPW N12LL W=360.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=360.00n L=60.00n
MM30 cn c VSS VPW N12LL W=300.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=300.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=440.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=500.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM38 s ps VDD VNW P12LL W=390.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=390.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=450.00n L=60.00n
MM29 cn c VDD VNW P12LL W=450.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=450.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=450.00n L=60.00n
.ENDS SNDRNHSV1
****Sub-Circuit for SNDRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRNHSV2 CKN D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=430.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=350.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=350.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=300.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=290.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=300.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=190.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM39 s ps net_099 VPW N12LL W=360.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=360.00n L=60.00n
MM30 cn c VSS VPW N12LL W=300.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=190.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=190.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=300.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=650.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=450.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=450.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM38 s ps VDD VNW P12LL W=390.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=390.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=445.00n L=60.00n
MM29 cn c VDD VNW P12LL W=450.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=450.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=450.00n L=60.00n
.ENDS SNDRNHSV2
****Sub-Circuit for SNDRNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRNHSV4 CKN D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=860.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=350.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=350.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=300.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=300.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=300.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM39 s ps net_099 VPW N12LL W=380.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=380.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=300.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=1.3u L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=500.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM38 s ps VDD VNW P12LL W=350.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=450.00n L=60.00n
MM29 cn c VDD VNW P12LL W=530.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn ps VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=450.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=450.00n L=60.00n
.ENDS SNDRNHSV4
****Sub-Circuit for SNDRSNHSV1, Mon May 30 19:16:43 CST 2011****
.SUBCKT SNDRSNHSV1 CKN D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=270.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=340.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=300.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=300.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=300.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=300.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=450.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=450.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=500.00n L=60.00n
MM29 cn c VDD VNW P12LL W=540.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=540.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=540.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=500.00n L=60.00n
.ENDS SNDRSNHSV1
****Sub-Circuit for SNDRSNHSV2, Mon May 30 17:13:17 CST 2011****
.SUBCKT SNDRSNHSV2 CKN D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=270.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=340.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=300.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=300.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=300.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=300.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=450.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=450.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=500.00n L=60.00n
MM29 cn c VDD VNW P12LL W=540.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=540.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=540.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=500.00n L=60.00n
.ENDS SNDRSNHSV2
****Sub-Circuit for SNDRSNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRSNHSV4 CKN D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=270.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=350.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=360.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=300.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=320.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=320.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=300.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=450.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=450.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=540.00n L=60.00n
MM29 cn c VDD VNW P12LL W=540.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=540.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=540.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=540.00n L=60.00n
.ENDS SNDRSNHSV4
****Sub-Circuit for SNDSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDSNHSV1 CKN D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=220.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=220.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=220.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=220.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=200.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=250.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=220.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=430.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=480.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=480.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=480.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=480.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=380.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=480.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=500.00n L=60.00n
.ENDS SNDSNHSV1
****Sub-Circuit for SNDSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDSNHSV2 CKN D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=220.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=220.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=220.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=220.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=250.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=220.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=430.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=480.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=480.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=480.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=480.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=480.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=500.00n L=60.00n
.ENDS SNDSNHSV2
****Sub-Circuit for SNDSNHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SNDSNHSV4 CKN D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=250.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=250.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=250.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=250.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=390.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=250.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=430.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=480.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=480.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=480.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=480.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM38 s net43 VDD VNW P12LL W=540.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=470.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=480.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=500.00n L=60.00n
.ENDS SNDSNHSV4
