//* No part of this file can be released without the consent of SMIC.
//*
//* Note: SMIC recommends that users use version 6.1.0 08/15/2006 15:48 (usimlx111), or version 6.2.0 09/04/2007 08:19 (usimlx110),
//* or Spectre 7.01ISR20 , or Spectre 7.1ISR6 , or Spectre version after 7.1ISR6. And please do not use Spectre version 6.2.1 32bit 05/29/2008 05:19 (sfrh56)  
//* until  the version before 7.01ISR20 to run simulation, because the mutual coupling coefficient K will be restricted to [-1,1] within these versions.
//* Note: SMIC recommends that users set options reltol=1e-2 if circuit is not convergence.
//******************************************************************************************
//* 0.11um Mixed Signal 1P8M with MIM Salicide 1.2V/3.3V RF SPICE Model (for SPECTRE only) *
//******************************************************************************************
//*
//* Release version    : 1.14
//*
//* Release date       : 03/30/2016
//*
//* Simulation tool    : Cadence spectre V6.0
//*
//*
//*  Inductor   :
//* *  *-----------------*-------------------------*-------------------------*-------------------------*-------------------------*
//*    |  Turn & Radius  |   Turn=1,rin=50~120um   |   Turn=2,rin=50~120um   |   Turn=3,rin=50~120um   |   Turn=4,rin=50~120um   |
//     *-------------------------------------------*-------------------------*-------------------------*-------------------------*
//*    |     Model Name  |   rf_3Tdiff_1talpa_t1   |   rf_3Tdiff_1talpa_t2   |   rf_3Tdiff_1talpa_t3   |   rf_3Tdiff_1talpa_t4   |
//*    *-----------------*-------------------------*-------------------------*-------------------------*-------------------------*
//*    |  Turn & Radius  |   Turn=5,rin=50~120um   |   Turn=6,rin=50~120um   |   Turn=7,rin=50~120um   |                          
//     *-------------------------------------------*-------------------------*-------------------------*                          
//*    |     Model Name  |   rf_3Tdiff_1talpa_t5   |   rf_3Tdiff_1talpa_t6   |   rf_3Tdiff_1talpa_t7   |                          
//*    *-----------------*-------------------------*-------------------------*-------------------------*                          
//*Temperature range: -40~125 Celsius Degree
//
//*** 0.11um Three Port Differential Inductor 
simulator lang=spectre  insensitive=yes
//*********************************************** 
subckt rf_3Tdiff_1talpa_t1 (PLUS MINUS CT)
// ***********************************************************************************
//***PLUS=port1, MINUS=port2**//
//***0.11um 1 turns 3-T differential inductor scalable model**//
//***R= inner radius; N=turns; W=width; S=spacing**//
//***In this model, R is scalalbe, N=1, S=2.0um, W=15um**//
// ***********************************************************************************
parameters R=50.0e-6 N=1 
+Ldc1=3.4052e-6*R-2.969e-11                    
+Rdc1=1948.3*R+0.037897                        
+Ldc2=Ldc1                                     
+Rdc2=Rdc1                                     
+Cox1=2e-10*R+1e-14                            
+Csub1=6e-15                                   
+Rsub1=700                                     
+Cox2=Cox1                                     
+Csub2=Csub1                                   
+Rsub2=Rsub1                                   
+Cf=1.25e-10*R+2.5e-16                         
+mm=0.55                                       
+Lsshort=7.7302e-11*exp(6886.7*R)              
+Rsshort=0.21                                  
+Krssk=5                                       
+Klssk=1                                       
+Krp=46.946*pwr(R,0.50372)                     
+Klp=0.22                                      
+Ls1=1/(1+Klp/pwr(1+Krp,2))*Ldc1/2             
+Ls2=1/(1+Klp/pwr(1+Krp,2))*Ldc2/2             
+Rs1=(1+1/Krp)*Rdc1/2                          
+Rs2=(1+1/Krp)*Rdc2/2                          
+Rp1=Krp*Rs1                                   
+Rp2=Krp*Rs2                                   
+Lp1=Klp*Ls1                                   
+Lp2=Klp*Ls2                                   
+Lshort=Lsshort                                
+Lssk=Lsshort*Klssk                            
+Rshort=Rsshort                                
+Rssk=Rsshort*Krssk                            

//***equivalent circuit

Cf_Ind     (PLUS  MINUS) capacitor c=Cf
Ls1_Ind    (12  23) inductor l=Ls1*(1+dls_3Tdiff_1talpa)
Rs1_Ind    (PLUS 12) resistor r=Rs1*(1+drs_3Tdiff_1talpa) tc1=0.003
Ls2_Ind    (23  34) inductor l=Ls2*(1+dls_3Tdiff_1talpa)
Rs2_Ind    (34 MINUS) resistor r=Rs2*(1+drs_3Tdiff_1talpa) tc1=0.003
Lp1_Ind    (56 12) inductor l=Lp1
Rp1_Ind    (PLUS 56) resistor r=Rp1 tc1=0.003
Lp2_Ind    (78 MINUS) inductor l=Lp2
Rp2_Ind    (34 78) resistor r=Rp2 tc1=0.003
Cox1_Ind   (PLUS  11) capacitor c=Cox1
Rsub1_Ind  (11  0) resistor r=Rsub1
Csub1_Ind  (11  0) capacitor c=Csub1
Cox2_Ind   (MINUS  22) capacitor c=Cox2
Rsub2_Ind  (22  0) resistor r=Rsub2
Csub2_Ind  (22  0) capacitor c=Csub2
Lshort_Ind   (23  31) inductor l=Lshort
Rshort_Ind  (31  CT) resistor r=Rshort*(1+drs_3Tdiff_1talpa) tc1=0.003
Rssk_Ind  (31  32) resistor r=Rssk tc1=0.003  
Lssk_Ind  (32  CT) inductor l=Lssk  
Klm1      mutual_inductor coupling=mm ind1=Ls1_Ind ind2=Ls2_Ind

ends rf_3Tdiff_1talpa_t1

subckt rf_3Tdiff_1talpa_t2 (PLUS MINUS CT)
// ***********************************************************************************
//***PLUS=port1, MINUS=port2**//
//***0.11um 2 turns 3-T differential inductor scalable model**//
//***R= inner radius; N=turns; W=width; S=spacing**//
//***In this model, R is scalalbe, N=2, S=2.0um, W=15um**//
// ***********************************************************************************
parameters R=50.0e-6 N=2 
+Ldc1=1.2664e-5*R-1.0517e-10
+Rdc1=3879.3*R+0.20276 
+Ldc2=Ldc1
+Rdc2=4000*R+0.08 
+Cox1=6e-14
+Csub1=4.5e-10*R+1.75e-14
+Rsub1=650
+Cox2=Cox1
+Csub2=Csub1
+Rsub2=Rsub1 
+Cf=4.0172e-10*R+1.0345E-16
+mm=0.45
+Lsshort=8.0343e-11*log(R)+9.3491e-10
+Rsshort=7827.6*R+0.34466
+Krssk=5 
+Klssk=0.5 
+Krp=14.916*pwr(R,0.36985) 
+Klp=0.0019321*pwr(R,-0.50312) 
+Ls1=1/(1+Klp/pwr(1+Krp,2))*Ldc1/2
+Ls2=1/(1+Klp/pwr(1+Krp,2))*Ldc2/2
+Rs1=(1+1/Krp)*Rdc1/2
+Rs2=(1+1/Krp)*Rdc2/2
+Rp1=Krp*Rs1
+Rp2=Krp*Rs2
+Lp1=Klp*Ls1
+Lp2=Klp*Ls2
+Lshort=Lsshort
+Lssk=Lsshort*Klssk
+Rshort=Rsshort
+Rssk=Rsshort*Krssk
//***equivalent circuit
Cf_Ind     (PLUS  MINUS) capacitor c=Cf
Ls1_Ind    (12  23) inductor l=Ls1*(1+dls_3Tdiff_1talpa)
Rs1_Ind    (PLUS 12) resistor r=Rs1*(1+drs_3Tdiff_1talpa) tc1=0.003
Ls2_Ind    (23  34) inductor l=Ls2*(1+dls_3Tdiff_1talpa)
Rs2_Ind    (34 MINUS) resistor r=Rs2*(1+drs_3Tdiff_1talpa) tc1=0.003
Lp1_Ind    (56 12) inductor l=Lp1
Rp1_Ind    (PLUS 56) resistor r=Rp1 tc1=0.003
Lp2_Ind    (78 MINUS) inductor l=Lp2
Rp2_Ind    (34 78) resistor r=Rp2 tc1=0.003
Cox1_Ind   (PLUS  11) capacitor c=Cox1
Rsub1_Ind  (11  0) resistor r=Rsub1
Csub1_Ind  (11  0) capacitor c=Csub1
Cox2_Ind   (MINUS  22) capacitor c=Cox2
Rsub2_Ind  (22  0) resistor r=Rsub2
Csub2_Ind  (22  0) capacitor c=Csub2
Lshort_Ind   (23  31) inductor l=Lshort
Rshort_Ind  (31  CT) resistor r=Rshort*(1+drs_3Tdiff_1talpa) tc1=0.003
Rssk_Ind  (31  32) resistor r=Rssk tc1=0.003  
Lssk_Ind  (32  CT) inductor l=Lssk  
Klm1      mutual_inductor coupling=mm ind1=Ls1_Ind ind2=Ls2_Ind

ends rf_3Tdiff_1talpa_t2
 
subckt rf_3Tdiff_1talpa_t3 (PLUS MINUS CT)
// ***********************************************************************************
//***PLUS=port1, MINUS=port2**//
//***0.11um 3 turns 3-T differential inductor scalable model**//
//***R=inner radius; N=turns; W=width; S=spacing**//
//***In this model, R is scalalbe, N=3, S=2.0um, W=15um**//
// ***********************************************************************************
parameters R=50.0e-6 N=3 
+Ldc1=6.6156e-5*pwr(R,1.1142)
+Rdc1=5758.6*R+0.30052 
+Ldc2=Ldc1
+Rdc2=Rdc1 
+Cox1=6e-14
+Csub1=5e-10*R+4.5e-14
+Rsub1=-5000000*R+1200
+Cox2=Cox1
+Csub2=Csub1
+Rsub2=Rsub1 
+Cf=7.3103e-10*R+1.7362e-14
+mm=0.55
+Lsshort=1.8813e-10*exp(-18594*R)
+Rsshort=0.37
+Krssk=5 
+Klssk=1 
+Krp=0.32307*log(R)+3.5207 
+Klp=0.23 
+Ls1=1/(1+Klp/pwr(1+Krp,2))*Ldc1/2
+Ls2=1/(1+Klp/pwr(1+Krp,2))*Ldc2/2
+Rs1=(1+1/Krp)*Rdc1/2
+Rs2=(1+1/Krp)*Rdc2/2
+Rp1=Krp*Rs1
+Rp2=Krp*Rs2
+Lp1=Klp*Ls1
+Lp2=Klp*Ls2
+Lshort=Lsshort
+Lssk=Lsshort*Klssk
+Rshort=Rsshort
+Rssk=Rsshort*Krssk
//***equivalent circuit
Cf_Ind     (PLUS  MINUS) capacitor c=Cf
Ls1_Ind    (12  23) inductor l=Ls1*(1+dls_3Tdiff_1talpa)
Rs1_Ind    (PLUS 12) resistor r=Rs1*(1+drs_3Tdiff_1talpa) tc1=0.003
Ls2_Ind    (23  34) inductor l=Ls2*(1+dls_3Tdiff_1talpa)
Rs2_Ind    (34 MINUS) resistor r=Rs2*(1+drs_3Tdiff_1talpa) tc1=0.003
Lp1_Ind    (56 12) inductor l=Lp1
Rp1_Ind    (PLUS 56) resistor r=Rp1 tc1=0.003
Lp2_Ind    (78 MINUS) inductor l=Lp2
Rp2_Ind    (34 78) resistor r=Rp2 tc1=0.003
Cox1_Ind   (PLUS  11) capacitor c=Cox1
Rsub1_Ind  (11  0) resistor r=Rsub1
Csub1_Ind  (11  0) capacitor c=Csub1
Cox2_Ind   (MINUS  22) capacitor c=Cox2
Rsub2_Ind  (22  0) resistor r=Rsub2
Csub2_Ind  (22  0) capacitor c=Csub2
Lshort_Ind   (23  31) inductor l=Lshort
Rshort_Ind  (31  CT) resistor r=Rshort*(1+drs_3Tdiff_1talpa) tc1=0.003
Rssk_Ind  (31  32) resistor r=Rssk tc1=0.003  
Lssk_Ind  (32  CT) inductor l=Lssk  
Klm1      mutual_inductor coupling=mm ind1=Ls1_Ind ind2=Ls2_Ind

ends rf_3Tdiff_1talpa_t3

subckt rf_3Tdiff_1talpa_t4 (PLUS MINUS CT)
// ***********************************************************************************
//***PLUS=port1, MINUS=port2**//
//***0.11um 4 turns 3-T differential inductor scalable model**//
//***R=inner radius; N=turns; W=width; S=spacing**//
//***In this model, R is scalalbe, N=4, S=2.0um, W=15um**//
// ***********************************************************************************
parameters R=50.0e-6 N=4 
+Ldc1=4.2336e-5*R-1.2983e-10
+Rdc1=7551.7*R+0.5131 
+Ldc2=Ldc1
+Rdc2=7172.4*R+0.43534 
+Cox1=7.5e-14
+Csub1=5e-10*R+3e-14
+Rsub1=900
+Cox2=Cox1
+Csub2=Csub1
+Rsub2=Rsub1 
+Cf=1.1259e-9*R+3.8052e-14
+mm=0.55
+Lsshort=-6.7241e-7*R+1.1966e-10
+Rsshort=0.65047*exp(6275.5*R)
+Krssk=5 
+Klssk=1 
+Krp=0.39777*log(R)+4.3174 
+Klp=0.32 
+Ls1=1/(1+Klp/pwr(1+Krp,2))*Ldc1/2
+Ls2=1/(1+Klp/pwr(1+Krp,2))*Ldc2/2
+Rs1=(1+1/Krp)*Rdc1/2
+Rs2=(1+1/Krp)*Rdc2/2
+Rp1=Krp*Rs1
+Rp2=Krp*Rs2
+Lp1=Klp*Ls1
+Lp2=Klp*Ls2
+Lshort=Lsshort
+Lssk=Lsshort*Klssk
+Rshort=Rsshort
+Rssk=Rsshort*Krssk

//***equivalent circuit
Cf_Ind     (PLUS  MINUS) capacitor c=Cf
Ls1_Ind    (12  23) inductor l=Ls1*(1+dls_3Tdiff_1talpa)
Rs1_Ind    (PLUS 12) resistor r=Rs1*(1+drs_3Tdiff_1talpa) tc1=0.003
Ls2_Ind    (23  34) inductor l=Ls2*(1+dls_3Tdiff_1talpa)
Rs2_Ind    (34 MINUS) resistor r=Rs2*(1+drs_3Tdiff_1talpa) tc1=0.003
Lp1_Ind    (56 12) inductor l=Lp1
Rp1_Ind    (PLUS 56) resistor r=Rp1 tc1=0.003
Lp2_Ind    (78 MINUS) inductor l=Lp2
Rp2_Ind    (34 78) resistor r=Rp2 tc1=0.003
Cox1_Ind   (PLUS  11) capacitor c=Cox1
Rsub1_Ind  (11  0) resistor r=Rsub1
Csub1_Ind  (11  0) capacitor c=Csub1
Cox2_Ind   (MINUS  22) capacitor c=Cox2
Rsub2_Ind  (22  0) resistor r=Rsub2
Csub2_Ind  (22  0) capacitor c=Csub2
Lshort_Ind   (23  31) inductor l=Lshort
Rshort_Ind  (31  CT) resistor r=Rshort*(1+drs_3Tdiff_1talpa) tc1=0.003
Rssk_Ind  (31  32) resistor r=Rssk tc1=0.003  
Lssk_Ind  (32  CT) inductor l=Lssk  
Klm1      mutual_inductor coupling=mm ind1=Ls1_Ind ind2=Ls2_Ind

ends rf_3Tdiff_1talpa_t4

subckt rf_3Tdiff_1talpa_t5 (PLUS MINUS CT)
// ***********************************************************************************
//***PLUS=port1, MINUS=port2**//
//***0.11um 5 turns 3-T differential inductor scalable model**//
//***R=inner radius; N=turns; W=width; S=spacing**//
//***In this model, R is scalalbe, N=5, S=2.0um, W=15um**//
// ***********************************************************************************
parameters R=50.0e-6 N=5 
+Ldc1=5.5638e-5*R+1.9328e-10
+Rdc1=8793.1*R+0.70259 
+Ldc2=Ldc1
+Rdc2=Rdc1 
+Cox1=9.5e-14
+Csub1=5e-10*R+5e-14
+Rsub1=900
+Cox2=Cox1
+Csub2=Csub1
+Rsub2=Rsub1 
+Cf=1.5017e-9*R+6.2603e-14
+mm=0.75
+Lsshort=8.5e-11
+Rsshort=0.5
+Krssk=5 
+Klssk=1 
+Krp=627.38*pwr(R,0.7376) 
+Klp=0.39 
+Ls1=1/(1+Klp/pwr(1+Krp,2))*Ldc1/2
+Ls2=1/(1+Klp/pwr(1+Krp,2))*Ldc2/2
+Rs1=(1+1/Krp)*Rdc1/2
+Rs2=(1+1/Krp)*Rdc2/2
+Rp1=Krp*Rs1
+Rp2=Krp*Rs2
+Lp1=Klp*Ls1
+Lp2=Klp*Ls2
+Lshort=Lsshort
+Lssk=Lsshort*Klssk
+Rshort=Rsshort
+Rssk=Rsshort*Krssk

//***equivalent circuit

Cf_Ind     (PLUS  MINUS) capacitor c=Cf
Ls1_Ind    (12  23) inductor l=Ls1*(1+dls_3Tdiff_1talpa)
Rs1_Ind    (PLUS 12) resistor r=Rs1*(1+drs_3Tdiff_1talpa) tc1=0.003
Ls2_Ind    (23  34) inductor l=Ls2*(1+dls_3Tdiff_1talpa)
Rs2_Ind    (34 MINUS) resistor r=Rs2*(1+drs_3Tdiff_1talpa) tc1=0.003
Lp1_Ind    (56 12) inductor l=Lp1
Rp1_Ind    (PLUS 56) resistor r=Rp1 tc1=0.003
Lp2_Ind    (78 MINUS) inductor l=Lp2
Rp2_Ind    (34 78) resistor r=Rp2 tc1=0.003
Cox1_Ind   (PLUS  11) capacitor c=Cox1
Rsub1_Ind  (11  0) resistor r=Rsub1
Csub1_Ind  (11  0) capacitor c=Csub1
Cox2_Ind   (MINUS  22) capacitor c=Cox2
Rsub2_Ind  (22  0) resistor r=Rsub2
Csub2_Ind  (22  0) capacitor c=Csub2
Lshort_Ind   (23  31) inductor l=Lshort
Rshort_Ind  (31  CT) resistor r=Rshort*(1+drs_3Tdiff_1talpa) tc1=0.003
Rssk_Ind  (31  32) resistor r=Rssk tc1=0.003  
Lssk_Ind  (32  CT) inductor l=Lssk  
Klm1      mutual_inductor coupling=mm ind1=Ls1_Ind ind2=Ls2_Ind

ends rf_3Tdiff_1talpa_t5


subckt rf_3Tdiff_1talpa_t6 (PLUS MINUS CT)
// ***********************************************************************************
//***PLUS=port1, MINUS=port2**//
//***0.11um 6 turns 3-T differential inductor scalable model**//
//***R=inner radius; N=turns; W=width; S=spacing**//
//***In this model, R is scalalbe, N=6, S=2.0um, W=15um**//
// ***********************************************************************************
parameters R=50.0e-6 N=6 
+Ldc1=7.5897e-5*R+5.8879e-10
+Rdc1=11052*R+0.9831 
+Ldc2=Ldc1
+Rdc2=11224*R+0.85845 
+Cox1=1.05e-13
+Csub1=5e-10*R+5.5e-14
+Rsub1=1200
+Cox2=Cox1
+Csub2=Csub1
+Rsub2=Rsub1 
+Cf=2.0362e-9*R+8.9172e-14
+mm=0.75
+Lsshort=1.2e-10
+Rsshort=7327.6*R+0.61466
+Krssk=5 
+Klssk=1 
+Krp=2055.5*pwr(R,0.86997) 
+Klp=-413.79*R+0.36017 
+Ls1=1/(1+Klp/pwr(1+Krp,2))*Ldc1/2
+Ls2=1/(1+Klp/pwr(1+Krp,2))*Ldc2/2
+Rs1=(1+1/Krp)*Rdc1/2
+Rs2=(1+1/Krp)*Rdc2/2
+Rp1=Krp*Rs1
+Rp2=Krp*Rs2
+Lp1=Klp*Ls1
+Lp2=Klp*Ls2
+Lshort=Lsshort
+Lssk=Lsshort*Klssk
+Rshort=Rsshort
+Rssk=Rsshort*Krssk

//***equivalent circuit

Cf_Ind     (PLUS  MINUS) capacitor c=Cf
Ls1_Ind    (12  23) inductor l=Ls1*(1+dls_3Tdiff_1talpa)
Rs1_Ind    (PLUS 12) resistor r=Rs1*(1+drs_3Tdiff_1talpa) tc1=0.003
Ls2_Ind    (23  34) inductor l=Ls2*(1+dls_3Tdiff_1talpa)
Rs2_Ind    (34 MINUS) resistor r=Rs2*(1+drs_3Tdiff_1talpa) tc1=0.003
Lp1_Ind    (56 12) inductor l=Lp1
Rp1_Ind    (PLUS 56) resistor r=Rp1 tc1=0.003
Lp2_Ind    (78 MINUS) inductor l=Lp2
Rp2_Ind    (34 78) resistor r=Rp2 tc1=0.003
Cox1_Ind   (PLUS  11) capacitor c=Cox1
Rsub1_Ind  (11  0) resistor r=Rsub1
Csub1_Ind  (11  0) capacitor c=Csub1
Cox2_Ind   (MINUS  22) capacitor c=Cox2
Rsub2_Ind  (22  0) resistor r=Rsub2
Csub2_Ind  (22  0) capacitor c=Csub2
Lshort_Ind   (23  31) inductor l=Lshort
Rshort_Ind  (31  CT) resistor r=Rshort*(1+drs_3Tdiff_1talpa) tc1=0.003
Rssk_Ind  (31  32) resistor r=Rssk tc1=0.003  
Lssk_Ind  (32  CT) inductor l=Lssk  
Klm1      mutual_inductor coupling=mm ind1=Ls1_Ind ind2=Ls2_Ind

ends rf_3Tdiff_1talpa_t6

subckt rf_3Tdiff_1talpa_t7 (PLUS MINUS CT)
// ***********************************************************************************
//***PLUS=port1, MINUS=port2**//
//***0.11um 7 turns 3-T differential inductor scalable model**//
//***R=inner radius; N=turns; W=width; S=spacing**//
//***In this model, R is scalalbe, N=7, S=2.0um, W=15um**//
// ***********************************************************************************
parameters R=50.0e-6 N=7 
+Ldc1=8.6469e-5*R+1.3984e-9
+Rdc1=1.3449*exp(6031.1*R) 
+Ldc2=Ldc1
+Rdc2=Rdc1 
+Cox1=7.5e-14
+Csub1=7.5e-14
+Rsub1=800
+Cox2=Cox1
+Csub2=Csub1
+Rsub2=Rsub1 
+Cf=5.6495e-11*pwr(R,0.54411)
+mm=0.98
+Lsshort=1.4916e-10*exp(6337.4*R)
+Rsshort=0.6
+Krssk=5 
+Klssk=1 
+Krp=3423.1*R+0.20859 
+Klp=-1153.8*R+0.41718 
+Ls1=1/(1+Klp/pwr(1+Krp,2))*Ldc1/2
+Ls2=1/(1+Klp/pwr(1+Krp,2))*Ldc2/2
+Rs1=(1+1/Krp)*Rdc1/2
+Rs2=(1+1/Krp)*Rdc2/2
+Rp1=Krp*Rs1
+Rp2=Krp*Rs2
+Lp1=Klp*Ls1
+Lp2=Klp*Ls2
+Lshort=Lsshort
+Lssk=Lsshort*Klssk
+Rshort=Rsshort
+Rssk=Rsshort*Krssk

//***equivalent circuit

Cf_Ind     (PLUS  MINUS) capacitor c=Cf
Ls1_Ind    (12  23) inductor l=Ls1*(1+dls_3Tdiff_1talpa)
Rs1_Ind    (PLUS 12) resistor r=Rs1*(1+drs_3Tdiff_1talpa) tc1=0.003
Ls2_Ind    (23  34) inductor l=Ls2*(1+dls_3Tdiff_1talpa)
Rs2_Ind    (34 MINUS) resistor r=Rs2*(1+drs_3Tdiff_1talpa) tc1=0.003
Lp1_Ind    (56 12) inductor l=Lp1
Rp1_Ind    (PLUS 56) resistor r=Rp1 tc1=0.003
Lp2_Ind    (78 MINUS) inductor l=Lp2
Rp2_Ind    (34 78) resistor r=Rp2 tc1=0.003
Cox1_Ind   (PLUS  11) capacitor c=Cox1
Rsub1_Ind  (11  0) resistor r=Rsub1
Csub1_Ind  (11  0) capacitor c=Csub1
Cox2_Ind   (MINUS  22) capacitor c=Cox2
Rsub2_Ind  (22  0) resistor r=Rsub2
Csub2_Ind  (22  0) capacitor c=Csub2
Lshort_Ind   (23  31) inductor l=Lshort
Rshort_Ind  (31  CT) resistor r=Rshort*(1+drs_3Tdiff_1talpa) tc1=0.003
Rssk_Ind  (31  32) resistor r=Rssk tc1=0.003  
Lssk_Ind  (32  CT) inductor l=Lssk  
Klm1      mutual_inductor coupling=mm ind1=Ls1_Ind ind2=Ls2_Ind

ends rf_3Tdiff_1talpa_t7