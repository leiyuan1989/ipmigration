****Sub-Circuit for AC1CINHSV1, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC1CINHSV1 A B CIN CO VDD VSS
MM41 net0196 CIN net78 VPW N12LL W=180.00n L=60.00n
MM42 net0144 cinn net78 VPW N12LL W=180.00n L=60.00n
MM3 net0144 A VSS VPW N12LL W=180.00n L=60.00n
MM2 net0144 B VSS VPW N12LL W=180.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=220.00n L=60.00n
MM11 net0196 A net0124 VPW N12LL W=220.00n L=60.00n
MM27 cinn CIN VSS VPW N12LL W=180.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=350.00n L=60.00n
MM43 net0196 cinn net78 VNW P12LL W=220.00n L=60.00n
MM44 net0144 CIN net78 VNW P12LL W=220.00n L=60.00n
MM12 net0196 A VDD VNW P12LL W=180.00n L=60.00n
MM13 net0196 B VDD VNW P12LL W=180.00n L=60.00n
MM28 cinn CIN VDD VNW P12LL W=220.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=440.00n L=60.00n
MM4 net0144 A net0215 VNW P12LL W=250.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=250.00n L=60.00n
.ENDS AC1CINHSV1
****Sub-Circuit for AC1CINHSV2, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC1CINHSV2 A B CIN CO VDD VSS
MM41 net0196 CIN net78 VPW N12LL W=220.00n L=60.00n
MM42 net0144 cinn net78 VPW N12LL W=220.00n L=60.00n
MM3 net0144 A VSS VPW N12LL W=180.00n L=60.00n
MM2 net0144 B VSS VPW N12LL W=180.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=260.00n L=60.00n
MM11 net0196 A net0124 VPW N12LL W=260.00n L=60.00n
MM27 cinn CIN VSS VPW N12LL W=220.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=430.00n L=60.00n
MM43 net0196 cinn net78 VNW P12LL W=270.00n L=60.00n
MM44 net0144 CIN net78 VNW P12LL W=270.00n L=60.00n
MM12 net0196 A VDD VNW P12LL W=220.00n L=60.00n
MM13 net0196 B VDD VNW P12LL W=220.00n L=60.00n
MM28 cinn CIN VDD VNW P12LL W=270.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=540.00n L=60.00n
MM4 net0144 A net0215 VNW P12LL W=280.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=280.00n L=60.00n
.ENDS AC1CINHSV2
****Sub-Circuit for AC1CINHSV4, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC1CINHSV4 A B CIN CO VDD VSS
MM41 net0196 CIN net78 VPW N12LL W=430.00n L=60.00n
MM42 net0144 cinn net78 VPW N12LL W=430.00n L=60.00n
MM3 net0144 A VSS VPW N12LL W=240.00n L=60.00n
MM2 net0144 B VSS VPW N12LL W=240.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=430.00n L=60.00n
MM11 net0196 A net0124 VPW N12LL W=430.00n L=60.00n
MM27 cinn CIN VSS VPW N12LL W=220.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=860.00n L=60.00n
MM43 net0196 cinn net78 VNW P12LL W=540.00n L=60.00n
MM44 net0144 CIN net78 VNW P12LL W=540.00n L=60.00n
MM12 net0196 A VDD VNW P12LL W=420.00n L=60.00n
MM13 net0196 B VDD VNW P12LL W=420.00n L=60.00n
MM28 cinn CIN VDD VNW P12LL W=270.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=1.08u L=60.00n
MM4 net0144 A net0215 VNW P12LL W=440.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=440.00n L=60.00n
.ENDS AC1CINHSV4
****Sub-Circuit for AC1CONHSV1, Thu May 19 13:57:40 CST 2011****
.SUBCKT AC1CONHSV1 A B CI CON VDD VSS
MM16 net0133 net0286 VSS VPW N12LL W=180.00n L=60.00n
MM41 net0196 cin net78 VPW N12LL W=180.00n L=60.00n
MM42 net0133 CI net78 VPW N12LL W=180.00n L=60.00n
MM3 net0286 A VSS VPW N12LL W=180.00n L=60.00n
MM2 net0286 B VSS VPW N12LL W=180.00n L=60.00n
MM14 net0196 net0193 VSS VPW N12LL W=180.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=220.00n L=60.00n
MM11 net0193 A net0124 VPW N12LL W=220.00n L=60.00n
MM27 cin CI VSS VPW N12LL W=180.00n L=60.00n
MM22 CON net78 VSS VPW N12LL W=350.00n L=60.00n
MM17 net0133 net0286 VDD VNW P12LL W=220.00n L=60.00n
MM43 net0196 CI net78 VNW P12LL W=220.00n L=60.00n
MM44 net0133 cin net78 VNW P12LL W=220.00n L=60.00n
MM15 net0196 net0193 VDD VNW P12LL W=220.00n L=60.00n
MM12 net0193 A VDD VNW P12LL W=180.00n L=60.00n
MM13 net0193 B VDD VNW P12LL W=180.00n L=60.00n
MM28 cin CI VDD VNW P12LL W=220.00n L=60.00n
MM21 CON net78 VDD VNW P12LL W=440.00n L=60.00n
MM4 net0286 A net0215 VNW P12LL W=250.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=250.00n L=60.00n
.ENDS AC1CONHSV1
****Sub-Circuit for AC1CONHSV2, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC1CONHSV2 A B CI CON VDD VSS
MM16 net0133 net0286 VSS VPW N12LL W=220.00n L=60.00n
MM41 net0196 cin net78 VPW N12LL W=220.00n L=60.00n
MM42 net0133 CI net78 VPW N12LL W=220.00n L=60.00n
MM3 net0286 A VSS VPW N12LL W=180.00n L=60.00n
MM2 net0286 B VSS VPW N12LL W=180.00n L=60.00n
MM14 net0196 net0193 VSS VPW N12LL W=220.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=260.00n L=60.00n
MM11 net0193 A net0124 VPW N12LL W=260.00n L=60.00n
MM27 cin CI VSS VPW N12LL W=220.00n L=60.00n
MM22 CON net78 VSS VPW N12LL W=430.00n L=60.00n
MM17 net0133 net0286 VDD VNW P12LL W=270.00n L=60.00n
MM43 net0196 CI net78 VNW P12LL W=270.00n L=60.00n
MM44 net0133 cin net78 VNW P12LL W=270.00n L=60.00n
MM15 net0196 net0193 VDD VNW P12LL W=270.00n L=60.00n
MM12 net0193 A VDD VNW P12LL W=220.00n L=60.00n
MM13 net0193 B VDD VNW P12LL W=220.00n L=60.00n
MM28 cin CI VDD VNW P12LL W=270.00n L=60.00n
MM21 CON net78 VDD VNW P12LL W=540.00n L=60.00n
MM4 net0286 A net0215 VNW P12LL W=280.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=280.00n L=60.00n
.ENDS AC1CONHSV2
****Sub-Circuit for AC1CONHSV4, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC1CONHSV4 A B CI CON VDD VSS
MM16 net0133 net0286 VSS VPW N12LL W=430.00n L=60.00n
MM41 net0196 cin net78 VPW N12LL W=430.00n L=60.00n
MM42 net0133 CI net78 VPW N12LL W=430.00n L=60.00n
MM3 net0286 A VSS VPW N12LL W=240.00n L=60.00n
MM2 net0286 B VSS VPW N12LL W=240.00n L=60.00n
MM14 net0196 net0193 VSS VPW N12LL W=430.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=430.00n L=60.00n
MM11 net0193 A net0124 VPW N12LL W=430.00n L=60.00n
MM27 cin CI VSS VPW N12LL W=220.00n L=60.00n
MM22 CON net78 VSS VPW N12LL W=860.00n L=60.00n
MM17 net0133 net0286 VDD VNW P12LL W=540.00n L=60.00n
MM43 net0196 CI net78 VNW P12LL W=540.00n L=60.00n
MM44 net0133 cin net78 VNW P12LL W=540.00n L=60.00n
MM15 net0196 net0193 VDD VNW P12LL W=540.00n L=60.00n
MM12 net0193 A VDD VNW P12LL W=440.00n L=60.00n
MM13 net0193 B VDD VNW P12LL W=440.00n L=60.00n
MM28 cin CI VDD VNW P12LL W=270.00n L=60.00n
MM21 CON net78 VDD VNW P12LL W=1.08u L=60.00n
MM4 net0286 A net0215 VNW P12LL W=440.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=440.00n L=60.00n
.ENDS AC1CONHSV4
****Sub-Circuit for AC2CINHSV1, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC2CINHSV1 A B CI0N CI1N CO0 CO1 VDD VSS
MM51 ci1nn CI1N VSS VPW N12LL W=180.00n L=60.00n
MM48 ci0nn CI0N VSS VPW N12LL W=180.00n L=60.00n
MM3 norab A VSS VPW N12LL W=180.00n L=60.00n
MM18 net0132 B VSS VPW N12LL W=260.00n L=60.00n
MM23 nandab A net0132 VPW N12LL W=260.00n L=60.00n
MM2 norab B VSS VPW N12LL W=180.00n L=60.00n
MM26 nandab CI0N net0143 VPW N12LL W=180.00n L=60.00n
MM29 norab ci0nn net0143 VPW N12LL W=180.00n L=60.00n
MM30 CO0 net0143 VSS VPW N12LL W=350.00n L=60.00n
MM34 nandab CI1N net0155 VPW N12LL W=180.00n L=60.00n
MM35 norab ci1nn net0155 VPW N12LL W=180.00n L=60.00n
MM37 CO1 net0155 VSS VPW N12LL W=350.00n L=60.00n
MM50 ci1nn CI1N VDD VNW P12LL W=220.00n L=60.00n
MM49 ci0nn CI0N VDD VNW P12LL W=220.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=220.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=220.00n L=60.00n
MM31 nandab ci0nn net0143 VNW P12LL W=220.00n L=60.00n
MM32 norab CI0N net0143 VNW P12LL W=220.00n L=60.00n
MM33 CO0 net0143 VDD VNW P12LL W=440.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=280.00n L=60.00n
MM45 nandab ci1nn net0155 VNW P12LL W=220.00n L=60.00n
MM46 norab CI1N net0155 VNW P12LL W=220.00n L=60.00n
MM47 CO1 net0155 VDD VNW P12LL W=440.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=280.00n L=60.00n
.ENDS AC2CINHSV1
****Sub-Circuit for AC2CINHSV2, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC2CINHSV2 A B CI0N CI1N CO0 CO1 VDD VSS
MM51 ci1nn CI1N VSS VPW N12LL W=220.00n L=60.00n
MM48 ci0nn CI0N VSS VPW N12LL W=220.00n L=60.00n
MM3 norab A VSS VPW N12LL W=240.00n L=60.00n
MM18 net0132 B VSS VPW N12LL W=430.00n L=60.00n
MM23 nandab A net0132 VPW N12LL W=430.00n L=60.00n
MM2 norab B VSS VPW N12LL W=240.00n L=60.00n
MM26 nandab CI0N net0143 VPW N12LL W=220.00n L=60.00n
MM29 norab ci0nn net0143 VPW N12LL W=220.00n L=60.00n
MM30 CO0 net0143 VSS VPW N12LL W=430.00n L=60.00n
MM34 nandab CI1N net0155 VPW N12LL W=220.00n L=60.00n
MM35 norab ci1nn net0155 VPW N12LL W=220.00n L=60.00n
MM37 CO1 net0155 VSS VPW N12LL W=430.00n L=60.00n
MM50 ci1nn CI1N VDD VNW P12LL W=270.00n L=60.00n
MM49 ci0nn CI0N VDD VNW P12LL W=270.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=440.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=440.00n L=60.00n
MM31 nandab ci0nn net0143 VNW P12LL W=270.00n L=60.00n
MM32 norab CI0N net0143 VNW P12LL W=270.00n L=60.00n
MM33 CO0 net0143 VDD VNW P12LL W=540.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=440.00n L=60.00n
MM45 nandab ci1nn net0155 VNW P12LL W=270.00n L=60.00n
MM46 norab CI1N net0155 VNW P12LL W=270.00n L=60.00n
MM47 CO1 net0155 VDD VNW P12LL W=540.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=440.00n L=60.00n
.ENDS AC2CINHSV2
****Sub-Circuit for AC2CINHSV4, Mon Jan 24 17:06:27 CST 2011****
.SUBCKT AC2CINHSV4 A B CI0N CI1N CO0 CO1 VDD VSS
MM51 ci1nn CI1N VSS VPW N12LL W=220.00n L=60.00n
MM48 ci0nn CI0N VSS VPW N12LL W=220.00n L=60.00n
MM3 norab A VSS VPW N12LL W=480.00n L=60.00n
MM18 net0132 B VSS VPW N12LL W=860.00n L=60.00n
MM23 nandab A net0132 VPW N12LL W=860.00n L=60.00n
MM2 norab B VSS VPW N12LL W=480.00n L=60.00n
MM26 nandab CI0N net0143 VPW N12LL W=430.00n L=60.00n
MM29 norab ci0nn net0143 VPW N12LL W=430.00n L=60.00n
MM30 CO0 net0143 VSS VPW N12LL W=860.00n L=60.00n
MM34 nandab CI1N net0155 VPW N12LL W=430.00n L=60.00n
MM35 norab ci1nn net0155 VPW N12LL W=430.00n L=60.00n
MM37 CO1 net0155 VSS VPW N12LL W=860.00n L=60.00n
MM50 ci1nn CI1N VDD VNW P12LL W=270.00n L=60.00n
MM49 ci0nn CI0N VDD VNW P12LL W=270.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=880.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=880.00n L=60.00n
MM31 nandab ci0nn net0143 VNW P12LL W=540.00n L=60.00n
MM32 norab CI0N net0143 VNW P12LL W=540.00n L=60.00n
MM33 CO0 net0143 VDD VNW P12LL W=1.08u L=60.00n
MM4 norab A net0215 VNW P12LL W=880.00n L=60.00n
MM45 nandab ci1nn net0155 VNW P12LL W=540.00n L=60.00n
MM46 norab CI1N net0155 VNW P12LL W=540.00n L=60.00n
MM47 CO1 net0155 VDD VNW P12LL W=1.08u L=60.00n
MM5 net0215 B VDD VNW P12LL W=880.00n L=60.00n
.ENDS AC2CINHSV4
****Sub-Circuit for AC2CONHSV1, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC2CONHSV1 A B CI0 CI1 CO0N CO1N VDD VSS
MM50 ci1n CI1 VDD VNW P12LL W=220.00n L=60.00n
MM49 ci0n CI0 VDD VNW P12LL W=220.00n L=60.00n
MM77 andab nandab VDD VNW P12LL W=220.00n L=60.00n
MM76 orab norab VDD VNW P12LL W=220.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=220.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=220.00n L=60.00n
MM45 andab CI1 net176 VNW P12LL W=220.00n L=60.00n
MM46 orab ci1n net176 VNW P12LL W=220.00n L=60.00n
MM47 CO1N net176 VDD VNW P12LL W=440.00n L=60.00n
MM31 andab CI0 net188 VNW P12LL W=220.00n L=60.00n
MM32 orab ci0n net188 VNW P12LL W=220.00n L=60.00n
MM33 CO0N net188 VDD VNW P12LL W=440.00n L=60.00n
MM4 norab A net144 VNW P12LL W=280.00n L=60.00n
MM5 net144 B VDD VNW P12LL W=280.00n L=60.00n
MM51 ci1n CI1 VSS VPW N12LL W=180.00n L=60.00n
MM48 ci0n CI0 VSS VPW N12LL W=180.00n L=60.00n
MM26 andab ci0n net188 VPW N12LL W=180.00n L=60.00n
MM29 orab CI0 net188 VPW N12LL W=180.00n L=60.00n
MM30 CO0N net188 VSS VPW N12LL W=350.00n L=60.00n
MM34 andab ci1n net176 VPW N12LL W=180.00n L=60.00n
MM35 orab CI1 net176 VPW N12LL W=180.00n L=60.00n
MM37 CO1N net176 VSS VPW N12LL W=350.00n L=60.00n
MM75 andab nandab VSS VPW N12LL W=180.00n L=60.00n
MM74 orab norab VSS VPW N12LL W=180.00n L=60.00n
MM3 norab A VSS VPW N12LL W=180.00n L=60.00n
MM2 norab B VSS VPW N12LL W=180.00n L=60.00n
MM18 net209 B VSS VPW N12LL W=260.00n L=60.00n
MM23 nandab A net209 VPW N12LL W=260.00n L=60.00n
.ENDS AC2CONHSV1
****Sub-Circuit for AC2CONHSV2, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC2CONHSV2 A B CI0 CI1 CO0N CO1N VDD VSS
MM50 ci1n CI1 VDD VNW P12LL W=270.00n L=60.00n
MM49 ci0n CI0 VDD VNW P12LL W=270.00n L=60.00n
MM77 andab nandab VDD VNW P12LL W=270.00n L=60.00n
MM76 orab norab VDD VNW P12LL W=270.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=440.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=440.00n L=60.00n
MM45 andab CI1 net176 VNW P12LL W=270.00n L=60.00n
MM46 orab ci1n net176 VNW P12LL W=270.00n L=60.00n
MM47 CO1N net176 VDD VNW P12LL W=540.00n L=60.00n
MM31 andab CI0 net188 VNW P12LL W=270.00n L=60.00n
MM32 orab ci0n net188 VNW P12LL W=270.00n L=60.00n
MM33 CO0N net188 VDD VNW P12LL W=540.00n L=60.00n
MM4 norab A net144 VNW P12LL W=440.00n L=60.00n
MM5 net144 B VDD VNW P12LL W=440.00n L=60.00n
MM51 ci1n CI1 VSS VPW N12LL W=220.00n L=60.00n
MM48 ci0n CI0 VSS VPW N12LL W=220.00n L=60.00n
MM26 andab ci0n net188 VPW N12LL W=220.00n L=60.00n
MM29 orab CI0 net188 VPW N12LL W=220.00n L=60.00n
MM30 CO0N net188 VSS VPW N12LL W=430.00n L=60.00n
MM34 andab ci1n net176 VPW N12LL W=220.00n L=60.00n
MM35 orab CI1 net176 VPW N12LL W=220.00n L=60.00n
MM37 CO1N net176 VSS VPW N12LL W=430.00n L=60.00n
MM75 andab nandab VSS VPW N12LL W=220.00n L=60.00n
MM74 orab norab VSS VPW N12LL W=220.00n L=60.00n
MM3 norab A VSS VPW N12LL W=240.00n L=60.00n
MM2 norab B VSS VPW N12LL W=240.00n L=60.00n
MM18 net209 B VSS VPW N12LL W=430.00n L=60.00n
MM23 nandab A net209 VPW N12LL W=430.00n L=60.00n
.ENDS AC2CONHSV2
****Sub-Circuit for AC2CONHSV4, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AC2CONHSV4 A B CI0 CI1 CO0N CO1N VDD VSS
MM50 ci1n CI1 VDD VNW P12LL W=270.00n L=60.00n
MM49 ci0n CI0 VDD VNW P12LL W=270.00n L=60.00n
MM77 andab nandab VDD VNW P12LL W=540.00n L=60.00n
MM76 orab norab VDD VNW P12LL W=540.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=880.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=880.00n L=60.00n
MM45 andab CI1 net176 VNW P12LL W=540.00n L=60.00n
MM46 orab ci1n net176 VNW P12LL W=540.00n L=60.00n
MM47 CO1N net176 VDD VNW P12LL W=1.08u L=60.00n
MM31 andab CI0 net188 VNW P12LL W=540.00n L=60.00n
MM32 orab ci0n net188 VNW P12LL W=540.00n L=60.00n
MM33 CO0N net188 VDD VNW P12LL W=1.08u L=60.00n
MM4 norab A net144 VNW P12LL W=880.00n L=60.00n
MM5 net144 B VDD VNW P12LL W=880.00n L=60.00n
MM51 ci1n CI1 VSS VPW N12LL W=220.00n L=60.00n
MM48 ci0n CI0 VSS VPW N12LL W=220.00n L=60.00n
MM26 andab ci0n net188 VPW N12LL W=430.00n L=60.00n
MM29 orab CI0 net188 VPW N12LL W=430.00n L=60.00n
MM30 CO0N net188 VSS VPW N12LL W=860.00n L=60.00n
MM34 andab ci1n net176 VPW N12LL W=430.00n L=60.00n
MM35 orab CI1 net176 VPW N12LL W=430.00n L=60.00n
MM37 CO1N net176 VSS VPW N12LL W=860.00n L=60.00n
MM75 andab nandab VSS VPW N12LL W=430.00n L=60.00n
MM74 orab norab VSS VPW N12LL W=430.00n L=60.00n
MM3 norab A VSS VPW N12LL W=480.00n L=60.00n
MM2 norab B VSS VPW N12LL W=480.00n L=60.00n
MM18 net209 B VSS VPW N12LL W=860.00n L=60.00n
MM23 nandab A net209 VPW N12LL W=860.00n L=60.00n
.ENDS AC2CONHSV4
****Sub-Circuit for ACH2CONHSV1, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT ACH2CONHSV1 A B CO0N CO1N VDD VSS
MM5 net50 B VDD VNW P12LL W=520.00n L=60.00n
MM4 CO1N A net50 VNW P12LL W=520.00n L=60.00n
MM13 CO0N B VDD VNW P12LL W=390.00n L=60.00n
MM12 CO0N A VDD VNW P12LL W=390.00n L=60.00n
MM11 CO0N A net83 VPW N12LL W=430.00n L=60.00n
MM10 net83 B VSS VPW N12LL W=430.00n L=60.00n
MM2 CO1N B VSS VPW N12LL W=280.00n L=60.00n
MM3 CO1N A VSS VPW N12LL W=280.00n L=60.00n
.ENDS ACH2CONHSV1
****Sub-Circuit for ACH2CONHSV2, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT ACH2CONHSV2 A B CO0N CO1N VDD VSS
MM5 net50 B VDD VNW P12LL W=650.00n L=60.00n
MM4 CO1N A net50 VNW P12LL W=650.00n L=60.00n
MM13 CO0N B VDD VNW P12LL W=420.00n L=60.00n
MM12 CO0N A VDD VNW P12LL W=420.00n L=60.00n
MM11 CO0N A net83 VPW N12LL W=430.00n L=60.00n
MM10 net83 B VSS VPW N12LL W=430.00n L=60.00n
MM2 CO1N B VSS VPW N12LL W=350.00n L=60.00n
MM3 CO1N A VSS VPW N12LL W=350.00n L=60.00n
.ENDS ACH2CONHSV2
****Sub-Circuit for ACH2CONHSV4, Thu May 19 15:02:12 CST 2011****
.SUBCKT ACH2CONHSV4 A B CO0N CO1N VDD VSS
MM5 net50 B VDD VNW P12LL W=1.03u L=60.00n
MM4 CO1N A net50 VNW P12LL W=1.03u L=60.00n
MM13 CO0N B VDD VNW P12LL W=960.00n L=60.00n
MM12 CO0N A VDD VNW P12LL W=960.00n L=60.00n
MM11 CO0N A net83 VPW N12LL W=860n L=60.00n
MM10 net83 B VSS VPW N12LL W=860n L=60.00n
MM2 CO1N B VSS VPW N12LL W=700.00n L=60.00n
MM3 CO1N A VSS VPW N12LL W=700.00n L=60.00n
.ENDS ACH2CONHSV4
****Sub-Circuit for AD142HSV1, Thu May 19 13:57:40 CST 2011****
.SUBCKT AD142HSV1 A B C CI CO D ICO S VDD VSS
MM66 cin CI VSS VPW N12LL W=180.00n L=60.00n
MM65 cinn cin VSS VPW N12LL W=180.00n L=60.00n
MM61 cin xorabcd net0135 VPW N12LL W=180.00n L=60.00n
MM60 dn xnorabcd net0135 VPW N12LL W=180.00n L=60.00n
MM59 CO net0135 VSS VPW N12LL W=350.00n L=60.00n
MM57 S net0147 VSS VPW N12LL W=350.00n L=60.00n
MM54 cin xnorabcd net0147 VPW N12LL W=180.00n L=60.00n
MM53 cinn xorabcd net0147 VPW N12LL W=180.00n L=60.00n
MM52 xorab xnorab VSS VPW N12LL W=180.00n L=60.00n
MM49 xnorabcd xorabcd VSS VPW N12LL W=180.00n L=60.00n
MM47 xorabcd xnorab net0179 VPW N12LL W=180.00n L=60.00n
MM14 net0196 B VSS VPW N12LL W=210.00n L=60.00n
MM15 nandab A net0196 VPW N12LL W=210.00n L=60.00n
MM69 dn D VSS VPW N12LL W=180.00n L=60.00n
MM32 net0172 cn VSS VPW N12LL W=180.00n L=60.00n
MM26 net0204 A VSS VPW N12LL W=250.00n L=60.00n
MM29 net0204 B VSS VPW N12LL W=250.00n L=60.00n
MM31 xnorab nandab net0204 VPW N12LL W=180.00n L=60.00n
MM34 cn D net0179 VPW N12LL W=180.00n L=60.00n
MM27 cn C VSS VPW N12LL W=220.00n L=60.00n
MM33 net0172 dn net0179 VPW N12LL W=180.00n L=60.00n
MM19 ICO net108 VSS VPW N12LL W=350.00n L=60.00n
MM45 xorabcd net0179 xnorab VPW N12LL W=180.00n L=60.00n
MM36 nandab xnorab net108 VPW N12LL W=180.00n L=60.00n
MM38 cn xorab net108 VPW N12LL W=180.00n L=60.00n
MM68 cin CI VDD VNW P12LL W=220.00n L=60.00n
MM67 cinn cin VDD VNW P12LL W=220.00n L=60.00n
MM64 cin xnorabcd net0135 VNW P12LL W=220.00n L=60.00n
MM63 dn xorabcd net0135 VNW P12LL W=220.00n L=60.00n
MM62 CO net0135 VDD VNW P12LL W=440.00n L=60.00n
MM58 S net0147 VDD VNW P12LL W=440.00n L=60.00n
MM56 cin xorabcd net0147 VNW P12LL W=220.00n L=60.00n
MM55 cinn xnorabcd net0147 VNW P12LL W=220.00n L=60.00n
MM51 xorab xnorab VDD VNW P12LL W=220.00n L=60.00n
MM50 xnorabcd xorabcd VDD VNW P12LL W=220.00n L=60.00n
MM48 xorabcd xorab net0179 VNW P12LL W=220.00n L=60.00n
MM16 nandab A VDD VNW P12LL W=180.00n L=60.00n
MM17 nandab B VDD VNW P12LL W=180.00n L=60.00n
MM70 dn D VDD VNW P12LL W=220.00n L=60.00n
MM30 net0172 cn VDD VNW P12LL W=220.00n L=60.00n
MM18 xnorab A net0307 VNW P12LL W=200.00n L=60.00n
MM23 xnorab nandab VDD VNW P12LL W=200.00n L=60.00n
MM25 net0307 B VDD VNW P12LL W=200.00n L=60.00n
MM35 net0172 D net0179 VNW P12LL W=220.00n L=60.00n
MM37 cn dn net0179 VNW P12LL W=220.00n L=60.00n
MM28 cn C VDD VNW P12LL W=270.00n L=60.00n
MM20 ICO net108 VDD VNW P12LL W=440.00n L=60.00n
MM46 xorabcd net0179 xorab VNW P12LL W=220.00n L=60.00n
MM39 nandab xorab net108 VNW P12LL W=220.00n L=60.00n
MM40 cn xnorab net108 VNW P12LL W=220.00n L=60.00n
.ENDS AD142HSV1
****Sub-Circuit for AD142HSV2, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD142HSV2 A B C CI CO D ICO S VDD VSS
MM66 cin CI VSS VPW N12LL W=280.00n L=60.00n
MM65 cinn cin VSS VPW N12LL W=220.00n L=60.00n
MM61 cin xorabcd net0135 VPW N12LL W=220.00n L=60.00n
MM60 dn xnorabcd net0135 VPW N12LL W=220.00n L=60.00n
MM59 CO net0135 VSS VPW N12LL W=430.00n L=60.00n
MM57 S net0147 VSS VPW N12LL W=430.00n L=60.00n
MM54 cin xnorabcd net0147 VPW N12LL W=220.00n L=60.00n
MM53 cinn xorabcd net0147 VPW N12LL W=220.00n L=60.00n
MM52 xorab xnorab VSS VPW N12LL W=220.00n L=60.00n
MM49 xnorabcd xorabcd VSS VPW N12LL W=220.00n L=60.00n
MM47 xorabcd xnorab net0179 VPW N12LL W=220.00n L=60.00n
MM14 net0196 B VSS VPW N12LL W=430.00n L=60.00n
MM15 nandab A net0196 VPW N12LL W=430.00n L=60.00n
MM69 dn D VSS VPW N12LL W=280.00n L=60.00n
MM32 net0172 cn VSS VPW N12LL W=220.00n L=60.00n
MM26 net0204 A VSS VPW N12LL W=320.00n L=60.00n
MM29 net0204 B VSS VPW N12LL W=320.00n L=60.00n
MM31 xnorab nandab net0204 VPW N12LL W=180.00n L=60.00n
MM34 cn D net0179 VPW N12LL W=220.00n L=60.00n
MM27 cn C VSS VPW N12LL W=280.00n L=60.00n
MM33 net0172 dn net0179 VPW N12LL W=220.00n L=60.00n
MM19 ICO net108 VSS VPW N12LL W=430.00n L=60.00n
MM45 xorabcd net0179 xnorab VPW N12LL W=220.00n L=60.00n
MM36 nandab xnorab net108 VPW N12LL W=220.00n L=60.00n
MM38 cn xorab net108 VPW N12LL W=220.00n L=60.00n
MM68 cin CI VDD VNW P12LL W=350.00n L=60.00n
MM67 cinn cin VDD VNW P12LL W=270.00n L=60.00n
MM64 cin xnorabcd net0135 VNW P12LL W=270.00n L=60.00n
MM63 dn xorabcd net0135 VNW P12LL W=270.00n L=60.00n
MM62 CO net0135 VDD VNW P12LL W=540.00n L=60.00n
MM58 S net0147 VDD VNW P12LL W=540.00n L=60.00n
MM56 cin xorabcd net0147 VNW P12LL W=270.00n L=60.00n
MM55 cinn xnorabcd net0147 VNW P12LL W=270.00n L=60.00n
MM51 xorab xnorab VDD VNW P12LL W=270.00n L=60.00n
MM50 xnorabcd xorabcd VDD VNW P12LL W=270.00n L=60.00n
MM48 xorabcd xorab net0179 VNW P12LL W=270.00n L=60.00n
MM16 nandab A VDD VNW P12LL W=420.00n L=60.00n
MM17 nandab B VDD VNW P12LL W=420.00n L=60.00n
MM70 dn D VDD VNW P12LL W=350.00n L=60.00n
MM30 net0172 cn VDD VNW P12LL W=270.00n L=60.00n
MM18 xnorab A net0307 VNW P12LL W=220.00n L=60.00n
MM23 xnorab nandab VDD VNW P12LL W=220.00n L=60.00n
MM25 net0307 B VDD VNW P12LL W=220.00n L=60.00n
MM35 net0172 D net0179 VNW P12LL W=270.00n L=60.00n
MM37 cn dn net0179 VNW P12LL W=270.00n L=60.00n
MM28 cn C VDD VNW P12LL W=350.00n L=60.00n
MM20 ICO net108 VDD VNW P12LL W=540.00n L=60.00n
MM46 xorabcd net0179 xorab VNW P12LL W=270.00n L=60.00n
MM39 nandab xorab net108 VNW P12LL W=270.00n L=60.00n
MM40 cn xnorab net108 VNW P12LL W=270.00n L=60.00n
.ENDS AD142HSV2
****Sub-Circuit for AD142HSV4, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD142HSV4 A B C CI CO D ICO S VDD VSS
MM66 cin CI VSS VPW N12LL W=430.00n L=60.00n
MM65 cinn cin VSS VPW N12LL W=350.00n L=60.00n
MM61 cin xorabcd net0135 VPW N12LL W=430.00n L=60.00n
MM60 dn xnorabcd net0135 VPW N12LL W=430.00n L=60.00n
MM59 CO net0135 VSS VPW N12LL W=860.00n L=60.00n
MM57 S net0147 VSS VPW N12LL W=860.00n L=60.00n
MM54 cin xnorabcd net0147 VPW N12LL W=430.00n L=60.00n
MM53 cinn xorabcd net0147 VPW N12LL W=430.00n L=60.00n
MM52 xorab xnorab VSS VPW N12LL W=430.00n L=60.00n
MM49 xnorabcd xorabcd VSS VPW N12LL W=430.00n L=60.00n
MM47 xorabcd xnorab net0179 VPW N12LL W=430.00n L=60.00n
MM14 net0196 B VSS VPW N12LL W=430.00n L=60.00n
MM15 nandab A net0196 VPW N12LL W=430.00n L=60.00n
MM69 dn D VSS VPW N12LL W=430.00n L=60.00n
MM32 net0172 cn VSS VPW N12LL W=430.00n L=60.00n
MM26 net0204 A VSS VPW N12LL W=320.00n L=60.00n
MM29 net0204 B VSS VPW N12LL W=320.00n L=60.00n
MM31 xnorab nandab net0204 VPW N12LL W=180.00n L=60.00n
MM34 cn D net0179 VPW N12LL W=430.00n L=60.00n
MM27 cn C VSS VPW N12LL W=430.00n L=60.00n
MM33 net0172 dn net0179 VPW N12LL W=430.00n L=60.00n
MM19 ICO net108 VSS VPW N12LL W=860.00n L=60.00n
MM45 xorabcd net0179 xnorab VPW N12LL W=430.00n L=60.00n
MM36 nandab xnorab net108 VPW N12LL W=430.00n L=60.00n
MM38 cn xorab net108 VPW N12LL W=430.00n L=60.00n
MM68 cin CI VDD VNW P12LL W=540.00n L=60.00n
MM67 cinn cin VDD VNW P12LL W=440.00n L=60.00n
MM64 cin xnorabcd net0135 VNW P12LL W=540.00n L=60.00n
MM63 dn xorabcd net0135 VNW P12LL W=540.00n L=60.00n
MM62 CO net0135 VDD VNW P12LL W=1.08u L=60.00n
MM58 S net0147 VDD VNW P12LL W=1.08u L=60.00n
MM56 cin xorabcd net0147 VNW P12LL W=540.00n L=60.00n
MM55 cinn xnorabcd net0147 VNW P12LL W=540.00n L=60.00n
MM51 xorab xnorab VDD VNW P12LL W=540.00n L=60.00n
MM50 xnorabcd xorabcd VDD VNW P12LL W=540.00n L=60.00n
MM48 xorabcd xorab net0179 VNW P12LL W=540.00n L=60.00n
MM16 nandab A VDD VNW P12LL W=420.00n L=60.00n
MM17 nandab B VDD VNW P12LL W=420.00n L=60.00n
MM70 dn D VDD VNW P12LL W=540.00n L=60.00n
MM30 net0172 cn VDD VNW P12LL W=540.00n L=60.00n
MM18 xnorab A net0307 VNW P12LL W=220.00n L=60.00n
MM23 xnorab nandab VDD VNW P12LL W=220.00n L=60.00n
MM25 net0307 B VDD VNW P12LL W=220.00n L=60.00n
MM35 net0172 D net0179 VNW P12LL W=540.00n L=60.00n
MM37 cn dn net0179 VNW P12LL W=540.00n L=60.00n
MM28 cn C VDD VNW P12LL W=540.00n L=60.00n
MM20 ICO net108 VDD VNW P12LL W=1.08u L=60.00n
MM46 xorabcd net0179 xorab VNW P12LL W=540.00n L=60.00n
MM39 nandab xorab net108 VNW P12LL W=540.00n L=60.00n
MM40 cn xnorab net108 VNW P12LL W=540.00n L=60.00n
.ENDS AD142HSV4
****Sub-Circuit for AD1CINHSV1, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1CINHSV1 A B CIN CO S VDD VSS
MM41 net0196 CIN net78 VPW N12LL W=180.00n L=60.00n
MM42 norab cinn net78 VPW N12LL W=180.00n L=60.00n
MMN1 xo norab VSS VPW N12LL W=390.00n L=60.00n
MM3 norab A VSS VPW N12LL W=300.00n L=60.00n
MM0 xo A net0164 VPW N12LL W=440.00n L=60.00n
MM2 norab B VSS VPW N12LL W=300.00n L=60.00n
MM7 net0164 B VSS VPW N12LL W=440.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=180.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=210.00n L=60.00n
MM11 net0196 A net0124 VPW N12LL W=210.00n L=60.00n
MM27 cinn CIN VSS VPW N12LL W=180.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=350.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=350.00n L=60.00n
MM36 xn CIN net108 VPW N12LL W=180.00n L=60.00n
MM38 xo cinn net108 VPW N12LL W=180.00n L=60.00n
MM43 net0196 cinn net78 VNW P12LL W=220.00n L=60.00n
MM44 norab CIN net78 VNW P12LL W=220.00n L=60.00n
MM12 net0196 A VDD VNW P12LL W=180.00n L=60.00n
MM13 net0196 B VDD VNW P12LL W=180.00n L=60.00n
MM28 cinn CIN VDD VNW P12LL W=220.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=440.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=440.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=550.00n L=60.00n
MMP1 net0223 A VDD VNW P12LL W=550.00n L=60.00n
MM1 xo norab net0223 VNW P12LL W=440.00n L=60.00n
MM6 net0223 B VDD VNW P12LL W=550.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=550.00n L=60.00n
MM9 xn xo VDD VNW P12LL W=220.00n L=60.00n
MM39 xn cinn net108 VNW P12LL W=220.00n L=60.00n
MM40 xo CIN net108 VNW P12LL W=220.00n L=60.00n
.ENDS AD1CINHSV1
****Sub-Circuit for AD1CINHSV2, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1CINHSV2 A B CIN CO S VDD VSS
MM41 net0196 CIN net78 VPW N12LL W=220.00n L=60.00n
MM42 norab cinn net78 VPW N12LL W=220.00n L=60.00n
MMN1 xo norab VSS VPW N12LL W=430.00n L=60.00n
MM3 norab A VSS VPW N12LL W=350.00n L=60.00n
MM0 xo A net0164 VPW N12LL W=430.00n L=60.00n
MM2 norab B VSS VPW N12LL W=350.00n L=60.00n
MM7 net0164 B VSS VPW N12LL W=430.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=220.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=260.00n L=60.00n
MM11 net0196 A net0124 VPW N12LL W=260.00n L=60.00n
MM27 cinn CIN VSS VPW N12LL W=220.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=430.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=430.00n L=60.00n
MM36 xn CIN net108 VPW N12LL W=220.00n L=60.00n
MM38 xo cinn net108 VPW N12LL W=220.00n L=60.00n
MM43 net0196 cinn net78 VNW P12LL W=270.00n L=60.00n
MM44 norab CIN net78 VNW P12LL W=270.00n L=60.00n
MM12 net0196 A VDD VNW P12LL W=220.00n L=60.00n
MM13 net0196 B VDD VNW P12LL W=220.00n L=60.00n
MM28 cinn CIN VDD VNW P12LL W=270.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=540.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=540.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=650.00n L=60.00n
MMP1 net0223 A VDD VNW P12LL W=650.00n L=60.00n
MM1 xo norab net0223 VNW P12LL W=540.00n L=60.00n
MM6 net0223 B VDD VNW P12LL W=650.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=650.00n L=60.00n
MM9 xn xo VDD VNW P12LL W=270.00n L=60.00n
MM39 xn cinn net108 VNW P12LL W=270.00n L=60.00n
MM40 xo CIN net108 VNW P12LL W=270.00n L=60.00n
.ENDS AD1CINHSV2
****Sub-Circuit for AD1CINHSV4, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1CINHSV4 A B CIN CO S VDD VSS
MM41 net0196 CIN net78 VPW N12LL W=430.00n L=60.00n
MM42 norab cinn net78 VPW N12LL W=430.00n L=60.00n
MMN1 xo norab VSS VPW N12LL W=880.00n L=60.00n
MM3 norab A VSS VPW N12LL W=700.00n L=60.00n
MM0 xo A net0164 VPW N12LL W=1.08u L=60.00n
MM2 norab B VSS VPW N12LL W=700.00n L=60.00n
MM7 net0164 B VSS VPW N12LL W=1.08u L=60.00n
MM8 xn xo VSS VPW N12LL W=430.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=520.00n L=60.00n
MM11 net0196 A net0124 VPW N12LL W=520.00n L=60.00n
MM27 cinn CIN VSS VPW N12LL W=220.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=860.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=860.00n L=60.00n
MM36 xn CIN net108 VPW N12LL W=430.00n L=60.00n
MM38 xo cinn net108 VPW N12LL W=430.00n L=60.00n
MM43 net0196 cinn net78 VNW P12LL W=540.00n L=60.00n
MM44 norab CIN net78 VNW P12LL W=540.00n L=60.00n
MM12 net0196 A VDD VNW P12LL W=440.00n L=60.00n
MM13 net0196 B VDD VNW P12LL W=440.00n L=60.00n
MM28 cinn CIN VDD VNW P12LL W=270.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=1.08u L=60.00n
MM20 S net108 VDD VNW P12LL W=1.08u L=60.00n
MM4 norab A net0215 VNW P12LL W=1.3u L=60.00n
MMP1 net0223 A VDD VNW P12LL W=1.3u L=60.00n
MM1 xo norab net0223 VNW P12LL W=1.08u L=60.00n
MM6 net0223 B VDD VNW P12LL W=1.3u L=60.00n
MM5 net0215 B VDD VNW P12LL W=1.3u L=60.00n
MM9 xn xo VDD VNW P12LL W=540.00n L=60.00n
MM39 xn cinn net108 VNW P12LL W=540.00n L=60.00n
MM40 xo CIN net108 VNW P12LL W=540.00n L=60.00n
.ENDS AD1CINHSV4
****Sub-Circuit for AD1CONHSV1, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1CONHSV1 A B CI CON S VDD VSS
MM16 net0133 norab VSS VPW N12LL W=180.00n L=60.00n
MM41 net0196 cin net78 VPW N12LL W=180.00n L=60.00n
MM42 net0133 CI net78 VPW N12LL W=180.00n L=60.00n
MMN1 xo norab VSS VPW N12LL W=390.00n L=60.00n
MM3 norab A VSS VPW N12LL W=300.00n L=60.00n
MM0 xo A net0164 VPW N12LL W=440.00n L=60.00n
MM2 norab B VSS VPW N12LL W=300.00n L=60.00n
MM7 net0164 B VSS VPW N12LL W=440.00n L=60.00n
MM14 net0196 net0193 VSS VPW N12LL W=180.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=180.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=210.00n L=60.00n
MM11 net0193 A net0124 VPW N12LL W=210.00n L=60.00n
MM27 cin CI VSS VPW N12LL W=180.00n L=60.00n
MM22 CON net78 VSS VPW N12LL W=350.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=350.00n L=60.00n
MM36 xn cin net108 VPW N12LL W=180.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=180.00n L=60.00n
MM17 net0133 norab VDD VNW P12LL W=220.00n L=60.00n
MM43 net0196 CI net78 VNW P12LL W=220.00n L=60.00n
MM44 net0133 cin net78 VNW P12LL W=220.00n L=60.00n
MM15 net0196 net0193 VDD VNW P12LL W=220.00n L=60.00n
MM12 net0193 A VDD VNW P12LL W=180.00n L=60.00n
MM13 net0193 B VDD VNW P12LL W=180.00n L=60.00n
MM28 cin CI VDD VNW P12LL W=220.00n L=60.00n
MM21 CON net78 VDD VNW P12LL W=440.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=440.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=550.00n L=60.00n
MMP1 net0223 A VDD VNW P12LL W=550.00n L=60.00n
MM1 xo norab net0223 VNW P12LL W=440.00n L=60.00n
MM6 net0223 B VDD VNW P12LL W=550.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=550.00n L=60.00n
MM9 xn xo VDD VNW P12LL W=220.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=220.00n L=60.00n
MM40 xo cin net108 VNW P12LL W=220.00n L=60.00n
.ENDS AD1CONHSV1
****Sub-Circuit for AD1CONHSV2, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1CONHSV2 A B CI CON S VDD VSS
MM17 net0133 norab VSS VPW N12LL W=220.00n L=60.00n
MM41 net0196 cin net78 VPW N12LL W=220.00n L=60.00n
MM42 net0133 CI net78 VPW N12LL W=220.00n L=60.00n
MMN1 xo norab VSS VPW N12LL W=430.00n L=60.00n
MM3 norab A VSS VPW N12LL W=350.00n L=60.00n
MM0 xo A net0164 VPW N12LL W=430.00n L=60.00n
MM2 norab B VSS VPW N12LL W=350.00n L=60.00n
MM7 net0164 B VSS VPW N12LL W=430.00n L=60.00n
MM14 net0196 net0193 VSS VPW N12LL W=220.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=220.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=260.00n L=60.00n
MM11 net0193 A net0124 VPW N12LL W=260.00n L=60.00n
MM27 cin CI VSS VPW N12LL W=220.00n L=60.00n
MM22 CON net78 VSS VPW N12LL W=430.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=430.00n L=60.00n
MM36 xn cin net108 VPW N12LL W=220.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=220.00n L=60.00n
MM16 net0133 norab VDD VNW P12LL W=270.00n L=60.00n
MM43 net0196 CI net78 VNW P12LL W=270.00n L=60.00n
MM44 net0133 cin net78 VNW P12LL W=270.00n L=60.00n
MM15 net0196 net0193 VDD VNW P12LL W=270.00n L=60.00n
MM12 net0193 A VDD VNW P12LL W=220.00n L=60.00n
MM13 net0193 B VDD VNW P12LL W=220.00n L=60.00n
MM28 cin CI VDD VNW P12LL W=270.00n L=60.00n
MM21 CON net78 VDD VNW P12LL W=540.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=540.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=650.00n L=60.00n
MMP1 net0223 A VDD VNW P12LL W=650.00n L=60.00n
MM1 xo norab net0223 VNW P12LL W=540.00n L=60.00n
MM6 net0223 B VDD VNW P12LL W=650.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=650.00n L=60.00n
MM9 xn xo VDD VNW P12LL W=270.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=270.00n L=60.00n
MM40 xo cin net108 VNW P12LL W=270.00n L=60.00n
.ENDS AD1CONHSV2
****Sub-Circuit for AD1CONHSV4, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1CONHSV4 A B CI CON S VDD VSS
MM41 net0196 cin net78 VPW N12LL W=430.00n L=60.00n
MM42 net0141 CI net78 VPW N12LL W=430.00n L=60.00n
MM17 net0141 norab VSS VPW N12LL W=430.00n L=60.00n
MMN1 xo norab VSS VPW N12LL W=880.00n L=60.00n
MM3 norab A VSS VPW N12LL W=700.00n L=60.00n
MM0 xo A net0164 VPW N12LL W=0.86u L=60.00n
MM2 norab B VSS VPW N12LL W=700.00n L=60.00n
MM7 net0164 B VSS VPW N12LL W=0.86u L=60.00n
MM14 net0196 net0193 VSS VPW N12LL W=430.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=430.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=430.00n L=60.00n
MM11 net0193 A net0124 VPW N12LL W=430.00n L=60.00n
MM27 cin CI VSS VPW N12LL W=220.00n L=60.00n
MM22 CON net78 VSS VPW N12LL W=860.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=860.00n L=60.00n
MM36 xn cin net108 VPW N12LL W=430.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=430.00n L=60.00n
MM16 net0141 norab VDD VNW P12LL W=540.00n L=60.00n
MM43 net0196 CI net78 VNW P12LL W=540.00n L=60.00n
MM44 net0141 cin net78 VNW P12LL W=540.00n L=60.00n
MM15 net0196 net0193 VDD VNW P12LL W=540.00n L=60.00n
MM12 net0193 A VDD VNW P12LL W=540.00n L=60.00n
MM13 net0193 B VDD VNW P12LL W=540.00n L=60.00n
MM28 cin CI VDD VNW P12LL W=270.00n L=60.00n
MM21 CON net78 VDD VNW P12LL W=1.08u L=60.00n
MM20 S net108 VDD VNW P12LL W=1.08u L=60.00n
MM4 norab A net0215 VNW P12LL W=1.3u L=60.00n
MMP1 net0223 A VDD VNW P12LL W=1.3u L=60.00n
MM1 xo norab net0223 VNW P12LL W=1.08u L=60.00n
MM6 net0223 B VDD VNW P12LL W=1.3u L=60.00n
MM5 net0215 B VDD VNW P12LL W=1.3u L=60.00n
MM9 xn xo VDD VNW P12LL W=540.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=540.00n L=60.00n
MM40 xo cin net108 VNW P12LL W=540.00n L=60.00n
.ENDS AD1CONHSV4
****Sub-Circuit for AD1HSV1, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AD1HSV1 A B CI CO S VDD VSS
MM41 net115 xo net78 VPW N12LL W=260.00n L=60.00n
MM42 net117 xn net78 VPW N12LL W=260.00n L=60.00n
MM31 net115 CI VSS VPW N12LL W=300.00n L=60.00n
MM30 net109 net117 VSS VPW N12LL W=340.00n L=60.00n
MM27 net117 B VSS VPW N12LL W=260.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=300.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=300.00n L=60.00n
MM17 net119 A VSS VPW N12LL W=400.00n L=60.00n
MM36 xn net115 net108 VPW N12LL W=260.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=260.00n L=60.00n
MM3 xn net117 net119 VPW N12LL W=260.00n L=60.00n
MM35 xo net119 net109 VPW N12LL W=260.00n L=60.00n
MM5 xo net109 net119 VPW N12LL W=260.00n L=60.00n
MM0 xn net119 net117 VPW N12LL W=240.00n L=60.00n
MM43 net115 xn net78 VNW P12LL W=400.00n L=60.00n
MM44 net117 xo net78 VNW P12LL W=400.00n L=60.00n
MM32 net115 CI VDD VNW P12LL W=450.00n L=60.00n
MM29 net109 net117 VDD VNW P12LL W=500.00n L=60.00n
MM28 net117 B VDD VNW P12LL W=400.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=450.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=450.00n L=60.00n
MM18 net119 A VDD VNW P12LL W=600.00n L=60.00n
MM37 xo net119 net117 VNW P12LL W=400.00n L=60.00n
MM4 xn net109 net119 VNW P12LL W=400.00n L=60.00n
MM6 xo net117 net119 VNW P12LL W=400.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=400.00n L=60.00n
MM40 xo net115 net108 VNW P12LL W=400.00n L=60.00n
MM1 xn net119 net109 VNW P12LL W=375.00n L=60.00n
.ENDS AD1HSV1
****Sub-Circuit for AD1HSV1C, Thu May 19 13:57:40 CST 2011****
.SUBCKT AD1HSV1C A B CI CO S VDD VSS
MM16 net0152 B VSS VPW N12LL W=250.00n L=60.00n
MM13 net0164 B VSS VPW N12LL W=180.00n L=60.00n
MM5 net100 CI net0144 VPW N12LL W=180.00n L=60.00n
MM39 net108 CI net0168 VPW N12LL W=180.00n L=60.00n
MM38 net108 net100 net0152 VPW N12LL W=180.00n L=60.00n
MM15 net0152 A VSS VPW N12LL W=250.00n L=60.00n
MM4 net0144 B VSS VPW N12LL W=250.00n L=60.00n
MM31 CO net100 VSS VPW N12LL W=350.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=350.00n L=60.00n
MM17 net100 A net0140 VPW N12LL W=180.00n L=60.00n
MM36 net0168 A net0164 VPW N12LL W=180.00n L=60.00n
MM37 net0140 B VSS VPW N12LL W=180.00n L=60.00n
MM14 net0152 CI VSS VPW N12LL W=250.00n L=60.00n
MM35 net0144 A VSS VPW N12LL W=250.00n L=60.00n
MM8 net108 CI net0227 VNW P12LL W=200.00n L=60.00n
MM7 net0231 B VDD VNW P12LL W=200.00n L=60.00n
MM6 net0227 A net0231 VNW P12LL W=200.00n L=60.00n
MM10 net0212 B VDD VNW P12LL W=290.00n L=60.00n
MM11 net0212 CI VDD VNW P12LL W=290.00n L=60.00n
MM2 net100 A net0183 VNW P12LL W=200.00n L=60.00n
MM3 net0183 B VDD VNW P12LL W=200.00n L=60.00n
MM32 CO net100 VDD VNW P12LL W=440.00n L=60.00n
MM12 net108 net100 net0212 VNW P12LL W=200.00n L=60.00n
MM9 net0212 A VDD VNW P12LL W=290.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=440.00n L=60.00n
MM18 net0203 A VDD VNW P12LL W=290.00n L=60.00n
MM1 net0203 B VDD VNW P12LL W=290.00n L=60.00n
MM0 net100 CI net0203 VNW P12LL W=200.00n L=60.00n
.ENDS AD1HSV1C
****Sub-Circuit for AD1HSV1R, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1HSV1R A B CI CO S VDD VSS
MM41 net0196 cin net78 VPW N12LL W=180.00n L=60.00n
MM42 norab CI net78 VPW N12LL W=180.00n L=60.00n
MMN1 xo norab VSS VPW N12LL W=390.00n L=60.00n
MM3 norab A VSS VPW N12LL W=300.00n L=60.00n
MM0 xo A net0164 VPW N12LL W=430.00n L=60.00n
MM2 norab B VSS VPW N12LL W=300.00n L=60.00n
MM7 net0164 B VSS VPW N12LL W=430.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=180.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=210.00n L=60.00n
MM11 net0196 A net0124 VPW N12LL W=210.00n L=60.00n
MM27 cin CI VSS VPW N12LL W=180.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=350.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=350.00n L=60.00n
MM36 xn cin net108 VPW N12LL W=180.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=180.00n L=60.00n
MM43 net0196 CI net78 VNW P12LL W=220.00n L=60.00n
MM44 norab cin net78 VNW P12LL W=220.00n L=60.00n
MM12 net0196 A VDD VNW P12LL W=180.00n L=60.00n
MM13 net0196 B VDD VNW P12LL W=180.00n L=60.00n
MM28 cin CI VDD VNW P12LL W=220.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=440.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=440.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=550.00n L=60.00n
MMP1 net0223 A VDD VNW P12LL W=550.00n L=60.00n
MM1 xo norab net0223 VNW P12LL W=440.00n L=60.00n
MM6 net0223 B VDD VNW P12LL W=550.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=550.00n L=60.00n
MM9 xn xo VDD VNW P12LL W=220.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=220.00n L=60.00n
MM40 xo cin net108 VNW P12LL W=220.00n L=60.00n
.ENDS AD1HSV1R
****Sub-Circuit for AD1HSV1T, Mon May 30 15:56:35 CST 2011****
.SUBCKT AD1HSV1T A B CI CO S VDD VSS
MM10 net117 B VSS VPW N12LL W=350.00n L=60.00n
MM41 cin xo net78 VPW N12LL W=180.00n L=60.00n
MM42 net117 xn net78 VPW N12LL W=180.00n L=60.00n
MMN1 xo net0164 VSS VPW N12LL W=290.00n L=60.00n
MM2 net0164 B VSS VPW N12LL W=290.00n L=60.00n
MM3 net0164 A VSS VPW N12LL W=290.00n L=60.00n
MM0 xo A net0176 VPW N12LL W=350.00n L=60.00n
MM7 net0176 B VSS VPW N12LL W=350.00n L=60.00n
MM31 cin CI VSS VPW N12LL W=350.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=360.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=350.00n L=60.00n
MM36 xn cin net108 VPW N12LL W=180.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=180.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=180.00n L=60.00n
MM11 net117 B VDD VNW P12LL W=440.00n L=60.00n
MM43 cin xn net78 VNW P12LL W=220.00n L=60.00n
MM44 net117 xo net78 VNW P12LL W=220.00n L=60.00n
MM4 net0164 A net0235 VNW P12LL W=540.00n L=60.00n
MMP1 net0227 A VDD VNW P12LL W=590.00n L=60.00n
MM1 xo net0164 net0227 VNW P12LL W=440.00n L=60.00n
MM6 net0227 B VDD VNW P12LL W=590.00n L=60.00n
MM5 net0235 B VDD VNW P12LL W=540.00n L=60.00n
MM32 cin CI VDD VNW P12LL W=440.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=440n L=60.00n
MM20 S net108 VDD VNW P12LL W=440n L=60.00n
MM9 xn xo VDD VNW P12LL W=220.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=220.00n L=60.00n
MM40 xo cin net108 VNW P12LL W=220.00n L=60.00n
.ENDS AD1HSV1T
****Sub-Circuit for AD1HSV2, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AD1HSV2 A B CI CO S VDD VSS
MM41 net115 xo net78 VPW N12LL W=380.00n L=60.00n
MM42 net117 xn net78 VPW N12LL W=380.00n L=60.00n
MM31 net115 CI VSS VPW N12LL W=430.00n L=60.00n
MM30 net109 net117 VSS VPW N12LL W=510.00n L=60.00n
MM27 net117 B VSS VPW N12LL W=390.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=430.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=430.00n L=60.00n
MM17 net119 A VSS VPW N12LL W=600.00n L=60.00n
MM36 xn net115 net108 VPW N12LL W=380.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=380.00n L=60.00n
MM3 xn net117 net119 VPW N12LL W=500.00n L=60.00n
MM35 xo net119 net109 VPW N12LL W=500.00n L=60.00n
MM5 xo net109 net119 VPW N12LL W=500.00n L=60.00n
MM0 xn net119 net117 VPW N12LL W=500.00n L=60.00n
MM43 net115 xn net78 VNW P12LL W=580.00n L=60.00n
MM44 net117 xo net78 VNW P12LL W=580.00n L=60.00n
MM32 net115 CI VDD VNW P12LL W=650.00n L=60.00n
MM29 net109 net117 VDD VNW P12LL W=760.00n L=60.00n
MM28 net117 B VDD VNW P12LL W=600.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=650.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=650.00n L=60.00n
MM18 net119 A VDD VNW P12LL W=920.00n L=60.00n
MM37 xo net119 net117 VNW P12LL W=780.00n L=60.00n
MM4 xn net109 net119 VNW P12LL W=780.00n L=60.00n
MM6 xo net117 net119 VNW P12LL W=780.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=580.00n L=60.00n
MM40 xo net115 net108 VNW P12LL W=580.00n L=60.00n
MM1 xn net119 net109 VNW P12LL W=780.00n L=60.00n
.ENDS AD1HSV2
****Sub-Circuit for AD1HSV2C, Thu May 19 14:42:46 CST 2011****
.SUBCKT AD1HSV2C A B CI CO S VDD VSS
MM16 net0152 B VSS VPW N12LL W=320.00n L=60.00n
MM13 net0164 B VSS VPW N12LL W=180.00n L=60.00n
MM5 net100 CI net0144 VPW N12LL W=180.00n L=60.00n
MM39 net108 CI net0168 VPW N12LL W=180.00n L=60.00n
MM38 net108 net100 net0152 VPW N12LL W=180.00n L=60.00n
MM15 net0152 A VSS VPW N12LL W=320.00n L=60.00n
MM4 net0144 B VSS VPW N12LL W=320.00n L=60.00n
MM31 CO net100 VSS VPW N12LL W=430.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=430.00n L=60.00n
MM17 net100 A net0140 VPW N12LL W=180.00n L=60.00n
MM36 net0168 A net0164 VPW N12LL W=180.00n L=60.00n
MM37 net0140 B VSS VPW N12LL W=180.00n L=60.00n
MM14 net0152 CI VSS VPW N12LL W=320.00n L=60.00n
MM35 net0144 A VSS VPW N12LL W=320.00n L=60.00n
MM8 net108 CI net0227 VNW P12LL W=220.00n L=60.00n
MM7 net0231 B VDD VNW P12LL W=220.00n L=60.00n
MM6 net0227 A net0231 VNW P12LL W=220.00n L=60.00n
MM10 net0212 B VDD VNW P12LL W=350.00n L=60.00n
MM11 net0212 CI VDD VNW P12LL W=325.00n L=60.00n
MM2 net100 A net0183 VNW P12LL W=220.00n L=60.00n
MM3 net0183 B VDD VNW P12LL W=220.00n L=60.00n
MM32 CO net100 VDD VNW P12LL W=540.00n L=60.00n
MM12 net108 net100 net0212 VNW P12LL W=220.00n L=60.00n
MM9 net0212 A VDD VNW P12LL W=350.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=540.00n L=60.00n
MM18 net0203 A VDD VNW P12LL W=350.00n L=60.00n
MM1 net0203 B VDD VNW P12LL W=350.00n L=60.00n
MM0 net100 CI net0203 VNW P12LL W=220.00n L=60.00n
.ENDS AD1HSV2C
****Sub-Circuit for AD1HSV2R, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1HSV2R A B CI CO S VDD VSS
MM41 net0196 cin net78 VPW N12LL W=220.00n L=60.00n
MM42 norab CI net78 VPW N12LL W=220.00n L=60.00n
MMN1 xo norab VSS VPW N12LL W=430.00n L=60.00n
MM3 norab A VSS VPW N12LL W=350.00n L=60.00n
MM0 xo A net0164 VPW N12LL W=430.00n L=60.00n
MM2 norab B VSS VPW N12LL W=350.00n L=60.00n
MM7 net0164 B VSS VPW N12LL W=430.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=220.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=260.00n L=60.00n
MM11 net0196 A net0124 VPW N12LL W=260.00n L=60.00n
MM27 cin CI VSS VPW N12LL W=220.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=430.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=430.00n L=60.00n
MM36 xn cin net108 VPW N12LL W=220.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=220.00n L=60.00n
MM43 net0196 CI net78 VNW P12LL W=270.00n L=60.00n
MM44 norab cin net78 VNW P12LL W=270.00n L=60.00n
MM12 net0196 A VDD VNW P12LL W=220.00n L=60.00n
MM13 net0196 B VDD VNW P12LL W=220.00n L=60.00n
MM28 cin CI VDD VNW P12LL W=270.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=540.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=540.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=650.00n L=60.00n
MMP1 net0223 A VDD VNW P12LL W=650.00n L=60.00n
MM1 xo norab net0223 VNW P12LL W=540.00n L=60.00n
MM6 net0223 B VDD VNW P12LL W=650.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=650.00n L=60.00n
MM9 xn xo VDD VNW P12LL W=270.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=270.00n L=60.00n
MM40 xo cin net108 VNW P12LL W=270.00n L=60.00n
.ENDS AD1HSV2R
****Sub-Circuit for AD1HSV2T, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1HSV2T A B CI CO S VDD VSS
MM10 net117 B VSS VPW N12LL W=430.00n L=60.00n
MM41 cin xo net78 VPW N12LL W=220.00n L=60.00n
MM42 net117 xn net78 VPW N12LL W=220.00n L=60.00n
MMN1 xo net0164 VSS VPW N12LL W=350.00n L=60.00n
MM2 net0164 B VSS VPW N12LL W=350.00n L=60.00n
MM3 net0164 A VSS VPW N12LL W=350.00n L=60.00n
MM0 xo A net0176 VPW N12LL W=430.00n L=60.00n
MM7 net0176 B VSS VPW N12LL W=430.00n L=60.00n
MM31 cin CI VSS VPW N12LL W=430.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=430.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=430.00n L=60.00n
MM36 xn cin net108 VPW N12LL W=220.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=220.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=220.00n L=60.00n
MM11 net117 B VDD VNW P12LL W=540.00n L=60.00n
MM43 cin xn net78 VNW P12LL W=270.00n L=60.00n
MM44 net117 xo net78 VNW P12LL W=270.00n L=60.00n
MM4 net0164 A net0235 VNW P12LL W=650.00n L=60.00n
MMP1 net0227 A VDD VNW P12LL W=650.00n L=60.00n
MM1 xo net0164 net0227 VNW P12LL W=540.00n L=60.00n
MM6 net0227 B VDD VNW P12LL W=650.00n L=60.00n
MM5 net0235 B VDD VNW P12LL W=650.00n L=60.00n
MM32 cin CI VDD VNW P12LL W=540.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=540.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=540.00n L=60.00n
MM9 xn xo VDD VNW P12LL W=270.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=270.00n L=60.00n
MM40 xo cin net108 VNW P12LL W=270.00n L=60.00n
.ENDS AD1HSV2T
****Sub-Circuit for AD1HSV4, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AD1HSV4 A B CI CO S VDD VSS
MM41 net115 xo net78 VPW N12LL W=780.00n L=60.00n
MM42 net117 xn net78 VPW N12LL W=780.00n L=60.00n
MM31 net115 CI VSS VPW N12LL W=860.00n L=60.00n
MM30 net109 net117 VSS VPW N12LL W=960.00n L=60.00n
MM27 net117 B VSS VPW N12LL W=860.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=860.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=860.00n L=60.00n
MM17 net119 A VSS VPW N12LL W=860.00n L=60.00n
MM36 xn net115 net108 VPW N12LL W=780.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=780.00n L=60.00n
MM3 xn net117 net119 VPW N12LL W=780.00n L=60.00n
MM35 xo net119 net109 VPW N12LL W=780.00n L=60.00n
MM5 xo net109 net119 VPW N12LL W=780.00n L=60.00n
MM0 xn net119 net117 VPW N12LL W=780.00n L=60.00n
MM43 net115 xn net78 VNW P12LL W=1.2u L=60.00n
MM44 net117 xo net78 VNW P12LL W=1.2u L=60.00n
MM32 net115 CI VDD VNW P12LL W=1.3u L=60.00n
MM29 net109 net117 VDD VNW P12LL W=1.41u L=60.00n
MM28 net117 B VDD VNW P12LL W=1.3u L=60.00n
MM21 CO net78 VDD VNW P12LL W=1.3u L=60.00n
MM20 S net108 VDD VNW P12LL W=1.3u L=60.00n
MM18 net119 A VDD VNW P12LL W=1.3u L=60.00n
MM37 xo net119 net117 VNW P12LL W=1.18u L=60.00n
MM4 xn net109 net119 VNW P12LL W=1.18u L=60.00n
MM6 xo net117 net119 VNW P12LL W=1.18u L=60.00n
MM39 xn CI net108 VNW P12LL W=1.2u L=60.00n
MM40 xo net115 net108 VNW P12LL W=1.2u L=60.00n
MM1 xn net119 net109 VNW P12LL W=1.18u L=60.00n
.ENDS AD1HSV4
****Sub-Circuit for AD1HSV4C, Tue May 24 14:57:30 CST 2011****
.SUBCKT AD1HSV4C A B CI CO S VDD VSS
MM16 net0152 B VSS VPW N12LL W=430.00n L=60.00n
MM13 net0164 B VSS VPW N12LL W=300.00n L=60.00n
MM5 net100 CI net0144 VPW N12LL W=350.00n L=60.00n
MM39 net108 CI net0168 VPW N12LL W=300.00n L=60.00n
MM38 net108 net100 net0152 VPW N12LL W=300.00n L=60.00n
MM15 net0152 A VSS VPW N12LL W=430.00n L=60.00n
MM4 net0144 B VSS VPW N12LL W=430.00n L=60.00n
MM31 CO net100 VSS VPW N12LL W=860.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=860.00n L=60.00n
MM17 net100 A net0140 VPW N12LL W=350.00n L=60.00n
MM36 net0168 A net0164 VPW N12LL W=300.00n L=60.00n
MM37 net0140 B VSS VPW N12LL W=350.00n L=60.00n
MM14 net0152 CI VSS VPW N12LL W=430.00n L=60.00n
MM35 net0144 A VSS VPW N12LL W=430.00n L=60.00n
MM8 net108 CI net0227 VNW P12LL W=375.00n L=60.00n
MM7 net0231 B VDD VNW P12LL W=375.00n L=60.00n
MM6 net0227 A net0231 VNW P12LL W=375.00n L=60.00n
MM10 net0212 B VDD VNW P12LL W=640.00n L=60.00n
MM11 net0212 CI VDD VNW P12LL W=640.00n L=60.00n
MM2 net100 A net0183 VNW P12LL W=440.00n L=60.00n
MM3 net0183 B VDD VNW P12LL W=400.00n L=60.00n
MM32 CO net100 VDD VNW P12LL W=1.08u L=60.00n
MM12 net108 net100 net0212 VNW P12LL W=375.00n L=60.00n
MM9 net0212 A VDD VNW P12LL W=640.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=1.08u L=60.00n
MM18 net0203 A VDD VNW P12LL W=650.00n L=60.00n
MM1 net0203 B VDD VNW P12LL W=650.00n L=60.00n
MM0 net100 CI net0203 VNW P12LL W=440.00n L=60.00n
.ENDS AD1HSV4C
****Sub-Circuit for AD1HSV4R, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1HSV4R A B CI CO S VDD VSS
MM41 net0196 cin net78 VPW N12LL W=430.00n L=60.00n
MM42 norab CI net78 VPW N12LL W=430.00n L=60.00n
MMN1 xo norab VSS VPW N12LL W=880.00n L=60.00n
MM3 norab A VSS VPW N12LL W=700.00n L=60.00n
MM0 xo A net0164 VPW N12LL W=1.08u L=60.00n
MM2 norab B VSS VPW N12LL W=700.00n L=60.00n
MM7 net0164 B VSS VPW N12LL W=1.08u L=60.00n
MM8 xn xo VSS VPW N12LL W=430.00n L=60.00n
MM10 net0124 B VSS VPW N12LL W=520.00n L=60.00n
MM11 net0196 A net0124 VPW N12LL W=520.00n L=60.00n
MM27 cin CI VSS VPW N12LL W=220.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=860.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=860.00n L=60.00n
MM36 xn cin net108 VPW N12LL W=430.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=430.00n L=60.00n
MM43 net0196 CI net78 VNW P12LL W=540.00n L=60.00n
MM44 norab cin net78 VNW P12LL W=540.00n L=60.00n
MM12 net0196 A VDD VNW P12LL W=440.00n L=60.00n
MM13 net0196 B VDD VNW P12LL W=440.00n L=60.00n
MM28 cin CI VDD VNW P12LL W=270.00n L=60.00n
MM21 CO net78 VDD VNW P12LL W=1.08u L=60.00n
MM20 S net108 VDD VNW P12LL W=1.08u L=60.00n
MM4 norab A net0215 VNW P12LL W=1.3u L=60.00n
MMP1 net0223 A VDD VNW P12LL W=1.3u L=60.00n
MM1 xo norab net0223 VNW P12LL W=1.08u L=60.00n
MM6 net0223 B VDD VNW P12LL W=1.3u L=60.00n
MM5 net0215 B VDD VNW P12LL W=1.3u L=60.00n
MM9 xn xo VDD VNW P12LL W=540.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=540.00n L=60.00n
MM40 xo cin net108 VNW P12LL W=540.00n L=60.00n
.ENDS AD1HSV4R
****Sub-Circuit for AD1HSV4T, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT AD1HSV4T A B CI CO S VDD VSS
MM10 net117 B VSS VPW N12LL W=860.00n L=60.00n
MM41 cin xo net78 VPW N12LL W=430.00n L=60.00n
MM42 net117 xn net78 VPW N12LL W=430.00n L=60.00n
MMN1 xo net0164 VSS VPW N12LL W=700.00n L=60.00n
MM2 net0164 B VSS VPW N12LL W=700.00n L=60.00n
MM3 net0164 A VSS VPW N12LL W=700.00n L=60.00n
MM0 xo A net0176 VPW N12LL W=860.00n L=60.00n
MM7 net0176 B VSS VPW N12LL W=860.00n L=60.00n
MM31 cin CI VSS VPW N12LL W=860.00n L=60.00n
MM22 CO net78 VSS VPW N12LL W=860.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=860.00n L=60.00n
MM36 xn cin net108 VPW N12LL W=420.00n L=60.00n
MM38 xo CI net108 VPW N12LL W=420.00n L=60.00n
MM8 xn xo VSS VPW N12LL W=420.00n L=60.00n
MM11 net117 B VDD VNW P12LL W=1.08u L=60.00n
MM43 cin xn net78 VNW P12LL W=540.00n L=60.00n
MM44 net117 xo net78 VNW P12LL W=540.00n L=60.00n
MM4 net0164 A net0235 VNW P12LL W=1.3u L=60.00n
MMP1 net0227 A VDD VNW P12LL W=1.3u L=60.00n
MM1 xo net0164 net0227 VNW P12LL W=1.08u L=60.00n
MM6 net0227 B VDD VNW P12LL W=1.3u L=60.00n
MM5 net0235 B VDD VNW P12LL W=1.3u L=60.00n
MM32 cin CI VDD VNW P12LL W=1.08u L=60.00n
MM21 CO net78 VDD VNW P12LL W=1.08u L=60.00n
MM20 S net108 VDD VNW P12LL W=1.08u L=60.00n
MM9 xn xo VDD VNW P12LL W=530.00n L=60.00n
MM39 xn CI net108 VNW P12LL W=530.00n L=60.00n
MM40 xo cin net108 VNW P12LL W=530.00n L=60.00n
.ENDS AD1HSV4T
****Sub-Circuit for AD2CSCINHSV1, Wed May 25 11:46:50 CST 2011****
.SUBCKT AD2CSCINHSV1 A B CI0N CI1N CO0 CO1 CS S VDD VSS
MM79 ci0 CI0N VSS VPW N12LL W=180.00n L=60.00n
MM78 ci1 CI1N VSS VPW N12LL W=180.00n L=60.00n
MM68 net0415 norab VSS VPW N12LL W=350.00n L=60.00n
MM70 net0227 net0415 VSS VPW N12LL W=330.00n L=60.00n
MM71 net0327 nandab net0227 VPW N12LL W=330.00n L=60.00n
MM61 net0231 ci1 net0395 VPW N12LL W=180.00n L=60.00n
MM60 net0235 CI1N net0395 VPW N12LL W=180.00n L=60.00n
MM55 net0235 CI0N net0219 VPW N12LL W=180.00n L=60.00n
MM54 net0231 ci0 net0219 VPW N12LL W=180.00n L=60.00n
MM52 csn CS VSS VPW N12LL W=180.00n L=60.00n
MM51 ci1nn CI1N VSS VPW N12LL W=180.00n L=60.00n
MM48 ci0nn CI0N VSS VPW N12LL W=180.00n L=60.00n
MM3 norab A VSS VPW N12LL W=280.00n L=60.00n
MM18 net0132 B VSS VPW N12LL W=430.00n L=60.00n
MM23 nandab A net0132 VPW N12LL W=430.00n L=60.00n
MM2 norab B VSS VPW N12LL W=280.00n L=60.00n
MM26 nandab CI0N net0143 VPW N12LL W=180.00n L=60.00n
MM29 norab ci0nn net0143 VPW N12LL W=180.00n L=60.00n
MM8 net0235 net0231 VSS VPW N12LL W=180.00n L=60.00n
MM30 CO0 net0143 VSS VPW N12LL W=350.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=350.00n L=60.00n
MM62 net0231 net0327 VSS VPW N12LL W=350.00n L=60.00n
MM34 nandab CI1N net0155 VPW N12LL W=180.00n L=60.00n
MM35 norab ci1nn net0155 VPW N12LL W=180.00n L=60.00n
MM37 CO1 net0155 VSS VPW N12LL W=350.00n L=60.00n
MM36 net0219 csn net108 VPW N12LL W=180.00n L=60.00n
MM38 net0395 CS net108 VPW N12LL W=180.00n L=60.00n
MM80 ci0 CI0N VDD VNW P12LL W=220.00n L=60.00n
MM77 ci1 CI1N VDD VNW P12LL W=220.00n L=60.00n
MM69 net0415 norab VDD VNW P12LL W=440.00n L=60.00n
MM72 net0327 nandab VDD VNW P12LL W=280.00n L=60.00n
MM73 net0327 net0415 VDD VNW P12LL W=280.00n L=60.00n
MM59 net0231 CI1N net0395 VNW P12LL W=220.00n L=60.00n
MM58 net0235 ci1 net0395 VNW P12LL W=220.00n L=60.00n
MM57 net0235 ci0 net0219 VNW P12LL W=220.00n L=60.00n
MM56 net0231 CI0N net0219 VNW P12LL W=220.00n L=60.00n
MM53 csn CS VDD VNW P12LL W=220.00n L=60.00n
MM50 ci1nn CI1N VDD VNW P12LL W=220.00n L=60.00n
MM49 ci0nn CI0N VDD VNW P12LL W=220.00n L=60.00n
MM63 net0231 net0327 VDD VNW P12LL W=440.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=390.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=390.00n L=60.00n
MM31 nandab ci0nn net0143 VNW P12LL W=220.00n L=60.00n
MM32 norab CI0N net0143 VNW P12LL W=220.00n L=60.00n
MM33 CO0 net0143 VDD VNW P12LL W=440.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=440.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=520.00n L=60.00n
MM45 nandab ci1nn net0155 VNW P12LL W=220.00n L=60.00n
MM46 norab CI1N net0155 VNW P12LL W=220.00n L=60.00n
MM47 CO1 net0155 VDD VNW P12LL W=440.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=520.00n L=60.00n
MM9 net0235 net0231 VDD VNW P12LL W=220.00n L=60.00n
MM39 net0219 CS net108 VNW P12LL W=220.00n L=60.00n
MM40 net0395 csn net108 VNW P12LL W=220.00n L=60.00n
.ENDS AD2CSCINHSV1
****Sub-Circuit for AD2CSCINHSV2, Wed May 25 13:06:45 CST 2011****
.SUBCKT AD2CSCINHSV2 A B CI0N CI1N CO0 CO1 CS S VDD VSS
MM74 ci1 CI1N VSS VPW N12LL W=220.00n L=60.00n
MM75 ci0 CI0N VSS VPW N12LL W=220.00n L=60.00n
MM68 net0415 norab VSS VPW N12LL W=370.00n L=60.00n
MM70 net0227 net0415 VSS VPW N12LL W=330.00n L=60.00n
MM71 net0327 nandab net0227 VPW N12LL W=330.00n L=60.00n
MM61 net0231 ci1 net0395 VPW N12LL W=220.00n L=60.00n
MM60 net0235 CI1N net0395 VPW N12LL W=220.00n L=60.00n
MM55 net0235 CI0N net0219 VPW N12LL W=220.00n L=60.00n
MM54 net0231 ci0 net0219 VPW N12LL W=220.00n L=60.00n
MM52 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM51 ci1nn CI1N VSS VPW N12LL W=220.00n L=60.00n
MM48 ci0nn CI0N VSS VPW N12LL W=220.00n L=60.00n
MM3 norab A VSS VPW N12LL W=350.00n L=60.00n
MM18 net0132 B VSS VPW N12LL W=430.00n L=60.00n
MM23 nandab A net0132 VPW N12LL W=430.00n L=60.00n
MM2 norab B VSS VPW N12LL W=350.00n L=60.00n
MM26 nandab CI0N net0143 VPW N12LL W=220.00n L=60.00n
MM29 norab ci0nn net0143 VPW N12LL W=220.00n L=60.00n
MM8 net0235 net0231 VSS VPW N12LL W=220.00n L=60.00n
MM30 CO0 net0143 VSS VPW N12LL W=430.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=430.00n L=60.00n
MM62 net0231 net0327 VSS VPW N12LL W=350.00n L=60.00n
MM34 nandab CI1N net0155 VPW N12LL W=220.00n L=60.00n
MM35 norab ci1nn net0155 VPW N12LL W=220.00n L=60.00n
MM37 CO1 net0155 VSS VPW N12LL W=370.00n L=60.00n
MM36 net0219 csn net108 VPW N12LL W=220.00n L=60.00n
MM38 net0395 CS net108 VPW N12LL W=220.00n L=60.00n
MM76 ci1 CI1N VDD VNW P12LL W=270.00n L=60.00n
MM77 ci0 CI0N VDD VNW P12LL W=270.00n L=60.00n
MM69 net0415 norab VDD VNW P12LL W=515.00n L=60.00n
MM72 net0327 nandab VDD VNW P12LL W=280.00n L=60.00n
MM73 net0327 net0415 VDD VNW P12LL W=280.00n L=60.00n
MM59 net0231 CI1N net0395 VNW P12LL W=270.00n L=60.00n
MM58 net0235 ci1 net0395 VNW P12LL W=270.00n L=60.00n
MM57 net0235 ci0 net0219 VNW P12LL W=270.00n L=60.00n
MM56 net0231 CI0N net0219 VNW P12LL W=270.00n L=60.00n
MM53 csn CS VDD VNW P12LL W=270.00n L=60.00n
MM50 ci1nn CI1N VDD VNW P12LL W=270.00n L=60.00n
MM49 ci0nn CI0N VDD VNW P12LL W=270.00n L=60.00n
MM63 net0231 net0327 VDD VNW P12LL W=515.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=420.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=420.00n L=60.00n
MM31 nandab ci0nn net0143 VNW P12LL W=270.00n L=60.00n
MM32 norab CI0N net0143 VNW P12LL W=270.00n L=60.00n
MM33 CO0 net0143 VDD VNW P12LL W=540.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=540.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=650.00n L=60.00n
MM45 nandab ci1nn net0155 VNW P12LL W=270.00n L=60.00n
MM46 norab CI1N net0155 VNW P12LL W=270.00n L=60.00n
MM47 CO1 net0155 VDD VNW P12LL W=515.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=650.00n L=60.00n
MM9 net0235 net0231 VDD VNW P12LL W=270.00n L=60.00n
MM39 net0219 CS net108 VNW P12LL W=270.00n L=60.00n
MM40 net0395 csn net108 VNW P12LL W=270.00n L=60.00n
.ENDS AD2CSCINHSV2
****Sub-Circuit for AD2CSCINHSV4, Thu May 26 09:11:25 CST 2011****
.SUBCKT AD2CSCINHSV4 A B CI0N CI1N CO0 CO1 CS S VDD VSS
MM74 ci1 CI1N VSS VPW N12LL W=220.00n L=60.00n
MM75 ci0 CI0N VSS VPW N12LL W=220.00n L=60.00n
MM68 net0415 norab VSS VPW N12LL W=750.00n L=60.00n
MM70 net0227 net0415 VSS VPW N12LL W=750.00n L=60.00n
MM71 net0327 nandab net0227 VPW N12LL W=750.00n L=60.00n
MM61 net0231 ci1 net0395 VPW N12LL W=430.00n L=60.00n
MM60 net0235 CI1N net0395 VPW N12LL W=430.00n L=60.00n
MM55 net0235 CI0N net0219 VPW N12LL W=430.00n L=60.00n
MM54 net0231 ci0 net0219 VPW N12LL W=430.00n L=60.00n
MM52 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM51 ci1nn CI1N VSS VPW N12LL W=220.00n L=60.00n
MM48 ci0nn CI0N VSS VPW N12LL W=220.00n L=60.00n
MM3 norab A VSS VPW N12LL W=700.00n L=60.00n
MM18 net0132 B VSS VPW N12LL W=860.00n L=60.00n
MM23 nandab A net0132 VPW N12LL W=860.00n L=60.00n
MM2 norab B VSS VPW N12LL W=700.00n L=60.00n
MM26 nandab CI0N net0143 VPW N12LL W=430.00n L=60.00n
MM29 norab ci0nn net0143 VPW N12LL W=430.00n L=60.00n
MM8 net0235 net0231 VSS VPW N12LL W=375.00n L=60.00n
MM30 CO0 net0143 VSS VPW N12LL W=860.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=860.00n L=60.00n
MM62 net0231 net0327 VSS VPW N12LL W=750.00n L=60.00n
MM34 nandab CI1N net0155 VPW N12LL W=430.00n L=60.00n
MM35 norab ci1nn net0155 VPW N12LL W=430.00n L=60.00n
MM37 CO1 net0155 VSS VPW N12LL W=740.00n L=60.00n
MM36 net0219 csn net108 VPW N12LL W=430.00n L=60.00n
MM38 net0395 CS net108 VPW N12LL W=430.00n L=60.00n
MM76 ci1 CI1N VDD VNW P12LL W=270.00n L=60.00n
MM77 ci0 CI0N VDD VNW P12LL W=270.00n L=60.00n
MM69 net0415 norab VDD VNW P12LL W=1.03u L=60.00n
MM72 net0327 nandab VDD VNW P12LL W=560.00n L=60.00n
MM73 net0327 net0415 VDD VNW P12LL W=560.00n L=60.00n
MM59 net0231 CI1N net0395 VNW P12LL W=540.00n L=60.00n
MM58 net0235 ci1 net0395 VNW P12LL W=540.00n L=60.00n
MM57 net0235 ci0 net0219 VNW P12LL W=540.00n L=60.00n
MM56 net0231 CI0N net0219 VNW P12LL W=540.00n L=60.00n
MM53 csn CS VDD VNW P12LL W=270.00n L=60.00n
MM50 ci1nn CI1N VDD VNW P12LL W=270.00n L=60.00n
MM49 ci0nn CI0N VDD VNW P12LL W=270.00n L=60.00n
MM63 net0231 net0327 VDD VNW P12LL W=1.03u L=60.00n
MM24 nandab A VDD VNW P12LL W=960.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=960.00n L=60.00n
MM31 nandab ci0nn net0143 VNW P12LL W=515.00n L=60.00n
MM32 norab CI0N net0143 VNW P12LL W=515.00n L=60.00n
MM33 CO0 net0143 VDD VNW P12LL W=1.08u L=60.00n
MM20 S net108 VDD VNW P12LL W=1.08u L=60.00n
MM4 norab A net0215 VNW P12LL W=1.3u L=60.00n
MM45 nandab ci1nn net0155 VNW P12LL W=540.00n L=60.00n
MM46 norab CI1N net0155 VNW P12LL W=540.00n L=60.00n
MM47 CO1 net0155 VDD VNW P12LL W=1.03u L=60.00n
MM5 net0215 B VDD VNW P12LL W=1.3u L=60.00n
MM9 net0235 net0231 VDD VNW P12LL W=515.00n L=60.00n
MM39 net0219 CS net108 VNW P12LL W=540.00n L=60.00n
MM40 net0395 csn net108 VNW P12LL W=540.00n L=60.00n
.ENDS AD2CSCINHSV4
****Sub-Circuit for AD2CSCONHSV1, Thu May 26 14:23:16 CST 2011****
.SUBCKT AD2CSCONHSV1 A B CI0 CI1 CO0N CO1N CS S VDD VSS
MM78 ci1nnn CI1 VSS VPW N12LL W=180.00n L=60.00n
MM79 ci0nnn CI0 VSS VPW N12LL W=180.00n L=60.00n
MM75 andab nandab VSS VPW N12LL W=180.00n L=60.00n
MM70 net0227 orab VSS VPW N12LL W=330.00n L=60.00n
MM71 net0327 nandab net0227 VPW N12LL W=330.00n L=60.00n
MM61 net0231 ci1nnn net0395 VPW N12LL W=180.00n L=60.00n
MM60 net0235 CI1 net0395 VPW N12LL W=180.00n L=60.00n
MM55 net0235 CI0 net0219 VPW N12LL W=180.00n L=60.00n
MM54 net0231 ci0nnn net0219 VPW N12LL W=180.00n L=60.00n
MM52 csn CS VSS VPW N12LL W=180.00n L=60.00n
MM51 ci1n CI1 VSS VPW N12LL W=180.00n L=60.00n
MM48 ci0n CI0 VSS VPW N12LL W=180.00n L=60.00n
MM3 norab A VSS VPW N12LL W=280.00n L=60.00n
MM74 orab norab VSS VPW N12LL W=350.00n L=60.00n
MM18 net0132 B VSS VPW N12LL W=430.00n L=60.00n
MM23 nandab A net0132 VPW N12LL W=430.00n L=60.00n
MM2 norab B VSS VPW N12LL W=280.00n L=60.00n
MM26 andab ci0n net0143 VPW N12LL W=180.00n L=60.00n
MM29 orab CI0 net0143 VPW N12LL W=180.00n L=60.00n
MM8 net0231 net0235 VSS VPW N12LL W=180.00n L=60.00n
MM30 CO0N net0143 VSS VPW N12LL W=350.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=350.00n L=60.00n
MM62 net0235 net0327 VSS VPW N12LL W=345.00n L=60.00n
MM34 andab ci1n net0155 VPW N12LL W=180.00n L=60.00n
MM35 orab CI1 net0155 VPW N12LL W=180.00n L=60.00n
MM37 CO1N net0155 VSS VPW N12LL W=350.00n L=60.00n
MM36 net0219 csn net108 VPW N12LL W=180.00n L=60.00n
MM38 net0395 CS net108 VPW N12LL W=180.00n L=60.00n
MM80 ci1nnn CI1 VDD VNW P12LL W=220.00n L=60.00n
MM81 ci0nnn CI0 VDD VNW P12LL W=220.00n L=60.00n
MM77 andab nandab VDD VNW P12LL W=220.00n L=60.00n
MM72 net0327 nandab VDD VNW P12LL W=280.00n L=60.00n
MM73 net0327 orab VDD VNW P12LL W=280.00n L=60.00n
MM59 net0231 CI1 net0395 VNW P12LL W=220.00n L=60.00n
MM58 net0235 ci1nnn net0395 VNW P12LL W=220.00n L=60.00n
MM57 net0235 ci0nnn net0219 VNW P12LL W=220.00n L=60.00n
MM56 net0231 CI0 net0219 VNW P12LL W=220.00n L=60.00n
MM53 csn CS VDD VNW P12LL W=220.00n L=60.00n
MM50 ci1n CI1 VDD VNW P12LL W=220.00n L=60.00n
MM49 ci0n CI0 VDD VNW P12LL W=220.00n L=60.00n
MM76 orab norab VDD VNW P12LL W=440.00n L=60.00n
MM63 net0235 net0327 VDD VNW P12LL W=440.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=390.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=390.00n L=60.00n
MM31 andab CI0 net0143 VNW P12LL W=220.00n L=60.00n
MM32 orab ci0n net0143 VNW P12LL W=220.00n L=60.00n
MM33 CO0N net0143 VDD VNW P12LL W=440.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=440.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=520.00n L=60.00n
MM45 andab CI1 net0155 VNW P12LL W=220.00n L=60.00n
MM46 orab ci1n net0155 VNW P12LL W=220.00n L=60.00n
MM47 CO1N net0155 VDD VNW P12LL W=440.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=520.00n L=60.00n
MM9 net0231 net0235 VDD VNW P12LL W=220.00n L=60.00n
MM39 net0219 CS net108 VNW P12LL W=220.00n L=60.00n
MM40 net0395 csn net108 VNW P12LL W=220.00n L=60.00n
.ENDS AD2CSCONHSV1
****Sub-Circuit for AD2CSCONHSV2, Thu May 26 15:40:13 CST 2011****
.SUBCKT AD2CSCONHSV2 A B CI0 CI1 CO0N CO1N CS S VDD VSS
MM78 ci1nnn CI1 VSS VPW N12LL W=220.00n L=60.00n
MM79 ci0nnn CI0 VSS VPW N12LL W=220.00n L=60.00n
MM75 andab nandab VSS VPW N12LL W=220.00n L=60.00n
MM70 net0227 orab VSS VPW N12LL W=330.00n L=60.00n
MM71 net0327 nandab net0227 VPW N12LL W=330.00n L=60.00n
MM61 net0231 ci1nnn net0395 VPW N12LL W=220.00n L=60.00n
MM60 net0235 CI1 net0395 VPW N12LL W=220.00n L=60.00n
MM55 net0235 CI0 net0219 VPW N12LL W=220.00n L=60.00n
MM54 net0231 ci0nnn net0219 VPW N12LL W=220.00n L=60.00n
MM52 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM51 ci1n CI1 VSS VPW N12LL W=220.00n L=60.00n
MM48 ci0n CI0 VSS VPW N12LL W=220.00n L=60.00n
MM3 norab A VSS VPW N12LL W=350.00n L=60.00n
MM74 orab norab VSS VPW N12LL W=430.00n L=60.00n
MM18 net0132 B VSS VPW N12LL W=430.00n L=60.00n
MM23 nandab A net0132 VPW N12LL W=430.00n L=60.00n
MM2 norab B VSS VPW N12LL W=350.00n L=60.00n
MM26 andab ci0n net0143 VPW N12LL W=220.00n L=60.00n
MM29 orab CI0 net0143 VPW N12LL W=220.00n L=60.00n
MM8 net0231 net0235 VSS VPW N12LL W=220.00n L=60.00n
MM30 CO0N net0143 VSS VPW N12LL W=430.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=430.00n L=60.00n
MM62 net0235 net0327 VSS VPW N12LL W=345.00n L=60.00n
MM34 andab ci1n net0155 VPW N12LL W=220.00n L=60.00n
MM35 orab CI1 net0155 VPW N12LL W=220.00n L=60.00n
MM37 CO1N net0155 VSS VPW N12LL W=375.00n L=60.00n
MM36 net0219 csn net108 VPW N12LL W=220.00n L=60.00n
MM38 net0395 CS net108 VPW N12LL W=220.00n L=60.00n
MM80 ci1nnn CI1 VDD VNW P12LL W=270.00n L=60.00n
MM81 ci0nnn CI0 VDD VNW P12LL W=270.00n L=60.00n
MM77 andab nandab VDD VNW P12LL W=270.00n L=60.00n
MM72 net0327 nandab VDD VNW P12LL W=280.00n L=60.00n
MM73 net0327 orab VDD VNW P12LL W=280.00n L=60.00n
MM59 net0231 CI1 net0395 VNW P12LL W=270.00n L=60.00n
MM58 net0235 ci1nnn net0395 VNW P12LL W=270.00n L=60.00n
MM57 net0235 ci0nnn net0219 VNW P12LL W=270.00n L=60.00n
MM56 net0231 CI0 net0219 VNW P12LL W=270.00n L=60.00n
MM53 csn CS VDD VNW P12LL W=270.00n L=60.00n
MM50 ci1n CI1 VDD VNW P12LL W=270.00n L=60.00n
MM49 ci0n CI0 VDD VNW P12LL W=270.00n L=60.00n
MM76 orab norab VDD VNW P12LL W=540.00n L=60.00n
MM63 net0235 net0327 VDD VNW P12LL W=515.00n L=60.00n
MM24 nandab A VDD VNW P12LL W=420.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=420.00n L=60.00n
MM31 andab CI0 net0143 VNW P12LL W=270.00n L=60.00n
MM32 orab ci0n net0143 VNW P12LL W=270.00n L=60.00n
MM33 CO0N net0143 VDD VNW P12LL W=540.00n L=60.00n
MM20 S net108 VDD VNW P12LL W=540.00n L=60.00n
MM4 norab A net0215 VNW P12LL W=650.00n L=60.00n
MM45 andab CI1 net0155 VNW P12LL W=270.00n L=60.00n
MM46 orab ci1n net0155 VNW P12LL W=270.00n L=60.00n
MM47 CO1N net0155 VDD VNW P12LL W=515.00n L=60.00n
MM5 net0215 B VDD VNW P12LL W=650.00n L=60.00n
MM9 net0231 net0235 VDD VNW P12LL W=270.00n L=60.00n
MM39 net0219 CS net108 VNW P12LL W=270.00n L=60.00n
MM40 net0395 csn net108 VNW P12LL W=270.00n L=60.00n
.ENDS AD2CSCONHSV2
****Sub-Circuit for AD2CSCONHSV4, Fri May 27 09:16:23 CST 2011****
.SUBCKT AD2CSCONHSV4 A B CI0 CI1 CO0N CO1N CS S VDD VSS
MM78 ci1nnn CI1 VSS VPW N12LL W=220.00n L=60.00n
MM79 ci0nnn CI0 VSS VPW N12LL W=215.00n L=60.00n
MM75 andab nandab VSS VPW N12LL W=430.00n L=60.00n
MM70 net0227 orab VSS VPW N12LL W=750.00n L=60.00n
MM71 net0327 nandab net0227 VPW N12LL W=750.00n L=60.00n
MM61 net0231 ci1nnn net0395 VPW N12LL W=430.00n L=60.00n
MM60 net0235 CI1 net0395 VPW N12LL W=430.00n L=60.00n
MM55 net0235 CI0 net0219 VPW N12LL W=430.00n L=60.00n
MM54 net0231 ci0nnn net0219 VPW N12LL W=430.00n L=60.00n
MM52 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM51 ci1n CI1 VSS VPW N12LL W=220.00n L=60.00n
MM48 ci0n CI0 VSS VPW N12LL W=220.00n L=60.00n
MM3 norab A VSS VPW N12LL W=700.00n L=60.00n
MM74 orab norab VSS VPW N12LL W=860.00n L=60.00n
MM18 net0132 B VSS VPW N12LL W=860.00n L=60.00n
MM23 nandab A net0132 VPW N12LL W=860.00n L=60.00n
MM2 norab B VSS VPW N12LL W=700.00n L=60.00n
MM26 andab ci0n net0143 VPW N12LL W=430.00n L=60.00n
MM29 orab CI0 net0143 VPW N12LL W=430.00n L=60.00n
MM8 net0231 net0235 VSS VPW N12LL W=375.00n L=60.00n
MM30 CO0N net0143 VSS VPW N12LL W=860.00n L=60.00n
MM19 S net108 VSS VPW N12LL W=860.00n L=60.00n
MM62 net0235 net0327 VSS VPW N12LL W=750.00n L=60.00n
MM34 andab ci1n net0155 VPW N12LL W=430.00n L=60.00n
MM35 orab CI1 net0155 VPW N12LL W=430.00n L=60.00n
MM37 CO1N net0155 VSS VPW N12LL W=740.00n L=60.00n
MM36 net0219 csn net108 VPW N12LL W=430.00n L=60.00n
MM38 net0395 CS net108 VPW N12LL W=430.00n L=60.00n
MM80 ci1nnn CI1 VDD VNW P12LL W=270.00n L=60.00n
MM81 ci0nnn CI0 VDD VNW P12LL W=270.00n L=60.00n
MM77 andab nandab VDD VNW P12LL W=540.00n L=60.00n
MM72 net0327 nandab VDD VNW P12LL W=560.00n L=60.00n
MM73 net0327 orab VDD VNW P12LL W=560.00n L=60.00n
MM59 net0231 CI1 net0395 VNW P12LL W=540.00n L=60.00n
MM58 net0235 ci1nnn net0395 VNW P12LL W=540.00n L=60.00n
MM57 net0235 ci0nnn net0219 VNW P12LL W=540.00n L=60.00n
MM56 net0231 CI0 net0219 VNW P12LL W=540.00n L=60.00n
MM53 csn CS VDD VNW P12LL W=270.00n L=60.00n
MM50 ci1n CI1 VDD VNW P12LL W=270.00n L=60.00n
MM49 ci0n CI0 VDD VNW P12LL W=270.00n L=60.00n
MM76 orab norab VDD VNW P12LL W=1.08u L=60.00n
MM63 net0235 net0327 VDD VNW P12LL W=1.03u L=60.00n
MM24 nandab A VDD VNW P12LL W=960.00n L=60.00n
MM25 nandab B VDD VNW P12LL W=960.00n L=60.00n
MM31 andab CI0 net0143 VNW P12LL W=500.00n L=60.00n
MM32 orab ci0n net0143 VNW P12LL W=500.00n L=60.00n
MM33 CO0N net0143 VDD VNW P12LL W=1.08u L=60.00n
MM20 S net108 VDD VNW P12LL W=1.08u L=60.00n
MM4 norab A net0215 VNW P12LL W=1.3u L=60.00n
MM45 andab CI1 net0155 VNW P12LL W=540.00n L=60.00n
MM46 orab ci1n net0155 VNW P12LL W=540.00n L=60.00n
MM47 CO1N net0155 VDD VNW P12LL W=1.03u L=60.00n
MM5 net0215 B VDD VNW P12LL W=1.3u L=60.00n
MM9 net0231 net0235 VDD VNW P12LL W=515.00n L=60.00n
MM39 net0219 CS net108 VNW P12LL W=540.00n L=60.00n
MM40 net0395 csn net108 VNW P12LL W=540.00n L=60.00n
.ENDS AD2CSCONHSV4
****Sub-Circuit for ADH1CINHSV1, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1CINHSV1 A CIN CO S VDD VSS
MM45 net_072 net35 VDD VNW P12LL W=180.00n L=60.00n
MM46 net_072 A VDD VNW P12LL W=180.00n L=60.00n
MM48 net45 net35 S VNW P12LL W=440.00n L=60.00n
MM32 net35 CIN VDD VNW P12LL W=270.00n L=60.00n
MM29 net45 net46 VDD VNW P12LL W=440.00n L=60.00n
MM28 net46 A VDD VNW P12LL W=440.00n L=60.00n
MM39 net46 CIN S VNW P12LL W=440.00n L=60.00n
MM0 CO net_072 VDD VNW P12LL W=440.00n L=60.00n
MM27 net46 A VSS VPW N12LL W=350.00n L=60.00n
MM47 net45 CIN S VPW N12LL W=350.00n L=60.00n
MM30 net45 net46 VSS VPW N12LL W=350.00n L=60.00n
MM1 CO net_072 VSS VPW N12LL W=350.00n L=60.00n
MM43 net_072 A net_95 VPW N12LL W=210.00n L=60.00n
MM31 net35 CIN VSS VPW N12LL W=220.00n L=60.00n
MM44 net_95 net35 VSS VPW N12LL W=210.00n L=60.00n
MM36 net46 net35 S VPW N12LL W=350.00n L=60.00n
.ENDS ADH1CINHSV1
****Sub-Circuit for ADH1CINHSV1C, Thu May 19 13:57:40 CST 2011****
.SUBCKT ADH1CINHSV1C A CIN CO S VDD VSS
MM7 net85 A net88 VNW P12LL W=200.00n L=60.00n
MM32 net35 CIN VDD VNW P12LL W=270.00n L=60.00n
MM0 CO acinn VDD VNW P12LL W=440.00n L=60.00n
MM6 net88 net35 VDD VNW P12LL W=200.00n L=60.00n
MM10 S net85 VDD VNW P12LL W=440.00n L=60.00n
MM45 acinn net35 VDD VNW P12LL W=180.00n L=60.00n
MM46 acinn A VDD VNW P12LL W=180.00n L=60.00n
MM4 net85 acinn VDD VNW P12LL W=200.00n L=60.00n
MM8 net117 A VSS VPW N12LL W=180.00n L=60.00n
MM9 net117 net35 VSS VPW N12LL W=180.00n L=60.00n
MM1 CO acinn VSS VPW N12LL W=350.00n L=60.00n
MM43 acinn A net_079 VPW N12LL W=210.00n L=60.00n
MM31 net35 CIN VSS VPW N12LL W=220.00n L=60.00n
MM44 net_079 net35 VSS VPW N12LL W=210.00n L=60.00n
MM11 S net85 VSS VPW N12LL W=350.00n L=60.00n
MM5 net85 acinn net117 VPW N12LL W=180.00n L=60.00n
.ENDS ADH1CINHSV1C
****Sub-Circuit for ADH1CINHSV2, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1CINHSV2 A CIN CO S VDD VSS
MM45 net_072 net35 VDD VNW P12LL W=220.00n L=60.00n
MM46 net_072 A VDD VNW P12LL W=220.00n L=60.00n
MM48 net45 net35 S VNW P12LL W=540.00n L=60.00n
MM32 net35 CIN VDD VNW P12LL W=270.00n L=60.00n
MM29 net45 net46 VDD VNW P12LL W=540.00n L=60.00n
MM28 net46 A VDD VNW P12LL W=540.00n L=60.00n
MM39 net46 CIN S VNW P12LL W=540.00n L=60.00n
MM0 CO net_072 VDD VNW P12LL W=540.00n L=60.00n
MM27 net46 A VSS VPW N12LL W=430.00n L=60.00n
MM47 net45 CIN S VPW N12LL W=430.00n L=60.00n
MM30 net45 net46 VSS VPW N12LL W=430.00n L=60.00n
MM1 CO net_072 VSS VPW N12LL W=430.00n L=60.00n
MM43 net_072 A net_95 VPW N12LL W=260.00n L=60.00n
MM31 net35 CIN VSS VPW N12LL W=220.00n L=60.00n
MM44 net_95 net35 VSS VPW N12LL W=260.00n L=60.00n
MM36 net46 net35 S VPW N12LL W=430.00n L=60.00n
.ENDS ADH1CINHSV2
****Sub-Circuit for ADH1CINHSV2C, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1CINHSV2C A CIN CO S VDD VSS
MM7 net85 A net88 VNW P12LL W=220.00n L=60.00n
MM32 net35 CIN VDD VNW P12LL W=270.00n L=60.00n
MM0 CO acinn VDD VNW P12LL W=540.00n L=60.00n
MM6 net88 net35 VDD VNW P12LL W=220.00n L=60.00n
MM10 S net85 VDD VNW P12LL W=540.00n L=60.00n
MM45 acinn net35 VDD VNW P12LL W=220.00n L=60.00n
MM46 acinn A VDD VNW P12LL W=220.00n L=60.00n
MM4 net85 acinn VDD VNW P12LL W=220.00n L=60.00n
MM8 net117 A VSS VPW N12LL W=320.00n L=60.00n
MM9 net117 net35 VSS VPW N12LL W=320.00n L=60.00n
MM1 CO acinn VSS VPW N12LL W=430.00n L=60.00n
MM43 acinn A net_079 VPW N12LL W=260.00n L=60.00n
MM31 net35 CIN VSS VPW N12LL W=220.00n L=60.00n
MM44 net_079 net35 VSS VPW N12LL W=260.00n L=60.00n
MM11 S net85 VSS VPW N12LL W=430.00n L=60.00n
MM5 net85 acinn net117 VPW N12LL W=180.00n L=60.00n
.ENDS ADH1CINHSV2C
****Sub-Circuit for ADH1CINHSV4, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1CINHSV4 A CIN CO S VDD VSS
MM45 net_072 net35 VDD VNW P12LL W=440.00n L=60.00n
MM46 net_072 A VDD VNW P12LL W=440.00n L=60.00n
MM48 net45 net35 S VNW P12LL W=1.08u L=60.00n
MM32 net35 CIN VDD VNW P12LL W=430.00n L=60.00n
MM29 net45 net46 VDD VNW P12LL W=1.08u L=60.00n
MM28 net46 A VDD VNW P12LL W=1.08u L=60.00n
MM39 net46 CIN S VNW P12LL W=1.08u L=60.00n
MM0 CO net_072 VDD VNW P12LL W=1.08u L=60.00n
MM27 net46 A VSS VPW N12LL W=860.00n L=60.00n
MM47 net45 CIN S VPW N12LL W=860.00n L=60.00n
MM30 net45 net46 VSS VPW N12LL W=860.00n L=60.00n
MM1 CO net_072 VSS VPW N12LL W=860.00n L=60.00n
MM43 net_072 A net_95 VPW N12LL W=490.00n L=60.00n
MM31 net35 CIN VSS VPW N12LL W=350.00n L=60.00n
MM44 net_95 net35 VSS VPW N12LL W=490.00n L=60.00n
MM36 net46 net35 S VPW N12LL W=860.00n L=60.00n
.ENDS ADH1CINHSV4
****Sub-Circuit for ADH1CINHSV4C, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1CINHSV4C A CIN CO S VDD VSS
MM7 net85 A net88 VNW P12LL W=440.00n L=60.00n
MM32 net35 CIN VDD VNW P12LL W=430.00n L=60.00n
MM0 CO acinn VDD VNW P12LL W=1.08u L=60.00n
MM6 net88 net35 VDD VNW P12LL W=440.00n L=60.00n
MM10 S net85 VDD VNW P12LL W=1.08u L=60.00n
MM45 acinn net35 VDD VNW P12LL W=440.00n L=60.00n
MM46 acinn A VDD VNW P12LL W=440.00n L=60.00n
MM4 net85 acinn VDD VNW P12LL W=440.00n L=60.00n
MM8 net117 A VSS VPW N12LL W=430.00n L=60.00n
MM9 net117 net35 VSS VPW N12LL W=430.00n L=60.00n
MM1 CO acinn VSS VPW N12LL W=860.00n L=60.00n
MM43 acinn A net_079 VPW N12LL W=510.00n L=60.00n
MM31 net35 CIN VSS VPW N12LL W=350.00n L=60.00n
MM44 net_079 net35 VSS VPW N12LL W=510.00n L=60.00n
MM11 S net85 VSS VPW N12LL W=860.00n L=60.00n
MM5 net85 acinn net117 VPW N12LL W=350.00n L=60.00n
.ENDS ADH1CINHSV4C
****Sub-Circuit for ADH1CONHSV1, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1CONHSV1 A CI CON S VDD VSS
MM45 CON CI VDD VNW P12LL W=390.00n L=60.00n
MM46 CON A VDD VNW P12LL W=390.00n L=60.00n
MM48 net45 CI S VNW P12LL W=440.00n L=60.00n
MM32 net35 CI VDD VNW P12LL W=270.00n L=60.00n
MM29 net45 net46 VDD VNW P12LL W=440.00n L=60.00n
MM28 net46 A VDD VNW P12LL W=440.00n L=60.00n
MM39 net46 net35 S VNW P12LL W=440.00n L=60.00n
MM27 net46 A VSS VPW N12LL W=350.00n L=60.00n
MM47 net45 net35 S VPW N12LL W=350.00n L=60.00n
MM30 net45 net46 VSS VPW N12LL W=350.00n L=60.00n
MM43 CON A net_95 VPW N12LL W=430.00n L=60.00n
MM31 net35 CI VSS VPW N12LL W=220.00n L=60.00n
MM44 net_95 CI VSS VPW N12LL W=430.00n L=60.00n
MM36 net46 CI S VPW N12LL W=350.00n L=60.00n
.ENDS ADH1CONHSV1
****Sub-Circuit for ADH1CONHSV1C, Thu May 19 13:57:40 CST 2011****
.SUBCKT ADH1CONHSV1C A B CON S VDD VSS
MM7 net85 A net88 VNW P12LL W=200.00n L=60.00n
MM6 net88 B VDD VNW P12LL W=200.00n L=60.00n
MM10 S net85 VDD VNW P12LL W=440.00n L=60.00n
MM1 CON B VDD VNW P12LL W=300.00n L=60.00n
MM0 CON A VDD VNW P12LL W=300.00n L=60.00n
MM4 net85 CON VDD VNW P12LL W=200.00n L=60.00n
MM8 net117 A VSS VPW N12LL W=250.00n L=60.00n
MM9 net117 B VSS VPW N12LL W=250.00n L=60.00n
MM11 S net85 VSS VPW N12LL W=350.00n L=60.00n
MM2 net125 B VSS VPW N12LL W=350.00n L=60.00n
MM5 net85 CON net117 VPW N12LL W=180.00n L=60.00n
MM3 CON A net125 VPW N12LL W=350.00n L=60.00n
.ENDS ADH1CONHSV1C
****Sub-Circuit for ADH1CONHSV2, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1CONHSV2 A CI CON S VDD VSS
MM36 net46 CI S VPW N12LL W=430.00n L=60.00n
MM27 net46 A VSS VPW N12LL W=430.00n L=60.00n
MM30 net45 net46 VSS VPW N12LL W=430.00n L=60.00n
MM31 net35 CI VSS VPW N12LL W=220.00n L=60.00n
MM47 net45 net35 S VPW N12LL W=430.00n L=60.00n
MM44 net_43 CI VSS VPW N12LL W=430.00n L=60.00n
MM43 CON A net_43 VPW N12LL W=430.00n L=60.00n
MM28 net46 A VDD VNW P12LL W=540.00n L=60.00n
MM29 net45 net46 VDD VNW P12LL W=540.00n L=60.00n
MM48 net45 CI S VNW P12LL W=540.00n L=60.00n
MM46 CON A VDD VNW P12LL W=420.00n L=60.00n
MM32 net35 CI VDD VNW P12LL W=270.00n L=60.00n
MM45 CON CI VDD VNW P12LL W=420.00n L=60.00n
MM39 net46 net35 S VNW P12LL W=540.00n L=60.00n
.ENDS ADH1CONHSV2
****Sub-Circuit for ADH1CONHSV2C, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT ADH1CONHSV2C A B CON S VDD VSS
MM2 net81 B VSS VPW N12LL W=430.00n L=60.00n
MM5 net125 CON net97 VPW N12LL W=180.00n L=60.00n
MM3 CON A net81 VPW N12LL W=430.00n L=60.00n
MM8 net97 A VSS VPW N12LL W=320.00n L=60.00n
MM9 net97 B VSS VPW N12LL W=320.00n L=60.00n
MM11 S net125 VSS VPW N12LL W=430.00n L=60.00n
MM7 net125 A net128 VNW P12LL W=220.00n L=60.00n
MM6 net128 B VDD VNW P12LL W=220.00n L=60.00n
MM10 S net125 VDD VNW P12LL W=540.00n L=60.00n
MM1 CON B VDD VNW P12LL W=370.00n L=60.00n
MM0 CON A VDD VNW P12LL W=370.00n L=60.00n
MM4 net125 CON VDD VNW P12LL W=220.00n L=60.00n
.ENDS ADH1CONHSV2C
****Sub-Circuit for ADH1CONHSV4, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1CONHSV4 A CI CON S VDD VSS
MM28 net46 A VDD VNW P12LL W=1.08u L=60.00n
MM29 net45 net46 VDD VNW P12LL W=1.08u L=60.00n
MM48 net45 CI S VNW P12LL W=1.08u L=60.00n
MM46 CON A VDD VNW P12LL W=960.00n L=60.00n
MM32 net35 CI VDD VNW P12LL W=430.00n L=60.00n
MM45 CON CI VDD VNW P12LL W=960.00n L=60.00n
MM39 net46 net35 S VNW P12LL W=1.08u L=60.00n
MM44 net_71 CI VSS VPW N12LL W=860n L=60.00n
MM30 net45 net46 VSS VPW N12LL W=860.00n L=60.00n
MM36 net46 CI S VPW N12LL W=860.00n L=60.00n
MM47 net45 net35 S VPW N12LL W=860.00n L=60.00n
MM43 CON A net_71 VPW N12LL W=860n L=60.00n
MM31 net35 CI VSS VPW N12LL W=350.00n L=60.00n
MM27 net46 A VSS VPW N12LL W=860.00n L=60.00n
.ENDS ADH1CONHSV4
****Sub-Circuit for ADH1CONHSV4C, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT ADH1CONHSV4C A B CON S VDD VSS
MM7 net97 A net100 VNW P12LL W=440.00n L=60.00n
MM6 net100 B VDD VNW P12LL W=440.00n L=60.00n
MM10 S net97 VDD VNW P12LL W=1.08u L=60.00n
MM1 CON B VDD VNW P12LL W=740n L=60.00n
MM0 CON A VDD VNW P12LL W=740n L=60.00n
MM4 net97 CON VDD VNW P12LL W=440.00n L=60.00n
MM2 net121 B VSS VPW N12LL W=860.00n L=60.00n
MM5 net97 CON net109 VPW N12LL W=350.00n L=60.00n
MM3 CON A net121 VPW N12LL W=860.00n L=60.00n
MM8 net109 A VSS VPW N12LL W=430.00n L=60.00n
MM9 net109 B VSS VPW N12LL W=430.00n L=60.00n
MM11 S net97 VSS VPW N12LL W=860.00n L=60.00n
.ENDS ADH1CONHSV4C
****Sub-Circuit for ADH1CSCINHSV1, Mon Apr 11 16:55:11 CST 2011****
.SUBCKT ADH1CSCINHSV1 A CIN CO CS S VDD VSS
MM4 an cinn net172 VNW P12LL W=350n L=60.00n
MM6 net135 an VDD VNW P12LL W=270n L=60.00n
MM7 net172 CIN net135 VNW P12LL W=270n L=60.00n
MM0 cinn CIN VDD VNW P12LL W=440n L=60.00n
MM10 net123 an VDD VNW P12LL W=280n L=60.00n
MM11 CO CIN net123 VNW P12LL W=280n L=60.00n
MM48 net172 csn net163 VNW P12LL W=350n L=60.00n
MM32 csn CS VDD VNW P12LL W=270n L=60.00n
MM28 an A VDD VNW P12LL W=440n L=60.00n
MM39 an CS net163 VNW P12LL W=300n L=60.00n
MM2 S net163 VDD VNW P12LL W=440n L=60.00n
MM9 net180 an VSS VPW N12LL W=220.00n L=60.00n
MM8 net172 cinn net180 VPW N12LL W=220.00n L=60.00n
MM43 CO an VSS VPW N12LL W=220.00n L=60.00n
MM47 net172 CS net163 VPW N12LL W=280.00n L=60.00n
MM31 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM27 an A VSS VPW N12LL W=350.00n L=60.00n
MM36 an csn net163 VPW N12LL W=240.00n L=60.00n
MM3 S net163 VSS VPW N12LL W=350.00n L=60.00n
MM1 cinn CIN VSS VPW N12LL W=350.00n L=60.00n
MM44 CO CIN VSS VPW N12LL W=220.00n L=60.00n
MM5 an CIN net172 VPW N12LL W=280.00n L=60.00n
.ENDS ADH1CSCINHSV1
****Sub-Circuit for ADH1CSCINHSV2, Mon Apr 11 16:55:11 CST 2011****
.SUBCKT ADH1CSCINHSV2 A CIN CO CS S VDD VSS
MM5 na CIN net96 VPW N12LL W=350.00n L=60.00n
MM9 net100 na VSS VPW N12LL W=220.00n L=60.00n
MM1 cinn CIN VSS VPW N12LL W=430.00n L=60.00n
MM8 net96 cinn net100 VPW N12LL W=220.00n L=60.00n
MM43 CO na VSS VPW N12LL W=220.00n L=60.00n
MM44 CO CIN VSS VPW N12LL W=220.00n L=60.00n
MM47 net96 CS net123 VPW N12LL W=350.00n L=60.00n
MM31 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM27 na A VSS VPW N12LL W=430.00n L=60.00n
MM36 na csn net123 VPW N12LL W=280.00n L=60.00n
MM3 S net123 VSS VPW N12LL W=430.00n L=60.00n
MM4 na cinn net96 VNW P12LL W=440.00n L=60.00n
MM6 net144 na VDD VNW P12LL W=275.00n L=60.00n
MM7 net96 CIN net144 VNW P12LL W=275.00n L=60.00n
MM0 cinn CIN VDD VNW P12LL W=540n L=60.00n
MM10 net151 na VDD VNW P12LL W=280.00n L=60.00n
MM11 CO CIN net151 VNW P12LL W=280.00n L=60.00n
MM48 net96 csn net123 VNW P12LL W=440.00n L=60.00n
MM32 csn CS VDD VNW P12LL W=275.00n L=60.00n
MM28 na A VDD VNW P12LL W=540n L=60.00n
MM39 na CS net123 VNW P12LL W=350.00n L=60.00n
MM2 S net123 VDD VNW P12LL W=540n L=60.00n
.ENDS ADH1CSCINHSV2
****Sub-Circuit for ADH1CSCINHSV4, Mon Apr 11 16:55:11 CST 2011****
.SUBCKT ADH1CSCINHSV4 A CIN CO CS S VDD VSS
MM3 S net127 VSS VPW N12LL W=860.00n L=60.00n
MM36 an csn net127 VPW N12LL W=350.00n L=60.00n
MM27 an A VSS VPW N12LL W=430.00n L=60.00n
MM31 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM47 net112 CS net127 VPW N12LL W=430.00n L=60.00n
MM44 CO CIN VSS VPW N12LL W=240.00n L=60.00n
MM43 CO an VSS VPW N12LL W=240.00n L=60.00n
MM8 net112 cinn net104 VPW N12LL W=220.00n L=60.00n
MM1 cinn CIN VSS VPW N12LL W=430.00n L=60.00n
MM9 net104 an VSS VPW N12LL W=220.00n L=60.00n
MM5 an CIN net112 VPW N12LL W=430.00n L=60.00n
MM2 S net127 VDD VNW P12LL W=1.08u L=60.00n
MM39 an CS net127 VNW P12LL W=440.00n L=60.00n
MM28 an A VDD VNW P12LL W=540n L=60.00n
MM32 csn CS VDD VNW P12LL W=275.00n L=60.00n
MM48 net112 csn net127 VNW P12LL W=540.00n L=60.00n
MM11 CO CIN net167 VNW P12LL W=320.00n L=60.00n
MM10 net167 an VDD VNW P12LL W=320.00n L=60.00n
MM0 cinn CIN VDD VNW P12LL W=540n L=60.00n
MM7 net112 CIN net155 VNW P12LL W=275.00n L=60.00n
MM6 net155 an VDD VNW P12LL W=275.00n L=60.00n
MM4 an cinn net112 VNW P12LL W=540.00n L=60.00n
.ENDS ADH1CSCINHSV4
****Sub-Circuit for ADH1CSCONHSV1, Mon Apr 11 14:38:06 CST 2011****
.SUBCKT ADH1CSCONHSV1 A CI CON CS S VDD VSS
MM8 net119 an VDD VNW P12LL W=270.00n L=60.00n
MM4 an CI net156 VNW P12LL W=350.00n L=60.00n
MM6 net156 cin net119 VNW P12LL W=270.00n L=60.00n
MM0 cin CI VDD VNW P12LL W=440n L=60.00n
MM48 net156 csn net147 VNW P12LL W=350.00n L=60.00n
MM32 csn CS VDD VNW P12LL W=270.00n L=60.00n
MM28 an A VDD VNW P12LL W=440n L=60.00n
MM39 an CS net147 VNW P12LL W=300.00n L=60.00n
MM45 CON CI VDD VNW P12LL W=220.00n L=60.00n
MM2 S net147 VDD VNW P12LL W=440n L=60.00n
MM46 CON A VDD VNW P12LL W=220.00n L=60.00n
MM5 an cin net156 VPW N12LL W=280.00n L=60.00n
MM1 cin CI VSS VPW N12LL W=350.00n L=60.00n
MM9 net164 an VSS VPW N12LL W=220.00n L=60.00n
MM7 net156 CI net164 VPW N12LL W=220.00n L=60.00n
MM43 CON CI net148 VPW N12LL W=250.00n L=60.00n
MM44 net148 A VSS VPW N12LL W=250.00n L=60.00n
MM47 net156 CS net147 VPW N12LL W=280.00n L=60.00n
MM31 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM27 an A VSS VPW N12LL W=350.00n L=60.00n
MM36 an csn net147 VPW N12LL W=240.00n L=60.00n
MM3 S net147 VSS VPW N12LL W=350.00n L=60.00n
.ENDS ADH1CSCONHSV1
****Sub-Circuit for ADH1CSCONHSV2, Mon Apr 11 14:38:06 CST 2011****
.SUBCKT ADH1CSCONHSV2 A CI CON CS S VDD VSS
MM5 an cin net92 VPW N12LL W=350.00n L=60.00n
MM9 net_098 an VSS VPW N12LL W=220.00n L=60.00n
MM1 cin CI VSS VPW N12LL W=425.00n L=60.00n
MM7 net92 CI net_098 VPW N12LL W=220.00n L=60.00n
MM43 CON CI net_0137 VPW N12LL W=250.00n L=60.00n
MM44 net_0137 A VSS VPW N12LL W=250.00n L=60.00n
MM47 net92 CS net_0144 VPW N12LL W=350.00n L=60.00n
MM31 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM27 an A VSS VPW N12LL W=430.00n L=60.00n
MM36 an csn net_0144 VPW N12LL W=280.00n L=60.00n
MM3 S net_0144 VSS VPW N12LL W=430.00n L=60.00n
MM8 net_0145 an VDD VNW P12LL W=270.00n L=60.00n
MM4 an CI net92 VNW P12LL W=440.00n L=60.00n
MM6 net92 cin net_0145 VNW P12LL W=270.00n L=60.00n
MM0 cin CI VDD VNW P12LL W=540n L=60.00n
MM48 net92 csn net_0144 VNW P12LL W=440.00n L=60.00n
MM32 csn CS VDD VNW P12LL W=270.00n L=60.00n
MM28 an A VDD VNW P12LL W=540n L=60.00n
MM39 an CS net_0144 VNW P12LL W=350.00n L=60.00n
MM45 CON CI VDD VNW P12LL W=220.00n L=60.00n
MM2 S net_0144 VDD VNW P12LL W=540n L=60.00n
MM46 CON A VDD VNW P12LL W=220.00n L=60.00n
.ENDS ADH1CSCONHSV2
****Sub-Circuit for ADH1CSCONHSV4, Mon Apr 11 14:38:06 CST 2011****
.SUBCKT ADH1CSCONHSV4 A CI CON CS S VDD VSS
MM8 net119 an VDD VNW P12LL W=270.00n L=60.00n
MM4 an CI net156 VNW P12LL W=540.00n L=60.00n
MM6 net156 cin net119 VNW P12LL W=270.00n L=60.00n
MM0 cin CI VDD VNW P12LL W=540n L=60.00n
MM48 net156 csn net147 VNW P12LL W=540.00n L=60.00n
MM32 csn CS VDD VNW P12LL W=270.00n L=60.00n
MM28 an A VDD VNW P12LL W=540n L=60.00n
MM39 an CS net147 VNW P12LL W=440.00n L=60.00n
MM45 CON CI VDD VNW P12LL W=310.00n L=60.00n
MM2 S net147 VDD VNW P12LL W=1.08u L=60.00n
MM46 CON A VDD VNW P12LL W=310.00n L=60.00n
MM5 an cin net156 VPW N12LL W=430.00n L=60.00n
MM9 net164 an VSS VPW N12LL W=220.00n L=60.00n
MM1 cin CI VSS VPW N12LL W=425.00n L=60.00n
MM7 net156 CI net164 VPW N12LL W=220.00n L=60.00n
MM43 CON CI net148 VPW N12LL W=350.00n L=60.00n
MM44 net148 A VSS VPW N12LL W=350.00n L=60.00n
MM47 net156 CS net147 VPW N12LL W=430.00n L=60.00n
MM31 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM27 an A VSS VPW N12LL W=430.00n L=60.00n
MM36 an csn net147 VPW N12LL W=350.00n L=60.00n
MM3 S net147 VSS VPW N12LL W=860.00n L=60.00n
.ENDS ADH1CSCONHSV4
****Sub-Circuit for ADH1HSV1, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT ADH1HSV1 A B CO S VDD VSS
MM43 net_0163 B net_0135 VPW N12LL W=260.00n L=60.00n
MM44 net_0135 A VSS VPW N12LL W=260.00n L=60.00n
MM47 net45 net35 S VPW N12LL W=300.00n L=60.00n
MM31 net35 B VSS VPW N12LL W=330.00n L=60.00n
MM30 net45 net46 VSS VPW N12LL W=300.00n L=60.00n
MM27 net46 A VSS VPW N12LL W=430.00n L=60.00n
MM22 CO net_0163 VSS VPW N12LL W=300.00n L=60.00n
MM36 net46 B S VPW N12LL W=300.00n L=60.00n
MM45 net_0163 A VDD VNW P12LL W=300.00n L=60.00n
MM46 net_0163 B VDD VNW P12LL W=300.00n L=60.00n
MM48 net45 B S VNW P12LL W=450.00n L=60.00n
MM32 net35 B VDD VNW P12LL W=500.00n L=60.00n
MM29 net45 net46 VDD VNW P12LL W=450.00n L=60.00n
MM28 net46 A VDD VNW P12LL W=650n L=60.00n
MM21 CO net_0163 VDD VNW P12LL W=450.00n L=60.00n
MM39 net46 net35 S VNW P12LL W=450.00n L=60.00n
.ENDS ADH1HSV1
****Sub-Circuit for ADH1HSV1C, Thu May 19 13:57:40 CST 2011****
.SUBCKT ADH1HSV1C A B CO S VDD VSS
MM7 net85 A net88 VNW P12LL W=200.00n L=60.00n
MM6 net88 B VDD VNW P12LL W=200.00n L=60.00n
MM10 S net85 VDD VNW P12LL W=440.00n L=60.00n
MM1 abn B VDD VNW P12LL W=300.00n L=60.00n
MM0 abn A VDD VNW P12LL W=300.00n L=60.00n
MM12 CO abn VDD VNW P12LL W=440.00n L=60.00n
MM4 net85 abn VDD VNW P12LL W=200.00n L=60.00n
MM8 net117 A VSS VPW N12LL W=250.00n L=60.00n
MM9 net117 B VSS VPW N12LL W=250.00n L=60.00n
MM11 S net85 VSS VPW N12LL W=350.00n L=60.00n
MM13 CO abn VSS VPW N12LL W=350.00n L=60.00n
MM2 net125 B VSS VPW N12LL W=350.00n L=60.00n
MM5 net85 abn net117 VPW N12LL W=180.00n L=60.00n
MM3 abn A net125 VPW N12LL W=350.00n L=60.00n
.ENDS ADH1HSV1C
****Sub-Circuit for ADH1HSV2, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT ADH1HSV2 A B CO S VDD VSS
MM43 net_0163 B net_0135 VPW N12LL W=260.00n L=60.00n
MM44 net_0135 A VSS VPW N12LL W=260.00n L=60.00n
MM47 net45 net35 S VPW N12LL W=430.00n L=60.00n
MM31 net35 B VSS VPW N12LL W=500.00n L=60.00n
MM30 net45 net46 VSS VPW N12LL W=430.00n L=60.00n
MM27 net46 A VSS VPW N12LL W=560.00n L=60.00n
MM22 CO net_0163 VSS VPW N12LL W=430.00n L=60.00n
MM36 net46 B S VPW N12LL W=430.00n L=60.00n
MM45 net_0163 A VDD VNW P12LL W=300.00n L=60.00n
MM46 net_0163 B VDD VNW P12LL W=300.00n L=60.00n
MM48 net45 B S VNW P12LL W=640.00n L=60.00n
MM32 net35 B VDD VNW P12LL W=760.00n L=60.00n
MM29 net45 net46 VDD VNW P12LL W=650.00n L=60.00n
MM28 net46 A VDD VNW P12LL W=860n L=60.00n
MM21 CO net_0163 VDD VNW P12LL W=650.00n L=60.00n
MM39 net46 net35 S VNW P12LL W=645.00n L=60.00n
.ENDS ADH1HSV2
****Sub-Circuit for ADH1HSV2C, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1HSV2C A B CO S VDD VSS
MM13 CO abn VSS VPW N12LL W=430.00n L=60.00n
MM2 net81 B VSS VPW N12LL W=430.00n L=60.00n
MM5 net125 abn net97 VPW N12LL W=180.00n L=60.00n
MM3 abn A net81 VPW N12LL W=430.00n L=60.00n
MM8 net97 A VSS VPW N12LL W=320.00n L=60.00n
MM9 net97 B VSS VPW N12LL W=320.00n L=60.00n
MM11 S net125 VSS VPW N12LL W=430.00n L=60.00n
MM7 net125 A net128 VNW P12LL W=220.00n L=60.00n
MM6 net128 B VDD VNW P12LL W=220.00n L=60.00n
MM10 S net125 VDD VNW P12LL W=540.00n L=60.00n
MM1 abn B VDD VNW P12LL W=370.00n L=60.00n
MM0 abn A VDD VNW P12LL W=370.00n L=60.00n
MM12 CO abn VDD VNW P12LL W=540.00n L=60.00n
MM4 net125 abn VDD VNW P12LL W=220.00n L=60.00n
.ENDS ADH1HSV2C
****Sub-Circuit for ADH1HSV4, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT ADH1HSV4 A B CO S VDD VSS
MM43 net_0163 B net_0135 VPW N12LL W=430.00n L=60.00n
MM44 net_0135 A VSS VPW N12LL W=420.00n L=60.00n
MM47 net45 net35 S VPW N12LL W=390.00n L=60.00n
MM31 net35 B VSS VPW N12LL W=990.00n L=60.00n
MM30 net45 net46 VSS VPW N12LL W=860.00n L=60.00n
MM27 net46 A VSS VPW N12LL W=1.12u L=60.00n
MM22 CO net_0163 VSS VPW N12LL W=860.00n L=60.00n
MM36 net46 B S VPW N12LL W=380.00n L=60.00n
MM45 net_0163 A VDD VNW P12LL W=500.00n L=60.00n
MM46 net_0163 B VDD VNW P12LL W=500.00n L=60.00n
MM48 net45 B S VNW P12LL W=1.22u L=60.00n
MM32 net35 B VDD VNW P12LL W=1.52u L=60.00n
MM29 net45 net46 VDD VNW P12LL W=1.3u L=60.00n
MM28 net46 A VDD VNW P12LL W=1.72u L=60.00n
MM21 CO net_0163 VDD VNW P12LL W=1.3u L=60.00n
MM39 net46 net35 S VNW P12LL W=1.22u L=60.00n
.ENDS ADH1HSV4
****Sub-Circuit for ADH1HSV4C, Thu Jan 20 09:48:40 CST 2011****
.SUBCKT ADH1HSV4C A B CO S VDD VSS
MM7 net97 A net100 VNW P12LL W=440.00n L=60.00n
MM6 net100 B VDD VNW P12LL W=440.00n L=60.00n
MM10 S net97 VDD VNW P12LL W=1.08u L=60.00n
MM1 abn B VDD VNW P12LL W=740n L=60.00n
MM12 CO abn VDD VNW P12LL W=1.08u L=60.00n
MM0 abn A VDD VNW P12LL W=740n L=60.00n
MM4 net97 abn VDD VNW P12LL W=440.00n L=60.00n
MM13 CO abn VSS VPW N12LL W=860.00n L=60.00n
MM2 net121 B VSS VPW N12LL W=860.00n L=60.00n
MM5 net97 abn net109 VPW N12LL W=350.00n L=60.00n
MM3 abn A net121 VPW N12LL W=860.00n L=60.00n
MM8 net109 A VSS VPW N12LL W=430.00n L=60.00n
MM9 net109 B VSS VPW N12LL W=430.00n L=60.00n
MM11 S net97 VSS VPW N12LL W=860.00n L=60.00n
.ENDS ADH1HSV4C
****Sub-Circuit for ADH2CONHSV1, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT ADH2CONHSV1 A B CO0N CO1N CS S VDD VSS
MM14 xo csn net82 VNW P12LL W=220.00n L=60.00n
MM15 xn CS net82 VNW P12LL W=220.00n L=60.00n
MM16 xn xo VDD VNW P12LL W=220.00n L=60.00n
MM17 net18 B VDD VNW P12LL W=550.00n L=60.00n
MM18 xo CO1N net18 VNW P12LL W=440.00n L=60.00n
MM21 net18 A VDD VNW P12LL W=550.00n L=60.00n
MM22 S net82 VDD VNW P12LL W=440.00n L=60.00n
MM5 net50 B VDD VNW P12LL W=550.00n L=60.00n
MM4 CO1N A net50 VNW P12LL W=550.00n L=60.00n
MM28 csn CS VDD VNW P12LL W=220.00n L=60.00n
MM13 CO0N B VDD VNW P12LL W=180.00n L=60.00n
MM12 CO0N A VDD VNW P12LL W=180.00n L=60.00n
MM23 xo CS net82 VPW N12LL W=180.00n L=60.00n
MM24 xn csn net82 VPW N12LL W=180.00n L=60.00n
MM25 S net82 VSS VPW N12LL W=350.00n L=60.00n
MM26 xn xo VSS VPW N12LL W=180.00n L=60.00n
MM29 net63 B VSS VPW N12LL W=430.00n L=60.00n
MM30 xo A net63 VPW N12LL W=430.00n L=60.00n
MM31 xo CO1N VSS VPW N12LL W=390.00n L=60.00n
MM27 csn CS VSS VPW N12LL W=180.00n L=60.00n
MM11 CO0N A net83 VPW N12LL W=210.00n L=60.00n
MM10 net83 B VSS VPW N12LL W=210.00n L=60.00n
MM2 CO1N B VSS VPW N12LL W=300.00n L=60.00n
MM3 CO1N A VSS VPW N12LL W=300.00n L=60.00n
.ENDS ADH2CONHSV1
****Sub-Circuit for ADH2CONHSV2, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT ADH2CONHSV2 A B CO0N CO1N CS S VDD VSS
MM14 xo csn net82 VNW P12LL W=270.00n L=60.00n
MM15 xn CS net82 VNW P12LL W=270.00n L=60.00n
MM16 xn xo VDD VNW P12LL W=270.00n L=60.00n
MM17 net18 B VDD VNW P12LL W=650.00n L=60.00n
MM18 xo CO1N net18 VNW P12LL W=540.00n L=60.00n
MM21 net18 A VDD VNW P12LL W=650.00n L=60.00n
MM22 S net82 VDD VNW P12LL W=540.00n L=60.00n
MM5 net50 B VDD VNW P12LL W=650.00n L=60.00n
MM4 CO1N A net50 VNW P12LL W=650.00n L=60.00n
MM28 csn CS VDD VNW P12LL W=270.00n L=60.00n
MM13 CO0N B VDD VNW P12LL W=220.00n L=60.00n
MM12 CO0N A VDD VNW P12LL W=220.00n L=60.00n
MM23 xo CS net82 VPW N12LL W=220.00n L=60.00n
MM24 xn csn net82 VPW N12LL W=220.00n L=60.00n
MM25 S net82 VSS VPW N12LL W=430.00n L=60.00n
MM26 xn xo VSS VPW N12LL W=220.00n L=60.00n
MM29 net63 B VSS VPW N12LL W=430.00n L=60.00n
MM30 xo A net63 VPW N12LL W=430.00n L=60.00n
MM31 xo CO1N VSS VPW N12LL W=430.00n L=60.00n
MM27 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM11 CO0N A net83 VPW N12LL W=260.00n L=60.00n
MM10 net83 B VSS VPW N12LL W=260.00n L=60.00n
MM2 CO1N B VSS VPW N12LL W=350.00n L=60.00n
MM3 CO1N A VSS VPW N12LL W=350.00n L=60.00n
.ENDS ADH2CONHSV2
****Sub-Circuit for ADH2CONHSV4, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT ADH2CONHSV4 A B CO0N CO1N CS S VDD VSS
MM14 xo csn net82 VNW P12LL W=540.00n L=60.00n
MM15 xn CS net82 VNW P12LL W=540.00n L=60.00n
MM16 xn xo VDD VNW P12LL W=540.00n L=60.00n
MM17 net18 B VDD VNW P12LL W=1.3u L=60.00n
MM18 xo CO1N net18 VNW P12LL W=1.08u L=60.00n
MM21 net18 A VDD VNW P12LL W=1.3u L=60.00n
MM22 S net82 VDD VNW P12LL W=1.08u L=60.00n
MM5 net50 B VDD VNW P12LL W=1.3u L=60.00n
MM4 CO1N A net50 VNW P12LL W=1.3u L=60.00n
MM28 csn CS VDD VNW P12LL W=270.00n L=60.00n
MM13 CO0N B VDD VNW P12LL W=440.00n L=60.00n
MM12 CO0N A VDD VNW P12LL W=440.00n L=60.00n
MM23 xo CS net82 VPW N12LL W=430.00n L=60.00n
MM24 xn csn net82 VPW N12LL W=430.00n L=60.00n
MM25 S net82 VSS VPW N12LL W=860.00n L=60.00n
MM26 xn xo VSS VPW N12LL W=430.00n L=60.00n
MM29 net63 B VSS VPW N12LL W=1.08u L=60.00n
MM30 xo A net63 VPW N12LL W=1.08u L=60.00n
MM31 xo CO1N VSS VPW N12LL W=880.00n L=60.00n
MM27 csn CS VSS VPW N12LL W=220.00n L=60.00n
MM11 CO0N A net83 VPW N12LL W=430.00n L=60.00n
MM10 net83 B VSS VPW N12LL W=430.00n L=60.00n
MM2 CO1N B VSS VPW N12LL W=700.00n L=60.00n
MM3 CO1N A VSS VPW N12LL W=700.00n L=60.00n
.ENDS ADH2CONHSV4
****Sub-Circuit for AND2HSV0, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND2HSV0 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=200.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=300.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS AND2HSV0
****Sub-Circuit for AND2HSV0RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV0RD A1 A2 Z VDD VSS
MM4 Z net12 VDD VNW P12LL W=250n L=60n
MM2 net12 A2 VDD VNW P12LL W=200n L=60n
MM1 net12 A1 VDD VNW P12LL W=200n L=60n
MM5 Z net12 VSS VPW N12LL W=200n L=60n
MM3 net12 A2 net046 VPW N12LL W=200n L=60n
MM0 net046 A1 VSS VPW N12LL W=200n L=60n
.ENDS AND2HSV0RD
****Sub-Circuit for AND2HSV1, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND2HSV1 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=200.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=440.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS AND2HSV1
****Sub-Circuit for AND2HSV12, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV12 A1 A2 Z VDD VSS
MM0 net4 A1 VSS VPW N12LL W=1.29u L=60n
MM3 net16 A2 net4 VPW N12LL W=1.29u L=60n
MM5 Z net16 VSS VPW N12LL W=2.58u L=60n
MM1 net16 A1 VDD VNW P12LL W=1.32u L=60n
MM2 net16 A2 VDD VNW P12LL W=1.32u L=60n
MM4 Z net16 VDD VNW P12LL W=3.24u L=60n
.ENDS AND2HSV12
****Sub-Circuit for AND2HSV12RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV12RD A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=2.1u L=60n
MM0 net057 A1 VSS VPW N12LL W=2.1u L=60n
MM5 Z net16 VSS VPW N12LL W=2.58u L=60n
MM1 net16 A1 VDD VNW P12LL W=2.1u L=60n
MM2 net16 A2 VDD VNW P12LL W=2.1u L=60n
MM4 Z net16 VDD VNW P12LL W=3.24u L=60n
.ENDS AND2HSV12RD
****Sub-Circuit for AND2HSV12RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV12RQ A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=650n L=60n
MM0 net057 A1 VSS VPW N12LL W=650n L=60n
MM5 Z net16 VSS VPW N12LL W=2.58u L=60n
MM1 net16 A1 VDD VNW P12LL W=810n L=60n
MM2 net16 A2 VDD VNW P12LL W=810n L=60n
MM4 Z net16 VDD VNW P12LL W=3.24u L=60n
.ENDS AND2HSV12RQ
****Sub-Circuit for AND2HSV16, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV16 A1 A2 Z VDD VSS
MM0 net4 A1 VSS VPW N12LL W=1.72u L=60n
MM3 net16 A2 net4 VPW N12LL W=1.72u L=60n
MM5 Z net16 VSS VPW N12LL W=3.44u L=60n
MM1 net16 A1 VDD VNW P12LL W=1.76u L=60n
MM2 net16 A2 VDD VNW P12LL W=1.76u L=60n
MM4 Z net16 VDD VNW P12LL W=4.32u L=60n
.ENDS AND2HSV16
****Sub-Circuit for AND2HSV16RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV16RD A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=2.8u L=60n
MM0 net057 A1 VSS VPW N12LL W=2.8u L=60n
MM5 Z net16 VSS VPW N12LL W=3.44u L=60n
MM1 net16 A1 VDD VNW P12LL W=2.8u L=60n
MM2 net16 A2 VDD VNW P12LL W=2.8u L=60n
MM4 Z net16 VDD VNW P12LL W=4.32u L=60n
.ENDS AND2HSV16RD
****Sub-Circuit for AND2HSV16RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV16RQ A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=860n L=60n
MM0 net057 A1 VSS VPW N12LL W=860n L=60n
MM5 Z net16 VSS VPW N12LL W=3.44u L=60n
MM1 net16 A1 VDD VNW P12LL W=1.08u L=60n
MM2 net16 A2 VDD VNW P12LL W=1.08u L=60n
MM4 Z net16 VDD VNW P12LL W=4.32u L=60n
.ENDS AND2HSV16RQ
****Sub-Circuit for AND2HSV1RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV1RD A1 A2 Z VDD VSS
MM3 net16 A2 net030 VPW N12LL W=280n L=60n
MM0 net030 A1 VSS VPW N12LL W=280n L=60n
MM5 Z net16 VSS VPW N12LL W=350n L=60n
MM1 net16 A1 VDD VNW P12LL W=280n L=60n
MM2 net16 A2 VDD VNW P12LL W=280n L=60n
MM4 Z net16 VDD VNW P12LL W=440n L=60n
.ENDS AND2HSV1RD
****Sub-Circuit for AND2HSV2, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND2HSV2 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=200.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=650.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.0n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.0n L=60.00n
.ENDS AND2HSV2
****Sub-Circuit for AND2HSV20, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV20 A1 A2 Z VDD VSS
MM0 net4 A1 VSS VPW N12LL W=2.15u L=60n
MM3 net16 A2 net4 VPW N12LL W=2.15u L=60n
MM5 Z net16 VSS VPW N12LL W=4.3u L=60n
MM1 net16 A1 VDD VNW P12LL W=2.2u L=60n
MM2 net16 A2 VDD VNW P12LL W=2.2u L=60n
MM4 Z net16 VDD VNW P12LL W=5.4u L=60n
.ENDS AND2HSV20
****Sub-Circuit for AND2HSV20RD, Thu May 19 15:57:34 CST 2011****
.SUBCKT AND2HSV20RD A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=3.44u L=60n
MM0 net057 A1 VSS VPW N12LL W=3.44u L=60n
MM5 Z net16 VSS VPW N12LL W=4.3u L=60n
MM1 net16 A1 VDD VNW P12LL W=3.5u L=60n
MM2 net16 A2 VDD VNW P12LL W=3.5u L=60n
MM4 Z net16 VDD VNW P12LL W=5.4u L=60n
.ENDS AND2HSV20RD
****Sub-Circuit for AND2HSV20RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV20RQ A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=1.08u L=60n
MM0 net057 A1 VSS VPW N12LL W=1.08u L=60n
MM5 Z net16 VSS VPW N12LL W=4.3u L=60n
MM1 net16 A1 VDD VNW P12LL W=1.35u L=60n
MM2 net16 A2 VDD VNW P12LL W=1.35u L=60n
MM4 Z net16 VDD VNW P12LL W=5.4u L=60n
.ENDS AND2HSV20RQ
****Sub-Circuit for AND2HSV24, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV24 A1 A2 Z VDD VSS
MM0 net4 A1 VSS VPW N12LL W=2.58u L=60n
MM3 net16 A2 net4 VPW N12LL W=2.58u L=60n
MM5 Z net16 VSS VPW N12LL W=5.16u L=60n
MM1 net16 A1 VDD VNW P12LL W=2.64u L=60n
MM2 net16 A2 VDD VNW P12LL W=2.64u L=60n
MM4 Z net16 VDD VNW P12LL W=6.48u L=60n
.ENDS AND2HSV24
****Sub-Circuit for AND2HSV24RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV24RD A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=4.2u L=60n
MM0 net057 A1 VSS VPW N12LL W=4.2u L=60n
MM5 Z net16 VSS VPW N12LL W=5.16u L=60n
MM1 net16 A1 VDD VNW P12LL W=4.2u L=60n
MM2 net16 A2 VDD VNW P12LL W=4.2u L=60n
MM4 Z net16 VDD VNW P12LL W=6.48u L=60n
.ENDS AND2HSV24RD
****Sub-Circuit for AND2HSV24RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV24RQ A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=1.29u L=60n
MM0 net057 A1 VSS VPW N12LL W=1.29u L=60n
MM5 Z net16 VSS VPW N12LL W=5.16u L=60n
MM1 net16 A1 VDD VNW P12LL W=1.62u L=60n
MM2 net16 A2 VDD VNW P12LL W=1.62u L=60n
MM4 Z net16 VDD VNW P12LL W=6.48u L=60n
.ENDS AND2HSV24RQ
****Sub-Circuit for AND2HSV2RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV2RD A1 A2 Z VDD VSS
MM3 net16 A2 net030 VPW N12LL W=350n L=60n
MM0 net030 A1 VSS VPW N12LL W=350n L=60n
MM5 Z net16 VSS VPW N12LL W=430n L=60n
MM1 net16 A1 VDD VNW P12LL W=350n L=60n
MM2 net16 A2 VDD VNW P12LL W=350n L=60n
MM4 Z net16 VDD VNW P12LL W=540n L=60n
.ENDS AND2HSV2RD
****Sub-Circuit for AND2HSV32, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV32 A1 A2 Z VDD VSS
MM0 net4 A1 VSS VPW N12LL W=3.44u L=60n
MM3 net16 A2 net4 VPW N12LL W=3.44u L=60n
MM5 Z net16 VSS VPW N12LL W=6.88u L=60n
MM1 net16 A1 VDD VNW P12LL W=3.52u L=60n
MM2 net16 A2 VDD VNW P12LL W=3.52u L=60n
MM4 Z net16 VDD VNW P12LL W=8.64u L=60n
.ENDS AND2HSV32
****Sub-Circuit for AND2HSV4, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND2HSV4 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=350.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=860.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=350.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=1.3u L=60.00n
MM0 net11 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=520.00n L=60.00n
.ENDS AND2HSV4
****Sub-Circuit for AND2HSV40, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV40 A1 A2 Z VDD VSS
MM0 net4 A1 VSS VPW N12LL W=4.3u L=60n
MM3 net16 A2 net4 VPW N12LL W=4.3u L=60n
MM5 Z net16 VSS VPW N12LL W=8.6u L=60n
MM1 net16 A1 VDD VNW P12LL W=4.4u L=60n
MM2 net16 A2 VDD VNW P12LL W=4.4u L=60n
MM4 Z net16 VDD VNW P12LL W=10.8u L=60n
.ENDS AND2HSV40
****Sub-Circuit for AND2HSV48, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV48 A1 A2 Z VDD VSS
MM0 net4 A1 VSS VPW N12LL W=5.16u L=60n
MM3 net16 A2 net4 VPW N12LL W=5.16u L=60n
MM5 Z net16 VSS VPW N12LL W=10.32u L=60n
MM1 net16 A1 VDD VNW P12LL W=5.28u L=60n
MM2 net16 A2 VDD VNW P12LL W=5.28u L=60n
MM4 Z net16 VDD VNW P12LL W=12.96u L=60n
.ENDS AND2HSV48
****Sub-Circuit for AND2HSV4RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV4RD A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=700n L=60n
MM0 net057 A1 VSS VPW N12LL W=700n L=60n
MM5 Z net16 VSS VPW N12LL W=860n L=60n
MM1 net16 A1 VDD VNW P12LL W=700n L=60n
MM2 net16 A2 VDD VNW P12LL W=700n L=60n
MM4 Z net16 VDD VNW P12LL W=1.08u L=60n
.ENDS AND2HSV4RD
****Sub-Circuit for AND2HSV4RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV4RQ A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=270n L=60n
MM0 net057 A1 VSS VPW N12LL W=270n L=60n
MM5 Z net16 VSS VPW N12LL W=860n L=60n
MM1 net16 A1 VDD VNW P12LL W=270n L=60n
MM2 net16 A2 VDD VNW P12LL W=270n L=60n
MM4 Z net16 VDD VNW P12LL W=1.08u L=60n
.ENDS AND2HSV4RQ
****Sub-Circuit for AND2HSV64, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV64 A1 A2 Z VDD VSS
MM0 net4 A1 VSS VPW N12LL W=6.88u L=60n
MM3 net16 A2 net4 VPW N12LL W=6.88u L=60n
MM5 Z net16 VSS VPW N12LL W=13.76u L=60n
MM1 net16 A1 VDD VNW P12LL W=7.04u L=60n
MM2 net16 A2 VDD VNW P12LL W=7.04u L=60n
MM4 Z net16 VDD VNW P12LL W=17.28u L=60n
.ENDS AND2HSV64
****Sub-Circuit for AND2HSV8, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND2HSV8 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=700.0n L=60.00n
MM2 Z net11 VSS VPW N12LL W=1.72u L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=700.0n L=60.00n
MM3 Z net11 VDD VNW P12LL W=2.6u L=60.00n
MM0 net11 A2 VDD VNW P12LL W=1.04u L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=1.04u L=60.00n
.ENDS AND2HSV8
****Sub-Circuit for AND2HSV8RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV8RD A1 A2 Z VDD VSS
MM3 net16 A2 net030 VPW N12LL W=1.4u L=60n
MM0 net030 A1 VSS VPW N12LL W=1.4u L=60n
MM5 Z net16 VSS VPW N12LL W=1.72u L=60n
MM1 net16 A1 VDD VNW P12LL W=1.4u L=60n
MM2 net16 A2 VDD VNW P12LL W=1.4u L=60n
MM4 Z net16 VDD VNW P12LL W=2.16u L=60n
.ENDS AND2HSV8RD
****Sub-Circuit for AND2HSV8RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND2HSV8RQ A1 A2 Z VDD VSS
MM3 net16 A2 net057 VPW N12LL W=430n L=60n
MM0 net057 A1 VSS VPW N12LL W=430n L=60n
MM5 Z net16 VSS VPW N12LL W=1.72u L=60n
MM1 net16 A1 VDD VNW P12LL W=540n L=60n
MM2 net16 A2 VDD VNW P12LL W=540n L=60n
MM4 Z net16 VDD VNW P12LL W=2.16u L=60n
.ENDS AND2HSV8RQ
****Sub-Circuit for AND3HSV0, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND3HSV0 A1 A2 A3 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=200.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=200.00n L=60.00n
MM4 net_043 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 net_043 VPW N12LL W=200.00n L=60.00n
MM5 net11 A3 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=300.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS AND3HSV0
****Sub-Circuit for AND3HSV0RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV0RD A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=200.00n L=60.00n
MM4 net9 A2 net5 VPW N12LL W=200.00n L=60.00n
MM5 net25 A1 net9 VPW N12LL W=200.00n L=60.00n
MM9 net25 A2 VDD VNW P12LL W=200.00n L=60.00n
MM8 net25 A1 VDD VNW P12LL W=200.00n L=60.00n
MM7 net25 A3 VDD VNW P12LL W=200.00n L=60.00n
MM0 Z net25 VSS VPW N12LL W=200.00n L=60n
MM1 Z net25 VDD VNW P12LL W=250.00n L=60n
.ENDS AND3HSV0RD
****Sub-Circuit for AND3HSV1, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND3HSV1 A1 A2 A3 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=200.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=290.00n L=60.00n
MM4 net_043 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 net_043 VPW N12LL W=200.00n L=60.00n
MM5 net11 A3 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=440.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS AND3HSV1
****Sub-Circuit for AND3HSV12, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV12 A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=1.29u L=60.00n
MM4 net9 A2 net5 VPW N12LL W=1.29u L=60.00n
MM5 net25 A1 net9 VPW N12LL W=1.29u L=60.00n
MM9 net25 A2 VDD VNW P12LL W=1.32u L=60.00n
MM8 net25 A1 VDD VNW P12LL W=1.32u L=60.00n
MM7 net25 A3 VDD VNW P12LL W=1.32u L=60.00n
MM0 Z net25 VSS VPW N12LL W=2.58u L=60n
MM1 Z net25 VDD VNW P12LL W=3.24u L=60n
.ENDS AND3HSV12
****Sub-Circuit for AND3HSV12RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV12RD A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=2.58u L=60.00n
MM4 net9 A2 net5 VPW N12LL W=2.58u L=60.00n
MM5 net25 A1 net9 VPW N12LL W=2.58u L=60.00n
MM9 net25 A2 VDD VNW P12LL W=2.1u L=60.00n
MM8 net25 A1 VDD VNW P12LL W=2.1u L=60.00n
MM7 net25 A3 VDD VNW P12LL W=2.1u L=60.00n
MM0 Z net25 VSS VPW N12LL W=2.58u L=60n
MM1 Z net25 VDD VNW P12LL W=3.24u L=60n
.ENDS AND3HSV12RD
****Sub-Circuit for AND3HSV12RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV12RQ A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=650.00n L=60.00n
MM4 net9 A2 net5 VPW N12LL W=650.00n L=60.00n
MM5 net25 A1 net9 VPW N12LL W=650.00n L=60.00n
MM9 net25 A2 VDD VNW P12LL W=810.00n L=60.00n
MM8 net25 A1 VDD VNW P12LL W=810.00n L=60.00n
MM7 net25 A3 VDD VNW P12LL W=810.00n L=60.00n
MM0 Z net25 VSS VPW N12LL W=2.58u L=60n
MM1 Z net25 VDD VNW P12LL W=3.24u L=60n
.ENDS AND3HSV12RQ
****Sub-Circuit for AND3HSV16, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV16 A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=1.72u L=60.00n
MM4 net9 A2 net5 VPW N12LL W=1.72u L=60.00n
MM5 net25 A1 net9 VPW N12LL W=1.72u L=60.00n
MM9 net25 A2 VDD VNW P12LL W=1.76u L=60.00n
MM8 net25 A1 VDD VNW P12LL W=1.76u L=60.00n
MM7 net25 A3 VDD VNW P12LL W=1.76u L=60.00n
MM0 Z net25 VSS VPW N12LL W=3.44u L=60n
MM1 Z net25 VDD VNW P12LL W=4.32u L=60n
.ENDS AND3HSV16
****Sub-Circuit for AND3HSV16RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV16RD A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=3.44u L=60.00n
MM4 net9 A2 net5 VPW N12LL W=3.44u L=60.00n
MM5 net25 A1 net9 VPW N12LL W=3.44u L=60.00n
MM9 net25 A2 VDD VNW P12LL W=2.8u L=60.00n
MM8 net25 A1 VDD VNW P12LL W=2.8u L=60.00n
MM7 net25 A3 VDD VNW P12LL W=2.8u L=60.00n
MM0 Z net25 VSS VPW N12LL W=3.44u L=60n
MM1 Z net25 VDD VNW P12LL W=4.32u L=60n
.ENDS AND3HSV16RD
****Sub-Circuit for AND3HSV16RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV16RQ A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=860.00n L=60.00n
MM4 net9 A2 net5 VPW N12LL W=860.00n L=60.00n
MM5 net25 A1 net9 VPW N12LL W=860.00n L=60.00n
MM9 net25 A2 VDD VNW P12LL W=1.08u L=60.00n
MM8 net25 A1 VDD VNW P12LL W=1.08u L=60.00n
MM7 net25 A3 VDD VNW P12LL W=1.08u L=60.00n
MM0 Z net25 VSS VPW N12LL W=3.44u L=60n
MM1 Z net25 VDD VNW P12LL W=4.32u L=60n
.ENDS AND3HSV16RQ
****Sub-Circuit for AND3HSV1RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV1RD A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=410.00n L=60.00n
MM4 net9 A2 net5 VPW N12LL W=410.00n L=60.00n
MM5 net25 A1 net9 VPW N12LL W=410.00n L=60.00n
MM9 net25 A2 VDD VNW P12LL W=280.00n L=60.00n
MM8 net25 A1 VDD VNW P12LL W=280.00n L=60.00n
MM7 net25 A3 VDD VNW P12LL W=280.00n L=60.00n
MM0 Z net25 VSS VPW N12LL W=350.00n L=60n
MM1 Z net25 VDD VNW P12LL W=440.00n L=60n
.ENDS AND3HSV1RD
****Sub-Circuit for AND3HSV2, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND3HSV2 A1 A2 A3 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=200.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=430.00n L=60.00n
MM4 net_043 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 net_043 VPW N12LL W=200.00n L=60.00n
MM5 net11 A3 VDD VNW P12LL W=300.0n L=60.00n
MM3 Z net11 VDD VNW P12LL W=650.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.0n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.0n L=60.00n
.ENDS AND3HSV2
****Sub-Circuit for AND3HSV2RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV2RD A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=430.00n L=60.00n
MM4 net9 A2 net5 VPW N12LL W=430.00n L=60.00n
MM5 net25 A1 net9 VPW N12LL W=430.00n L=60.00n
MM9 net25 A2 VDD VNW P12LL W=350.00n L=60.00n
MM8 net25 A1 VDD VNW P12LL W=350.00n L=60.00n
MM7 net25 A3 VDD VNW P12LL W=350.00n L=60.00n
MM0 Z net25 VSS VPW N12LL W=430.00n L=60n
MM1 Z net25 VDD VNW P12LL W=540.00n L=60n
.ENDS AND3HSV2RD
****Sub-Circuit for AND3HSV4, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND3HSV4 A1 A2 A3 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=350.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=860.00n L=60.00n
MM4 net_043 A3 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net18 A2 net_043 VPW N12LL W=350.00n L=60.00n
MM5 net11 A3 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=1.3u L=60.00n
MM0 net11 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=520.00n L=60.00n
.ENDS AND3HSV4
****Sub-Circuit for AND3HSV4RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV4RD A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=860.00n L=60.00n
MM4 net9 A2 net5 VPW N12LL W=860.00n L=60.00n
MM5 net25 A1 net9 VPW N12LL W=860.00n L=60.00n
MM9 net25 A2 VDD VNW P12LL W=700.00n L=60.00n
MM8 net25 A1 VDD VNW P12LL W=700.00n L=60.00n
MM7 net25 A3 VDD VNW P12LL W=700.00n L=60.00n
MM0 Z net25 VSS VPW N12LL W=860.00n L=60n
MM1 Z net25 VDD VNW P12LL W=1.08u L=60n
.ENDS AND3HSV4RD
****Sub-Circuit for AND3HSV4RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV4RQ A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=270.00n L=60.00n
MM4 net9 A2 net5 VPW N12LL W=270.00n L=60.00n
MM5 net25 A1 net9 VPW N12LL W=270.00n L=60.00n
MM9 net25 A2 VDD VNW P12LL W=270.00n L=60.00n
MM8 net25 A1 VDD VNW P12LL W=270.00n L=60.00n
MM7 net25 A3 VDD VNW P12LL W=270.00n L=60.00n
MM0 Z net25 VSS VPW N12LL W=860.00n L=60n
MM1 Z net25 VDD VNW P12LL W=1.08u L=60n
.ENDS AND3HSV4RQ
****Sub-Circuit for AND3HSV8, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND3HSV8 A1 A2 A3 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=700.0n L=60.00n
MM2 Z net11 VSS VPW N12LL W=1.72u L=60.00n
MM4 net_043 A3 VSS VPW N12LL W=700.0n L=60.00n
MMN1 net18 A2 net_043 VPW N12LL W=700.0n L=60.00n
MM5 net11 A3 VDD VNW P12LL W=1.04u L=60.00n
MM3 Z net11 VDD VNW P12LL W=2.6u L=60.00n
MM0 net11 A2 VDD VNW P12LL W=1.04u L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=1.04u L=60.00n
.ENDS AND3HSV8
****Sub-Circuit for AND3HSV8RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV8RD A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=1.72u L=60.00n
MM4 net9 A2 net5 VPW N12LL W=1.72u L=60.00n
MM5 net25 A1 net9 VPW N12LL W=1.72u L=60.00n
MM9 net25 A2 VDD VNW P12LL W=1.4u L=60.00n
MM8 net25 A1 VDD VNW P12LL W=1.4u L=60.00n
MM7 net25 A3 VDD VNW P12LL W=1.4u L=60.00n
MM0 Z net25 VSS VPW N12LL W=1.72u L=60n
MM1 Z net25 VDD VNW P12LL W=2.16u L=60n
.ENDS AND3HSV8RD
****Sub-Circuit for AND3HSV8RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND3HSV8RQ A1 A2 A3 Z VDD VSS
MM6 net5 A3 VSS VPW N12LL W=430.00n L=60.00n
MM4 net9 A2 net5 VPW N12LL W=430.00n L=60.00n
MM5 net25 A1 net9 VPW N12LL W=430.00n L=60.00n
MM9 net25 A2 VDD VNW P12LL W=540.00n L=60.00n
MM8 net25 A1 VDD VNW P12LL W=540.00n L=60.00n
MM7 net25 A3 VDD VNW P12LL W=540.00n L=60.00n
MM0 Z net25 VSS VPW N12LL W=1.72u L=60n
MM1 Z net25 VDD VNW P12LL W=2.16u L=60n
.ENDS AND3HSV8RQ
****Sub-Circuit for AND4HSV0, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND4HSV0 A1 A2 A3 A4 Z VDD VSS
MM6 net_042 A4 VSS VPW N12LL W=200.00n L=60.00n
MM1 net11 A1 net18 VPW N12LL W=200.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=200.00n L=60.00n
MM4 net_054 A3 net_042 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 net_054 VPW N12LL W=200.00n L=60.00n
MM7 net11 A4 VDD VNW P12LL W=300.00n L=60.00n
MM5 net11 A3 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=300.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS AND4HSV0
****Sub-Circuit for AND4HSV0RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV0RD A1 A2 A3 A4 Z VDD VSS
MM1 Z net26 VDD VNW P12LL W=250.00n L=60n
MM0 Z net26 VSS VPW N12LL W=200.00n L=60n
MM7 net26 A3 VDD VNW P12LL W=200.00n L=60.00n
MM8 net26 A1 VDD VNW P12LL W=200.00n L=60.00n
MM9 net26 A2 VDD VNW P12LL W=200.00n L=60.00n
MM3 net26 A4 VDD VNW P12LL W=200.00n L=60.00n
MM5 net26 A1 net34 VPW N12LL W=200.00n L=60.00n
MM4 net34 A2 net38 VPW N12LL W=200.00n L=60.00n
MM6 net38 A3 net42 VPW N12LL W=200.00n L=60.00n
MM2 net42 A4 VSS VPW N12LL W=200.00n L=60.00n
.ENDS AND4HSV0RD
****Sub-Circuit for AND4HSV1, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND4HSV1 A1 A2 A3 A4 Z VDD VSS
MM6 net_042 A4 VSS VPW N12LL W=200.00n L=60.00n
MM1 net11 A1 net18 VPW N12LL W=200.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=290.00n L=60.00n
MM4 net_054 A3 net_042 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 net_054 VPW N12LL W=200.00n L=60.00n
MM7 net11 A4 VDD VNW P12LL W=300.00n L=60.00n
MM5 net11 A3 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=440.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS AND4HSV1
****Sub-Circuit for AND4HSV12, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV12 A1 A2 A3 A4 Z VDD VSS
MMP1 net59 net44 VDD VNW P12LL W=3.9u L=60.00n
MM9 Z net52 net59 VNW P12LL W=3.9u L=60.00n
MM5 net52 A2 VDD VNW P12LL W=1.56u L=60.00n
MM4 net52 A1 VDD VNW P12LL W=1.56u L=60.00n
MM3 net44 A4 VDD VNW P12LL W=1.56u L=60.00n
MM0 net44 A3 VDD VNW P12LL W=1.56u L=60.00n
MMN1 Z net52 VSS VPW N12LL W=2.1u L=60.00n
MM8 Z net44 VSS VPW N12LL W=2.1u L=60.00n
MM7 net76 A2 VSS VPW N12LL W=1.8u L=60.00n
MM6 net52 A1 net76 VPW N12LL W=1.8u L=60.00n
MM1 net68 A4 VSS VPW N12LL W=1.8u L=60.00n
MM2 net44 A3 net68 VPW N12LL W=1.8u L=60.00n
.ENDS AND4HSV12
****Sub-Circuit for AND4HSV12RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV12RD A1 A2 A3 A4 Z VDD VSS
MMP1 net59 net44 VDD VNW P12LL W=3.9u L=60.00n
MM9 Z net52 net59 VNW P12LL W=3.9u L=60.00n
MM5 net52 A2 VDD VNW P12LL W=2.52u L=60.00n
MM4 net52 A1 VDD VNW P12LL W=2.52u L=60.00n
MM3 net44 A4 VDD VNW P12LL W=2.52u L=60.00n
MM0 net44 A3 VDD VNW P12LL W=2.52u L=60.00n
MMN1 Z net52 VSS VPW N12LL W=2.1u L=60.00n
MM8 Z net44 VSS VPW N12LL W=2.1u L=60.00n
MM7 net76 A2 VSS VPW N12LL W=2.58u L=60.00n
MM6 net52 A1 net76 VPW N12LL W=2.58u L=60.00n
MM1 net68 A4 VSS VPW N12LL W=2.58u L=60.00n
MM2 net44 A3 net68 VPW N12LL W=2.58u L=60.00n
.ENDS AND4HSV12RD
****Sub-Circuit for AND4HSV12RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV12RQ A1 A2 A3 A4 Z VDD VSS
MMP1 net59 net44 VDD VNW P12LL W=3.9u L=60.00n
MM9 Z net52 net59 VNW P12LL W=3.9u L=60.00n
MM5 net52 A2 VDD VNW P12LL W=970.00n L=60.00n
MM4 net52 A1 VDD VNW P12LL W=970.00n L=60.00n
MM3 net44 A4 VDD VNW P12LL W=970.00n L=60.00n
MM0 net44 A3 VDD VNW P12LL W=970.00n L=60.00n
MMN1 Z net52 VSS VPW N12LL W=2.1u L=60.00n
MM8 Z net44 VSS VPW N12LL W=2.1u L=60.00n
MM7 net76 A2 VSS VPW N12LL W=860.00n L=60.00n
MM6 net52 A1 net76 VPW N12LL W=860.00n L=60.00n
MM1 net68 A4 VSS VPW N12LL W=860.00n L=60.00n
MM2 net44 A3 net68 VPW N12LL W=860.00n L=60.00n
.ENDS AND4HSV12RQ
****Sub-Circuit for AND4HSV16, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV16 A1 A2 A3 A4 Z VDD VSS
MMP1 net59 net44 VDD VNW P12LL W=5.2u L=60.00n
MM9 Z net52 net59 VNW P12LL W=5.2u L=60.00n
MM5 net52 A2 VDD VNW P12LL W=2.08u L=60.00n
MM4 net52 A1 VDD VNW P12LL W=2.08u L=60.00n
MM3 net44 A4 VDD VNW P12LL W=2.08u L=60.00n
MM0 net44 A3 VDD VNW P12LL W=2.08u L=60.00n
MMN1 Z net52 VSS VPW N12LL W=2.8u L=60.00n
MM8 Z net44 VSS VPW N12LL W=2.8u L=60.00n
MM7 net76 A2 VSS VPW N12LL W=2.4u L=60.00n
MM6 net52 A1 net76 VPW N12LL W=2.4u L=60.00n
MM1 net68 A4 VSS VPW N12LL W=2.4u L=60.00n
MM2 net44 A3 net68 VPW N12LL W=2.4u L=60.00n
.ENDS AND4HSV16
****Sub-Circuit for AND4HSV16RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV16RD A1 A2 A3 A4 Z VDD VSS
MMP1 net59 net44 VDD VNW P12LL W=5.2u L=60.00n
MM9 Z net52 net59 VNW P12LL W=5.2u L=60.00n
MM5 net52 A2 VDD VNW P12LL W=3.36u L=60.00n
MM4 net52 A1 VDD VNW P12LL W=3.36u L=60.00n
MM3 net44 A4 VDD VNW P12LL W=3.36u L=60.00n
MM0 net44 A3 VDD VNW P12LL W=3.36u L=60.00n
MMN1 Z net52 VSS VPW N12LL W=2.8u L=60.00n
MM8 Z net44 VSS VPW N12LL W=2.8u L=60.00n
MM7 net76 A2 VSS VPW N12LL W=3.44u L=60.00n
MM6 net52 A1 net76 VPW N12LL W=3.44u L=60.00n
MM1 net68 A4 VSS VPW N12LL W=3.44u L=60.00n
MM2 net44 A3 net68 VPW N12LL W=3.44u L=60.00n
.ENDS AND4HSV16RD
****Sub-Circuit for AND4HSV16RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV16RQ A1 A2 A3 A4 Z VDD VSS
MMP1 net59 net44 VDD VNW P12LL W=5.2u L=60.00n
MM9 Z net52 net59 VNW P12LL W=5.2u L=60.00n
MM5 net52 A2 VDD VNW P12LL W=1.3u L=60.00n
MM4 net52 A1 VDD VNW P12LL W=1.3u L=60.00n
MM3 net44 A4 VDD VNW P12LL W=1.3u L=60.00n
MM0 net44 A3 VDD VNW P12LL W=1.3u L=60.00n
MMN1 Z net52 VSS VPW N12LL W=2.8u L=60.00n
MM8 Z net44 VSS VPW N12LL W=2.8u L=60.00n
MM7 net76 A2 VSS VPW N12LL W=860.00n L=60.00n
MM6 net52 A1 net76 VPW N12LL W=860.00n L=60.00n
MM1 net68 A4 VSS VPW N12LL W=860.00n L=60.00n
MM2 net44 A3 net68 VPW N12LL W=860.00n L=60.00n
.ENDS AND4HSV16RQ
****Sub-Circuit for AND4HSV1RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV1RD A1 A2 A3 A4 Z VDD VSS
MM1 Z net26 VDD VNW P12LL W=440.00n L=60n
MM0 Z net26 VSS VPW N12LL W=350.00n L=60n
MM7 net26 A3 VDD VNW P12LL W=280.00n L=60.00n
MM8 net26 A1 VDD VNW P12LL W=280.00n L=60.00n
MM9 net26 A2 VDD VNW P12LL W=280.00n L=60.00n
MM3 net26 A4 VDD VNW P12LL W=280.00n L=60.00n
MM5 net26 A1 net34 VPW N12LL W=410.00n L=60.00n
MM4 net34 A2 net38 VPW N12LL W=410.00n L=60.00n
MM6 net38 A3 net42 VPW N12LL W=410.00n L=60.00n
MM2 net42 A4 VSS VPW N12LL W=410.00n L=60.00n
.ENDS AND4HSV1RD
****Sub-Circuit for AND4HSV2, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND4HSV2 A1 A2 A3 A4 Z VDD VSS
MM6 net_042 A4 VSS VPW N12LL W=200.00n L=60.00n
MM1 net11 A1 net18 VPW N12LL W=200.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=430.00n L=60.00n
MM4 net_054 A3 net_042 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 net_054 VPW N12LL W=200.00n L=60.00n
MM7 net11 A4 VDD VNW P12LL W=300.00n L=60.00n
MM5 net11 A3 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=650.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS AND4HSV2
****Sub-Circuit for AND4HSV2RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV2RD A1 A2 A3 A4 Z VDD VSS
MM1 Z net26 VDD VNW P12LL W=540.00n L=60n
MM0 Z net26 VSS VPW N12LL W=430.00n L=60n
MM7 net26 A3 VDD VNW P12LL W=350.00n L=60.00n
MM8 net26 A1 VDD VNW P12LL W=350.00n L=60.00n
MM9 net26 A2 VDD VNW P12LL W=350.00n L=60.00n
MM3 net26 A4 VDD VNW P12LL W=350.00n L=60.00n
MM5 net26 A1 net34 VPW N12LL W=430.00n L=60.00n
MM4 net34 A2 net38 VPW N12LL W=430.00n L=60.00n
MM6 net38 A3 net42 VPW N12LL W=430.00n L=60.00n
MM2 net42 A4 VSS VPW N12LL W=430.00n L=60.00n
.ENDS AND4HSV2RD
****Sub-Circuit for AND4HSV4, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND4HSV4 A1 A2 A3 A4 Z VDD VSS
MM6 net_042 A4 VSS VPW N12LL W=350.00n L=60.00n
MM1 net11 A1 net18 VPW N12LL W=350.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=860.00n L=60.00n
MM4 net_054 A3 net_042 VPW N12LL W=350.00n L=60.00n
MMN1 net18 A2 net_054 VPW N12LL W=350.00n L=60.00n
MM7 net11 A4 VDD VNW P12LL W=520.00n L=60.00n
MM5 net11 A3 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=1.3u L=60.00n
MM0 net11 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=520.00n L=60.00n
.ENDS AND4HSV4
****Sub-Circuit for AND4HSV4RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV4RD A1 A2 A3 A4 Z VDD VSS
MM1 Z net26 VDD VNW P12LL W=1.08u L=60n
MM0 Z net26 VSS VPW N12LL W=860.00n L=60n
MM7 net26 A3 VDD VNW P12LL W=700.00n L=60.00n
MM8 net26 A1 VDD VNW P12LL W=700.00n L=60.00n
MM9 net26 A2 VDD VNW P12LL W=700.00n L=60.00n
MM3 net26 A4 VDD VNW P12LL W=700.00n L=60.00n
MM5 net26 A1 net34 VPW N12LL W=860.00n L=60.00n
MM4 net34 A2 net38 VPW N12LL W=860.00n L=60.00n
MM6 net38 A3 net42 VPW N12LL W=860.00n L=60.00n
MM2 net42 A4 VSS VPW N12LL W=860.00n L=60.00n
.ENDS AND4HSV4RD
****Sub-Circuit for AND4HSV4RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV4RQ A1 A2 A3 A4 Z VDD VSS
MM1 Z net26 VDD VNW P12LL W=1.08u L=60n
MM0 Z net26 VSS VPW N12LL W=860.00n L=60n
MM7 net26 A3 VDD VNW P12LL W=270.00n L=60.00n
MM8 net26 A1 VDD VNW P12LL W=270.00n L=60.00n
MM9 net26 A2 VDD VNW P12LL W=270.00n L=60.00n
MM3 net26 A4 VDD VNW P12LL W=270.00n L=60.00n
MM5 net26 A1 net34 VPW N12LL W=430.00n L=60.00n
MM4 net34 A2 net38 VPW N12LL W=430.00n L=60.00n
MM6 net38 A3 net42 VPW N12LL W=430.00n L=60.00n
MM2 net42 A4 VSS VPW N12LL W=430.00n L=60.00n
.ENDS AND4HSV4RQ
****Sub-Circuit for AND4HSV8, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AND4HSV8 A1 A2 A3 A4 Z VDD VSS
MM6 net_042 A4 VSS VPW N12LL W=705.0n L=60.00n
MM1 net11 A1 net18 VPW N12LL W=705.0n L=60.00n
MM2 Z net11 VSS VPW N12LL W=1.72u L=60.00n
MM4 net_054 A3 net_042 VPW N12LL W=705.0n L=60.00n
MMN1 net18 A2 net_054 VPW N12LL W=705.0n L=60.00n
MM7 net11 A4 VDD VNW P12LL W=1.04u L=60.00n
MM5 net11 A3 VDD VNW P12LL W=1.04u L=60.00n
MM3 Z net11 VDD VNW P12LL W=2.6u L=60.00n
MM0 net11 A2 VDD VNW P12LL W=1.04u L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=1.04u L=60.00n
.ENDS AND4HSV8
****Sub-Circuit for AND4HSV8RD, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV8RD A1 A2 A3 A4 Z VDD VSS
MMP1 net59 net44 VDD VNW P12LL W=2.6u L=60.00n
MM9 Z net52 net59 VNW P12LL W=2.6u L=60.00n
MM5 net52 A2 VDD VNW P12LL W=1.68u L=60.00n
MM4 net52 A1 VDD VNW P12LL W=1.68u L=60.00n
MM3 net44 A4 VDD VNW P12LL W=1.68u L=60.00n
MM0 net44 A3 VDD VNW P12LL W=1.68u L=60.00n
MMN1 Z net52 VSS VPW N12LL W=1.4u L=60.00n
MM8 Z net44 VSS VPW N12LL W=1.4u L=60.00n
MM7 net76 A2 VSS VPW N12LL W=1.72u L=60.00n
MM6 net52 A1 net76 VPW N12LL W=1.72u L=60.00n
MM1 net68 A4 VSS VPW N12LL W=1.72u L=60.00n
MM2 net44 A3 net68 VPW N12LL W=1.72u L=60.00n
.ENDS AND4HSV8RD
****Sub-Circuit for AND4HSV8RQ, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND4HSV8RQ A1 A2 A3 A4 Z VDD VSS
MMP1 net59 net44 VDD VNW P12LL W=2.6u L=60.00n
MM9 Z net52 net59 VNW P12LL W=2.6u L=60.00n
MM5 net52 A2 VDD VNW P12LL W=650.00n L=60.00n
MM4 net52 A1 VDD VNW P12LL W=650.00n L=60.00n
MM3 net44 A4 VDD VNW P12LL W=650.00n L=60.00n
MM0 net44 A3 VDD VNW P12LL W=650.00n L=60.00n
MMN1 Z net52 VSS VPW N12LL W=1.4u L=60.00n
MM8 Z net44 VSS VPW N12LL W=1.4u L=60.00n
MM7 net76 A2 VSS VPW N12LL W=430.00n L=60.00n
MM6 net52 A1 net76 VPW N12LL W=430.00n L=60.00n
MM1 net68 A4 VSS VPW N12LL W=430.00n L=60.00n
MM2 net44 A3 net68 VPW N12LL W=430.00n L=60.00n
.ENDS AND4HSV8RQ
****Sub-Circuit for AND5HSV0, Thu May 19 13:57:40 CST 2011****
.SUBCKT AND5HSV0 A1 A2 A3 A4 A5 Z VDD VSS
MM11 Z net49 VSS VPW N12LL W=220.00n L=60.00n
MM10 Z net53 VSS VPW N12LL W=220.00n L=60.00n
MM6 net13 A5 VSS VPW N12LL W=250.00n L=60.00n
MM4 net17 A4 net13 VPW N12LL W=250.00n L=60.00n
MM5 net49 A3 net17 VPW N12LL W=250.00n L=60.00n
MM1 net25 A2 VSS VPW N12LL W=190.00n L=60.00n
MM2 net53 A1 net25 VPW N12LL W=190.00n L=60.00n
MM13 Z net53 net36 VNW P12LL W=280.00n L=60.00n
MM12 net36 net49 VDD VNW P12LL W=280.00n L=60.00n
MM9 net49 A4 VDD VNW P12LL W=180.00n L=60.00n
MM8 net49 A3 VDD VNW P12LL W=180.00n L=60.00n
MM7 net49 A5 VDD VNW P12LL W=180.00n L=60.00n
MM3 net53 A2 VDD VNW P12LL W=180.00n L=60.00n
MM0 net53 A1 VDD VNW P12LL W=180.00n L=60.00n
.ENDS AND5HSV0
****Sub-Circuit for AND5HSV0RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV0RD A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=180.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=180.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=180.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=180.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=180.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=280.00n L=60.00n
MM13 Z net11 net34 VNW P12LL W=280.00n L=60.00n
MM2 net11 A1 net39 VPW N12LL W=210.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=210.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=260.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=260.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=260.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=220.00n L=60.00n
MM11 Z net15 VSS VPW N12LL W=220.00n L=60.00n
.ENDS AND5HSV0RD
****Sub-Circuit for AND5HSV1, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND5HSV1 A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=210.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=210.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=210.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=210.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=210.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=520.00n L=60.00n
MM13 Z net11 net34 VNW P12LL W=520.00n L=60.00n
MM2 net11 A1 net39 VPW N12LL W=240.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=240.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=300.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=300.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=300.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=280.00n L=60.00n
MM11 Z net15 VSS VPW N12LL W=280.00n L=60.00n
.ENDS AND5HSV1
****Sub-Circuit for AND5HSV12, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV12 A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=1.56u L=60.00n
MM3 net11 A2 VDD VNW P12LL W=1.56u L=60.00n
MM7 net15 A5 VDD VNW P12LL W=1.56u L=60.00n
MM8 net15 A3 VDD VNW P12LL W=1.56u L=60.00n
MM9 net15 A4 VDD VNW P12LL W=1.56u L=60.00n
MM12 net34 net15 VDD VNW P12LL W=3.9u L=60.00n
MM13 Z net11 net34 VNW P12LL W=3.9u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=1.8u L=60.00n
MM1 net39 A2 VSS VPW N12LL W=1.8u L=60.00n
MM5 net15 A3 net47 VPW N12LL W=2.28u L=60.00n
MM4 net47 A4 net51 VPW N12LL W=2.28u L=60.00n
MM6 net51 A5 VSS VPW N12LL W=2.28u L=60.00n
MM10 Z net11 VSS VPW N12LL W=2.1u L=60.00n
MM11 Z net15 VSS VPW N12LL W=2.1u L=60.00n
.ENDS AND5HSV12
****Sub-Circuit for AND5HSV12RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV12RD A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=2.52u L=60.00n
MM3 net11 A2 VDD VNW P12LL W=2.52u L=60.00n
MM7 net15 A5 VDD VNW P12LL W=2.52u L=60.00n
MM8 net15 A3 VDD VNW P12LL W=2.52u L=60.00n
MM9 net15 A4 VDD VNW P12LL W=2.52u L=60.00n
MM12 net34 net15 VDD VNW P12LL W=3.9u L=60.00n
MM13 Z net11 net34 VNW P12LL W=3.9u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=2.58u L=60.00n
MM1 net39 A2 VSS VPW N12LL W=2.58u L=60.00n
MM5 net15 A3 net47 VPW N12LL W=2.58u L=60.00n
MM4 net47 A4 net51 VPW N12LL W=2.58u L=60.00n
MM6 net51 A5 VSS VPW N12LL W=2.58u L=60.00n
MM10 Z net11 VSS VPW N12LL W=2.1u L=60.00n
MM11 Z net15 VSS VPW N12LL W=2.1u L=60.00n
.ENDS AND5HSV12RD
****Sub-Circuit for AND5HSV12RQ, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV12RQ A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=970.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=970.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=970.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=970.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=970.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=3.9u L=60.00n
MM13 Z net11 net34 VNW P12LL W=3.9u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=860.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=860.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=860.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=860.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=860.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=2.1u L=60.00n
MM11 Z net15 VSS VPW N12LL W=2.1u L=60.00n
.ENDS AND5HSV12RQ
****Sub-Circuit for AND5HSV16, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV16 A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=2.08u L=60.00n
MM3 net11 A2 VDD VNW P12LL W=2.08u L=60.00n
MM7 net15 A5 VDD VNW P12LL W=2.08u L=60.00n
MM8 net15 A3 VDD VNW P12LL W=2.08u L=60.00n
MM9 net15 A4 VDD VNW P12LL W=2.08u L=60.00n
MM12 net34 net15 VDD VNW P12LL W=5.2u L=60.00n
MM13 Z net11 net34 VNW P12LL W=5.2u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=2.4u L=60.00n
MM1 net39 A2 VSS VPW N12LL W=2.4u L=60.00n
MM5 net15 A3 net47 VPW N12LL W=3.04u L=60.00n
MM4 net47 A4 net51 VPW N12LL W=3.04u L=60.00n
MM6 net51 A5 VSS VPW N12LL W=3.04u L=60.00n
MM10 Z net11 VSS VPW N12LL W=2.8u L=60.00n
MM11 Z net15 VSS VPW N12LL W=2.8u L=60.00n
.ENDS AND5HSV16
****Sub-Circuit for AND5HSV16RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV16RD A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=3.36u L=60.00n
MM3 net11 A2 VDD VNW P12LL W=3.36u L=60.00n
MM7 net15 A5 VDD VNW P12LL W=3.36u L=60.00n
MM8 net15 A3 VDD VNW P12LL W=3.36u L=60.00n
MM9 net15 A4 VDD VNW P12LL W=3.36u L=60.00n
MM12 net34 net15 VDD VNW P12LL W=5.2u L=60.00n
MM13 Z net11 net34 VNW P12LL W=5.2u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=3.44u L=60.00n
MM1 net39 A2 VSS VPW N12LL W=3.44u L=60.00n
MM5 net15 A3 net47 VPW N12LL W=3.44u L=60.00n
MM4 net47 A4 net51 VPW N12LL W=3.44u L=60.00n
MM6 net51 A5 VSS VPW N12LL W=3.44u L=60.00n
MM10 Z net11 VSS VPW N12LL W=2.8u L=60.00n
MM11 Z net15 VSS VPW N12LL W=2.8u L=60.00n
.ENDS AND5HSV16RD
****Sub-Circuit for AND5HSV16RQ, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV16RQ A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=1.3u L=60.00n
MM3 net11 A2 VDD VNW P12LL W=1.3u L=60.00n
MM7 net15 A5 VDD VNW P12LL W=1.3u L=60.00n
MM8 net15 A3 VDD VNW P12LL W=1.3u L=60.00n
MM9 net15 A4 VDD VNW P12LL W=1.3u L=60.00n
MM12 net34 net15 VDD VNW P12LL W=5.2u L=60.00n
MM13 Z net11 net34 VNW P12LL W=5.2u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=860.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=860.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=860.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=860.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=860.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=2.8u L=60.00n
MM11 Z net15 VSS VPW N12LL W=2.8u L=60.00n
.ENDS AND5HSV16RQ
****Sub-Circuit for AND5HSV1RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV1RD A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=340.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=340.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=340.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=340.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=340.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=520.00n L=60.00n
MM13 Z net11 net34 VNW P12LL W=520.00n L=60.00n
MM2 net11 A1 net39 VPW N12LL W=390.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=390.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=430.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=430.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=430.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=280.00n L=60.00n
MM11 Z net15 VSS VPW N12LL W=280.00n L=60.00n
.ENDS AND5HSV1RD
****Sub-Circuit for AND5HSV2, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND5HSV2 A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=260.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=260.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=260.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=260.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=260.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=650.00n L=60.00n
MM13 Z net11 net34 VNW P12LL W=650.00n L=60.00n
MM2 net11 A1 net39 VPW N12LL W=300.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=300.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=380.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=380.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=380.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=350.00n L=60.00n
MM11 Z net15 VSS VPW N12LL W=350.00n L=60.00n
.ENDS AND5HSV2
****Sub-Circuit for AND5HSV2RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV2RD A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=420.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=420.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=420.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=420.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=420.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=650.00n L=60.00n
MM13 Z net11 net34 VNW P12LL W=650.00n L=60.00n
MM2 net11 A1 net39 VPW N12LL W=430.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=430.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=430.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=430.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=430.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=350.00n L=60.00n
MM11 Z net15 VSS VPW N12LL W=350.00n L=60.00n
.ENDS AND5HSV2RD
****Sub-Circuit for AND5HSV4, Thu Dec 16 16:16:04 CST 2010****
.SUBCKT AND5HSV4 A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=520.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=520.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=520.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=520.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=520.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=1.3u L=60.00n
MM13 Z net11 net34 VNW P12LL W=1.3u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=600.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=600.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=760.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=760.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=760.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=700.00n L=60.00n
MM11 Z net15 VSS VPW N12LL W=700.00n L=60.00n
.ENDS AND5HSV4
****Sub-Circuit for AND5HSV4RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV4RD A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=840.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=840.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=840.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=840.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=840.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=1.3u L=60.00n
MM13 Z net11 net34 VNW P12LL W=1.3u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=860.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=860.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=860.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=860.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=860.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=700.00n L=60.00n
MM11 Z net15 VSS VPW N12LL W=700.00n L=60.00n
.ENDS AND5HSV4RD
****Sub-Circuit for AND5HSV4RQ, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV4RQ A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=320.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=320.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=320.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=320.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=320.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=1.3u L=60.00n
MM13 Z net11 net34 VNW P12LL W=1.3u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=370.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=370.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=370.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=370.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=370.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=700.00n L=60.00n
MM11 Z net15 VSS VPW N12LL W=700.00n L=60.00n
.ENDS AND5HSV4RQ
****Sub-Circuit for AND5HSV8, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV8 A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=1.04u L=60.00n
MM3 net11 A2 VDD VNW P12LL W=1.04u L=60.00n
MM7 net15 A5 VDD VNW P12LL W=1.04u L=60.00n
MM8 net15 A3 VDD VNW P12LL W=1.04u L=60.00n
MM9 net15 A4 VDD VNW P12LL W=1.04u L=60.00n
MM12 net34 net15 VDD VNW P12LL W=2.6u L=60.00n
MM13 Z net11 net34 VNW P12LL W=2.6u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=1.2u L=60.00n
MM1 net39 A2 VSS VPW N12LL W=1.2u L=60.00n
MM5 net15 A3 net47 VPW N12LL W=1.52u L=60.00n
MM4 net47 A4 net51 VPW N12LL W=1.52u L=60.00n
MM6 net51 A5 VSS VPW N12LL W=1.52u L=60.00n
MM10 Z net11 VSS VPW N12LL W=1.4u L=60.00n
MM11 Z net15 VSS VPW N12LL W=1.4u L=60.00n
.ENDS AND5HSV8
****Sub-Circuit for AND5HSV8RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV8RD A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=1.68u L=60.00n
MM3 net11 A2 VDD VNW P12LL W=1.68u L=60.00n
MM7 net15 A5 VDD VNW P12LL W=1.68u L=60.00n
MM8 net15 A3 VDD VNW P12LL W=1.68u L=60.00n
MM9 net15 A4 VDD VNW P12LL W=1.68u L=60.00n
MM12 net34 net15 VDD VNW P12LL W=2.6u L=60.00n
MM13 Z net11 net34 VNW P12LL W=2.6u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=1.72u L=60.00n
MM1 net39 A2 VSS VPW N12LL W=1.72u L=60.00n
MM5 net15 A3 net47 VPW N12LL W=1.72u L=60.00n
MM4 net47 A4 net51 VPW N12LL W=1.72u L=60.00n
MM6 net51 A5 VSS VPW N12LL W=1.72u L=60.00n
MM10 Z net11 VSS VPW N12LL W=1.4u L=60.00n
MM11 Z net15 VSS VPW N12LL W=1.4u L=60.00n
.ENDS AND5HSV8RD
****Sub-Circuit for AND5HSV8RQ, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND5HSV8RQ A1 A2 A3 A4 A5 Z VDD VSS
MM0 net11 A1 VDD VNW P12LL W=650.00n L=60.00n
MM3 net11 A2 VDD VNW P12LL W=650.00n L=60.00n
MM7 net15 A5 VDD VNW P12LL W=650.00n L=60.00n
MM8 net15 A3 VDD VNW P12LL W=650.00n L=60.00n
MM9 net15 A4 VDD VNW P12LL W=650.00n L=60.00n
MM12 net34 net15 VDD VNW P12LL W=2.6u L=60.00n
MM13 Z net11 net34 VNW P12LL W=2.6u L=60.00n
MM2 net11 A1 net39 VPW N12LL W=430.00n L=60.00n
MM1 net39 A2 VSS VPW N12LL W=430.00n L=60.00n
MM5 net15 A3 net47 VPW N12LL W=430.00n L=60.00n
MM4 net47 A4 net51 VPW N12LL W=430.00n L=60.00n
MM6 net51 A5 VSS VPW N12LL W=430.00n L=60.00n
MM10 Z net11 VSS VPW N12LL W=1.4u L=60.00n
MM11 Z net15 VSS VPW N12LL W=1.4u L=60.00n
.ENDS AND5HSV8RQ
****Sub-Circuit for AND6HSV0, Thu May 19 13:57:40 CST 2011****
.SUBCKT AND6HSV0 A1 A2 A3 A4 A5 A6 Z VDD VSS
MM0 net7 A3 VDD VNW P12LL W=180.00n L=60.00n
MM1 net7 A1 VDD VNW P12LL W=180.00n L=60.00n
MM7 net19 A6 VDD VNW P12LL W=180.00n L=60.00n
MM8 net19 A4 VDD VNW P12LL W=180.00n L=60.00n
MM9 net19 A5 VDD VNW P12LL W=180.00n L=60.00n
MM12 net38 net19 VDD VNW P12LL W=280.00n L=60.00n
MM13 Z net7 net38 VNW P12LL W=280.00n L=60.00n
MM2 net7 A2 VDD VNW P12LL W=180.00n L=60.00n
MM3 net7 A1 net43 VPW N12LL W=250.00n L=60.00n
MM5 net19 A4 net55 VPW N12LL W=250.00n L=60.00n
MM4 net55 A5 net59 VPW N12LL W=250.00n L=60.00n
MM6 net59 A6 VSS VPW N12LL W=250.00n L=60.00n
MM10 Z net7 VSS VPW N12LL W=220.00n L=60.00n
MM11 Z net19 VSS VPW N12LL W=220.00n L=60.00n
MM14 net43 A2 net47 VPW N12LL W=250.00n L=60.00n
MM15 net47 A3 VSS VPW N12LL W=250.00n L=60.00n
.ENDS AND6HSV0
****Sub-Circuit for AND6HSV0RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV0RD A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=220.00n L=60.00n
MM10 Z net68 VSS VPW N12LL W=220.00n L=60.00n
MM6 net16 A6 VSS VPW N12LL W=260.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=260.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=260.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=260.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=260.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=260.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=280.00n L=60.00n
MM12 net43 net56 VDD VNW P12LL W=280.00n L=60.00n
MM9 net56 A5 VDD VNW P12LL W=180.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=180.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=180.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=180.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=180.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=180.00n L=60.00n
.ENDS AND6HSV0RD
****Sub-Circuit for AND6HSV1, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV1 A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=280.00n L=60.00n
MM10 Z net68 VSS VPW N12LL W=280.00n L=60.00n
MM6 net16 A6 VSS VPW N12LL W=300.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=300.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=300.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=300.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=300.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=300.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=520.00n L=60.00n
MM12 net43 net56 VDD VNW P12LL W=520.00n L=60.00n
MM9 net56 A5 VDD VNW P12LL W=210.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=210.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=210.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=210.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=210.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=210.00n L=60.00n
.ENDS AND6HSV1
****Sub-Circuit for AND6HSV12, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV12 A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=2.1u L=60.00n
MM10 Z net68 VSS VPW N12LL W=2.1u L=60.00n
MM6 net16 A6 VSS VPW N12LL W=2.28u L=60.00n
MM4 net20 A5 net16 VPW N12LL W=2.28u L=60.00n
MM5 net56 A4 net20 VPW N12LL W=2.28u L=60.00n
MM15 net28 A3 VSS VPW N12LL W=2.28u L=60.00n
MM14 net32 A2 net28 VPW N12LL W=2.28u L=60.00n
MM3 net68 A1 net32 VPW N12LL W=2.28u L=60.00n
MM13 Z net68 net43 VNW P12LL W=3.9u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=3.9u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=1.56u L=60.00n
MM8 net56 A4 VDD VNW P12LL W=1.56u L=60.00n
MM7 net56 A6 VDD VNW P12LL W=1.56u L=60.00n
MM2 net68 A2 VDD VNW P12LL W=1.56u L=60.00n
MM1 net68 A1 VDD VNW P12LL W=1.56u L=60.00n
MM0 net68 A3 VDD VNW P12LL W=1.56u L=60.00n
.ENDS AND6HSV12
****Sub-Circuit for AND6HSV12RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV12RD A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=2.1u L=60.00n
MM10 Z net68 VSS VPW N12LL W=2.1u L=60.00n
MM6 net16 A6 VSS VPW N12LL W=2.58u L=60.00n
MM4 net20 A5 net16 VPW N12LL W=2.58u L=60.00n
MM5 net56 A4 net20 VPW N12LL W=2.58u L=60.00n
MM15 net28 A3 VSS VPW N12LL W=2.58u L=60.00n
MM14 net32 A2 net28 VPW N12LL W=2.58u L=60.00n
MM3 net68 A1 net32 VPW N12LL W=2.58u L=60.00n
MM13 Z net68 net43 VNW P12LL W=3.9u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=3.9u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=2.52u L=60.00n
MM8 net56 A4 VDD VNW P12LL W=2.52u L=60.00n
MM7 net56 A6 VDD VNW P12LL W=2.52u L=60.00n
MM2 net68 A2 VDD VNW P12LL W=2.52u L=60.00n
MM1 net68 A1 VDD VNW P12LL W=2.52u L=60.00n
MM0 net68 A3 VDD VNW P12LL W=2.52u L=60.00n
.ENDS AND6HSV12RD
****Sub-Circuit for AND6HSV12RQ, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV12RQ A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=2.1u L=60.00n
MM10 Z net68 VSS VPW N12LL W=2.1u L=60.00n
MM6 net16 A6 VSS VPW N12LL W=860.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=860.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=860.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=860.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=860.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=860.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=3.9u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=3.9u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=860.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=860.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=860.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=860.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=860.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=860.00n L=60.00n
.ENDS AND6HSV12RQ
****Sub-Circuit for AND6HSV16, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV16 A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=2.8u L=60.00n
MM10 Z net68 VSS VPW N12LL W=2.8u L=60.00n
MM6 net16 A6 VSS VPW N12LL W=3.04u L=60.00n
MM4 net20 A5 net16 VPW N12LL W=3.04u L=60.00n
MM5 net56 A4 net20 VPW N12LL W=3.04u L=60.00n
MM15 net28 A3 VSS VPW N12LL W=3.04u L=60.00n
MM14 net32 A2 net28 VPW N12LL W=3.04u L=60.00n
MM3 net68 A1 net32 VPW N12LL W=3.04u L=60.00n
MM13 Z net68 net43 VNW P12LL W=5.2u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=5.2u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=2.08u L=60.00n
MM8 net56 A4 VDD VNW P12LL W=2.08u L=60.00n
MM7 net56 A6 VDD VNW P12LL W=2.08u L=60.00n
MM2 net68 A2 VDD VNW P12LL W=2.08u L=60.00n
MM1 net68 A1 VDD VNW P12LL W=2.08u L=60.00n
MM0 net68 A3 VDD VNW P12LL W=2.08u L=60.00n
.ENDS AND6HSV16
****Sub-Circuit for AND6HSV16RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV16RD A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=2.8u L=60.00n
MM10 Z net68 VSS VPW N12LL W=2.8u L=60.00n
MM6 net16 A6 VSS VPW N12LL W=3.44u L=60.00n
MM4 net20 A5 net16 VPW N12LL W=3.44u L=60.00n
MM5 net56 A4 net20 VPW N12LL W=3.44u L=60.00n
MM15 net28 A3 VSS VPW N12LL W=3.44u L=60.00n
MM14 net32 A2 net28 VPW N12LL W=3.44u L=60.00n
MM3 net68 A1 net32 VPW N12LL W=3.44u L=60.00n
MM13 Z net68 net43 VNW P12LL W=5.2u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=5.2u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=3.36u L=60.00n
MM8 net56 A4 VDD VNW P12LL W=3.36u L=60.00n
MM7 net56 A6 VDD VNW P12LL W=3.36u L=60.00n
MM2 net68 A2 VDD VNW P12LL W=3.36u L=60.00n
MM1 net68 A1 VDD VNW P12LL W=3.36u L=60.00n
MM0 net68 A3 VDD VNW P12LL W=3.36u L=60.00n
.ENDS AND6HSV16RD
****Sub-Circuit for AND6HSV16RQ, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV16RQ A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=2.8u L=60.00n
MM10 Z net68 VSS VPW N12LL W=2.8u L=60.00n
MM6 net16 A6 VSS VPW N12LL W=860.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=860.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=860.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=860.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=860.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=860.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=5.2u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=5.2u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=1.3u L=60.00n
MM8 net56 A4 VDD VNW P12LL W=1.3u L=60.00n
MM7 net56 A6 VDD VNW P12LL W=1.3u L=60.00n
MM2 net68 A2 VDD VNW P12LL W=1.3u L=60.00n
MM1 net68 A1 VDD VNW P12LL W=1.3u L=60.00n
MM0 net68 A3 VDD VNW P12LL W=1.3u L=60.00n
.ENDS AND6HSV16RQ
****Sub-Circuit for AND6HSV1RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV1RD A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=280.00n L=60.00n
MM10 Z net68 VSS VPW N12LL W=280.00n L=60.00n
MM6 net16 A6 VSS VPW N12LL W=430.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=430.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=430.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=430.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=430.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=430.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=520.00n L=60.00n
MM12 net43 net56 VDD VNW P12LL W=520.00n L=60.00n
MM9 net56 A5 VDD VNW P12LL W=340.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=340.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=340.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=340.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=340.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=340.00n L=60.00n
.ENDS AND6HSV1RD
****Sub-Circuit for AND6HSV2, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV2 A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=350.00n L=60.00n
MM10 Z net68 VSS VPW N12LL W=350.00n L=60.00n
MM6 net16 A6 VSS VPW N12LL W=380.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=380.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=380.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=380.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=380.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=380.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=650.00n L=60.00n
MM12 net43 net56 VDD VNW P12LL W=650.00n L=60.00n
MM9 net56 A5 VDD VNW P12LL W=260.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=260.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=260.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=260.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=260.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=260.00n L=60.00n
.ENDS AND6HSV2
****Sub-Circuit for AND6HSV2RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV2RD A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=350.00n L=60.00n
MM10 Z net68 VSS VPW N12LL W=350.00n L=60.00n
MM6 net16 A6 VSS VPW N12LL W=430.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=430.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=430.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=430.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=430.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=430.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=650.00n L=60.00n
MM12 net43 net56 VDD VNW P12LL W=650.00n L=60.00n
MM9 net56 A5 VDD VNW P12LL W=420.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=420.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=420.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=420.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=420.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=420.00n L=60.00n
.ENDS AND6HSV2RD
****Sub-Circuit for AND6HSV4, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV4 A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=700.00n L=60.00n
MM10 Z net68 VSS VPW N12LL W=700.00n L=60.00n
MM6 net16 A6 VSS VPW N12LL W=760.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=760.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=760.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=760.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=760.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=760.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=1.3u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=1.3u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=520.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=520.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=520.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=520.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=520.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=520.00n L=60.00n
.ENDS AND6HSV4
****Sub-Circuit for AND6HSV4RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV4RD A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=700.00n L=60.00n
MM10 Z net68 VSS VPW N12LL W=700.00n L=60.00n
MM6 net16 A6 VSS VPW N12LL W=860.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=860.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=860.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=860.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=860.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=860.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=1.3u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=1.3u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=840.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=840.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=840.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=840.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=840.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=840.00n L=60.00n
.ENDS AND6HSV4RD
****Sub-Circuit for AND6HSV4RQ, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV4RQ A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=700.00n L=60.00n
MM10 Z net68 VSS VPW N12LL W=700.00n L=60.00n
MM6 net16 A6 VSS VPW N12LL W=370.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=370.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=370.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=370.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=370.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=370.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=1.3u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=1.3u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=320.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=320.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=320.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=320.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=320.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=320.00n L=60.00n
.ENDS AND6HSV4RQ
****Sub-Circuit for AND6HSV8, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV8 A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=1.4u L=60.00n
MM10 Z net68 VSS VPW N12LL W=1.4u L=60.00n
MM6 net16 A6 VSS VPW N12LL W=1.52u L=60.00n
MM4 net20 A5 net16 VPW N12LL W=1.52u L=60.00n
MM5 net56 A4 net20 VPW N12LL W=1.52u L=60.00n
MM15 net28 A3 VSS VPW N12LL W=1.52u L=60.00n
MM14 net32 A2 net28 VPW N12LL W=1.52u L=60.00n
MM3 net68 A1 net32 VPW N12LL W=1.52u L=60.00n
MM13 Z net68 net43 VNW P12LL W=2.6u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=2.6u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=1.04u L=60.00n
MM8 net56 A4 VDD VNW P12LL W=1.04u L=60.00n
MM7 net56 A6 VDD VNW P12LL W=1.04u L=60.00n
MM2 net68 A2 VDD VNW P12LL W=1.04u L=60.00n
MM1 net68 A1 VDD VNW P12LL W=1.04u L=60.00n
MM0 net68 A3 VDD VNW P12LL W=1.04u L=60.00n
.ENDS AND6HSV8
****Sub-Circuit for AND6HSV8RD, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV8RD A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=1.4u L=60.00n
MM10 Z net68 VSS VPW N12LL W=1.4u L=60.00n
MM6 net16 A6 VSS VPW N12LL W=1.72u L=60.00n
MM4 net20 A5 net16 VPW N12LL W=1.72u L=60.00n
MM5 net56 A4 net20 VPW N12LL W=1.72u L=60.00n
MM15 net28 A3 VSS VPW N12LL W=1.72u L=60.00n
MM14 net32 A2 net28 VPW N12LL W=1.72u L=60.00n
MM3 net68 A1 net32 VPW N12LL W=1.72u L=60.00n
MM13 Z net68 net43 VNW P12LL W=2.6u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=2.6u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=1.68u L=60.00n
MM8 net56 A4 VDD VNW P12LL W=1.68u L=60.00n
MM7 net56 A6 VDD VNW P12LL W=1.68u L=60.00n
MM2 net68 A2 VDD VNW P12LL W=1.68u L=60.00n
MM1 net68 A1 VDD VNW P12LL W=1.68u L=60.00n
MM0 net68 A3 VDD VNW P12LL W=1.68u L=60.00n
.ENDS AND6HSV8RD
****Sub-Circuit for AND6HSV8RQ, Thu Dec 16 16:16:05 CST 2010****
.SUBCKT AND6HSV8RQ A1 A2 A3 A4 A5 A6 Z VDD VSS
MM11 Z net56 VSS VPW N12LL W=1.4u L=60.00n
MM10 Z net68 VSS VPW N12LL W=1.4u L=60.00n
MM6 net16 A6 VSS VPW N12LL W=430.00n L=60.00n
MM4 net20 A5 net16 VPW N12LL W=430.00n L=60.00n
MM5 net56 A4 net20 VPW N12LL W=430.00n L=60.00n
MM15 net28 A3 VSS VPW N12LL W=430.00n L=60.00n
MM14 net32 A2 net28 VPW N12LL W=430.00n L=60.00n
MM3 net68 A1 net32 VPW N12LL W=430.00n L=60.00n
MM13 Z net68 net43 VNW P12LL W=2.6u L=60.00n
MM12 net43 net56 VDD VNW P12LL W=2.6u L=60.00n
MM9 net56 A5 VDD VNW P12LL W=650.00n L=60.00n
MM8 net56 A4 VDD VNW P12LL W=650.00n L=60.00n
MM7 net56 A6 VDD VNW P12LL W=650.00n L=60.00n
MM2 net68 A2 VDD VNW P12LL W=650.00n L=60.00n
MM1 net68 A1 VDD VNW P12LL W=650.00n L=60.00n
MM0 net68 A3 VDD VNW P12LL W=650.00n L=60.00n
.ENDS AND6HSV8RQ
****Sub-Circuit for AO211HSV0, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO211HSV0 A1 A2 B C Z VDD VSS
MM6 net1 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net1 A1 net4 VPW N12LL W=200.00n L=60.00n
MM2 Z net1 VSS VPW N12LL W=200.00n L=60.00n
MM4 net1 C VSS VPW N12LL W=200.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=200.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net1 VDD VNW P12LL W=300.00n L=60.00n
MM0 net2 B net3 VNW P12LL W=300.00n L=60.00n
MMP1 net1 C net2 VNW P12LL W=300.00n L=60.00n
.ENDS AO211HSV0
****Sub-Circuit for AO211HSV1, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO211HSV1 A1 A2 B C Z VDD VSS
MM6 net1 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net1 A1 net4 VPW N12LL W=200.00n L=60.00n
MM2 Z net1 VSS VPW N12LL W=290.00n L=60.00n
MM4 net1 C VSS VPW N12LL W=200.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=200.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net1 VDD VNW P12LL W=440.00n L=60.00n
MM0 net2 B net3 VNW P12LL W=300.00n L=60.00n
MMP1 net1 C net2 VNW P12LL W=300.00n L=60.00n
.ENDS AO211HSV1
****Sub-Circuit for AO211HSV2, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO211HSV2 A1 A2 B C Z VDD VSS
MM6 net1 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net1 A1 net4 VPW N12LL W=200.00n L=60.00n
MM2 Z net1 VSS VPW N12LL W=390.00n L=60.00n
MM4 net1 C VSS VPW N12LL W=200.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=200.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net1 VDD VNW P12LL W=650.00n L=60.00n
MM0 net2 B net3 VNW P12LL W=300.00n L=60.00n
MMP1 net1 C net2 VNW P12LL W=300.00n L=60.00n
.ENDS AO211HSV2
****Sub-Circuit for AO211HSV4, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO211HSV4 A1 A2 B C Z VDD VSS
MM6 net1 B VSS VPW N12LL W=350.00n L=60.00n
MM1 net1 A1 net4 VPW N12LL W=350.00n L=60.00n
MM2 Z net1 VSS VPW N12LL W=860.00n L=60.00n
MM4 net1 C VSS VPW N12LL W=350.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=350.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=520.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z net1 VDD VNW P12LL W=1.3u L=60.00n
MM0 net2 B net3 VNW P12LL W=520.00n L=60.00n
MMP1 net1 C net2 VNW P12LL W=520.00n L=60.00n
.ENDS AO211HSV4
****Sub-Circuit for AO21HSV0, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO21HSV0 A1 A2 B Z VDD VSS
MM6 N14 B VSS VPW N12LL W=200.00n L=60.00n
MM1 N14 A1 N3 VPW N12LL W=200.00n L=60.00n
MM2 Z N14 VSS VPW N12LL W=200.00n L=60.00n
MMN1 N3 A2 VSS VPW N12LL W=200.00n L=60.00n
MM7 N13 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N13 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z N14 VDD VNW P12LL W=300.00n L=60.00n
MM0 N14 B N13 VNW P12LL W=300.00n L=60.00n
.ENDS AO21HSV0
****Sub-Circuit for AO21HSV1, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO21HSV1 A1 A2 B Z VDD VSS
MM6 N14 B VSS VPW N12LL W=200.00n L=60.00n
MM1 N14 A1 N3 VPW N12LL W=200.00n L=60.00n
MM2 Z N14 VSS VPW N12LL W=260.00n L=60.00n
MMN1 N3 A2 VSS VPW N12LL W=200.00n L=60.00n
MM7 N13 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N13 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z N14 VDD VNW P12LL W=410.00n L=60.00n
MM0 N14 B N13 VNW P12LL W=300.00n L=60.00n
.ENDS AO21HSV1
****Sub-Circuit for AO21HSV2, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO21HSV2 A1 A2 B Z VDD VSS
MM6 N14 B VSS VPW N12LL W=200.00n L=60.00n
MM1 N14 A1 N3 VPW N12LL W=200.00n L=60.00n
MM2 Z N14 VSS VPW N12LL W=430.00n L=60.00n
MMN1 N3 A2 VSS VPW N12LL W=200.00n L=60.00n
MM7 N13 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N13 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z N14 VDD VNW P12LL W=650.00n L=60.00n
MM0 N14 B N13 VNW P12LL W=300.00n L=60.00n
.ENDS AO21HSV2
****Sub-Circuit for AO21HSV4, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO21HSV4 A1 A2 B Z VDD VSS
MM6 N14 B VSS VPW N12LL W=350.00n L=60.00n
MM1 N14 A1 N3 VPW N12LL W=350.00n L=60.00n
MM2 Z N14 VSS VPW N12LL W=860.00n L=60.00n
MMN1 N3 A2 VSS VPW N12LL W=350.00n L=60.00n
MM7 N13 A1 VDD VNW P12LL W=520.00n L=60.00n
MM5 N13 A2 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z N14 VDD VNW P12LL W=1.3u L=60.00n
MM0 N14 B N13 VNW P12LL W=520.00n L=60.00n
.ENDS AO21HSV4
****Sub-Circuit for AO221HSV0, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO221HSV0 A1 A2 B1 B2 C Z VDD VSS
MM6 N8 C VSS VPW N12LL W=200.00n L=60.00n
MM9 N3 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 N8 A1 N14 VPW N12LL W=200.00n L=60.00n
MM2 Z N8 VSS VPW N12LL W=200.00n L=60.00n
MM4 N8 B1 N3 VPW N12LL W=200.00n L=60.00n
MMN1 N14 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 N9 B1 N11 VNW P12LL W=300.00n L=60.00n
MM7 N11 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N11 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z N8 VDD VNW P12LL W=300.00n L=60.00n
MM0 N9 B2 N11 VNW P12LL W=300.00n L=60.00n
MMP1 N8 C N9 VNW P12LL W=300.00n L=60.00n
.ENDS AO221HSV0
****Sub-Circuit for AO221HSV1, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO221HSV1 A1 A2 B1 B2 C Z VDD VSS
MM6 N8 C VSS VPW N12LL W=200.00n L=60.00n
MM9 N3 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 N8 A1 N14 VPW N12LL W=200.00n L=60.00n
MM2 Z N8 VSS VPW N12LL W=290.00n L=60.00n
MM4 N8 B1 N3 VPW N12LL W=200.00n L=60.00n
MMN1 N14 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 N9 B1 N11 VNW P12LL W=300.00n L=60.00n
MM7 N11 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N11 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z N8 VDD VNW P12LL W=440.00n L=60.00n
MM0 N9 B2 N11 VNW P12LL W=300.00n L=60.00n
MMP1 N8 C N9 VNW P12LL W=300.00n L=60.00n
.ENDS AO221HSV1
****Sub-Circuit for AO221HSV2, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO221HSV2 A1 A2 B1 B2 C Z VDD VSS
MM6 N8 C VSS VPW N12LL W=200.00n L=60.00n
MM9 N3 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 N8 A1 N14 VPW N12LL W=200.00n L=60.00n
MM2 Z N8 VSS VPW N12LL W=430.00n L=60.00n
MM4 N8 B1 N3 VPW N12LL W=200.00n L=60.00n
MMN1 N14 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 N9 B1 N11 VNW P12LL W=300.00n L=60.00n
MM7 N11 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N11 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z N8 VDD VNW P12LL W=650.00n L=60.00n
MM0 N9 B2 N11 VNW P12LL W=300.00n L=60.00n
MMP1 N8 C N9 VNW P12LL W=300.00n L=60.00n
.ENDS AO221HSV2
****Sub-Circuit for AO221HSV4, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO221HSV4 A1 A2 B1 B2 C Z VDD VSS
MM6 N8 C VSS VPW N12LL W=350.00n L=60.00n
MM9 N3 B2 VSS VPW N12LL W=350.00n L=60.00n
MM1 N8 A1 N14 VPW N12LL W=350.00n L=60.00n
MM2 Z N8 VSS VPW N12LL W=860.00n L=60.00n
MM4 N8 B1 N3 VPW N12LL W=350.00n L=60.00n
MMN1 N14 A2 VSS VPW N12LL W=350.00n L=60.00n
MM8 N9 B1 N11 VNW P12LL W=520.00n L=60.00n
MM7 N11 A1 VDD VNW P12LL W=520.00n L=60.00n
MM5 N11 A2 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z N8 VDD VNW P12LL W=1.3u L=60.00n
MM0 N9 B2 N11 VNW P12LL W=520.00n L=60.00n
MMP1 N8 C N9 VNW P12LL W=520.00n L=60.00n
.ENDS AO221HSV4
****Sub-Circuit for AO222HSV0, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO222HSV0 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM6 net3 C1 net4 VPW N12LL W=200.00n L=60.00n
MM10 net4 C2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 net3 A1 net6 VPW N12LL W=200.00n L=60.00n
MM2 Z net3 VSS VPW N12LL W=200.00n L=60.00n
MM4 net3 B1 net5 VPW N12LL W=200.00n L=60.00n
MMN1 net6 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM11 net3 C2 net2 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net3 VDD VNW P12LL W=300.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
MMP1 net3 C1 net2 VNW P12LL W=300.00n L=60.00n
.ENDS AO222HSV0
****Sub-Circuit for AO222HSV1, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO222HSV1 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM6 net3 C1 net4 VPW N12LL W=200.00n L=60.00n
MM10 net4 C2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 net3 A1 net6 VPW N12LL W=200.00n L=60.00n
MM2 Z net3 VSS VPW N12LL W=290.00n L=60.00n
MM4 net3 B1 net5 VPW N12LL W=200.00n L=60.00n
MMN1 net6 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM11 net3 C2 net2 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net3 VDD VNW P12LL W=440.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
MMP1 net3 C1 net2 VNW P12LL W=300.00n L=60.00n
.ENDS AO222HSV1
****Sub-Circuit for AO222HSV2, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO222HSV2 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM6 net3 C1 net4 VPW N12LL W=200.00n L=60.00n
MM10 net4 C2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 net3 A1 net6 VPW N12LL W=200.00n L=60.00n
MM2 Z net3 VSS VPW N12LL W=430.00n L=60.00n
MM4 net3 B1 net5 VPW N12LL W=200.00n L=60.00n
MMN1 net6 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM11 net3 C2 net2 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net3 VDD VNW P12LL W=650.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
MMP1 net3 C1 net2 VNW P12LL W=300.00n L=60.00n
.ENDS AO222HSV2
****Sub-Circuit for AO222HSV4, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO222HSV4 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM6 net3 C1 net4 VPW N12LL W=350.00n L=60.00n
MM10 net4 C2 VSS VPW N12LL W=350.00n L=60.00n
MM9 net5 B2 VSS VPW N12LL W=350.00n L=60.00n
MM1 net3 A1 net6 VPW N12LL W=350.00n L=60.00n
MM2 Z net3 VSS VPW N12LL W=860.00n L=60.00n
MM4 net3 B1 net5 VPW N12LL W=350.00n L=60.00n
MMN1 net6 A2 VSS VPW N12LL W=350.00n L=60.00n
MM8 net2 B2 net1 VNW P12LL W=520.00n L=60.00n
MM11 net3 C2 net2 VNW P12LL W=520.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=520.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z net3 VDD VNW P12LL W=1.3u L=60.00n
MM0 net2 B1 net1 VNW P12LL W=520.00n L=60.00n
MMP1 net3 C1 net2 VNW P12LL W=520.00n L=60.00n
.ENDS AO222HSV4
****Sub-Circuit for AO22HSV0, Wed Dec  8 11:21:13 CST 2010****
.SUBCKT AO22HSV0 A1 A2 B1 B2 Z VDD VSS
MM9 N64 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 N62 A1 N49 VPW N12LL W=200.00n L=60.00n
MM2 Z N62 VSS VPW N12LL W=200.00n L=60.00n
MM4 N62 B1 N64 VPW N12LL W=200.00n L=60.00n
MMN1 N49 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 N62 B2 N69 VNW P12LL W=300.00n L=60.00n
MM7 N69 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N69 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z N62 VDD VNW P12LL W=300.00n L=60.00n
MM0 N62 B1 N69 VNW P12LL W=300.00n L=60.00n
.ENDS AO22HSV0
****Sub-Circuit for AO22HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO22HSV1 A1 A2 B1 B2 Z VDD VSS
MM9 N64 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 N62 A1 N49 VPW N12LL W=200.00n L=60.00n
MM2 Z N62 VSS VPW N12LL W=290.00n L=60.00n
MM4 N62 B1 N64 VPW N12LL W=200.00n L=60.00n
MMN1 N49 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 N62 B2 N69 VNW P12LL W=300.00n L=60.00n
MM7 N69 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N69 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z N62 VDD VNW P12LL W=440.00n L=60.00n
MM0 N62 B1 N69 VNW P12LL W=300.00n L=60.00n
.ENDS AO22HSV1
****Sub-Circuit for AO22HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO22HSV2 A1 A2 B1 B2 Z VDD VSS
MM9 N64 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 N62 A1 N49 VPW N12LL W=200.00n L=60.00n
MM2 Z N62 VSS VPW N12LL W=430.00n L=60.00n
MM4 N62 B1 N64 VPW N12LL W=200.00n L=60.00n
MMN1 N49 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 N62 B2 N69 VNW P12LL W=300.00n L=60.00n
MM7 N69 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N69 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z N62 VDD VNW P12LL W=650.00n L=60.00n
MM0 N62 B1 N69 VNW P12LL W=300.00n L=60.00n
.ENDS AO22HSV2
****Sub-Circuit for AO22HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO22HSV4 A1 A2 B1 B2 Z VDD VSS
MM9 N64 B2 VSS VPW N12LL W=350.00n L=60.00n
MM1 N62 A1 N49 VPW N12LL W=350.00n L=60.00n
MM2 Z N62 VSS VPW N12LL W=860.00n L=60.00n
MM4 N62 B1 N64 VPW N12LL W=350.00n L=60.00n
MMN1 N49 A2 VSS VPW N12LL W=350.00n L=60.00n
MM8 N62 B2 N69 VNW P12LL W=520.00n L=60.00n
MM7 N69 A1 VDD VNW P12LL W=520.00n L=60.00n
MM5 N69 A2 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z N62 VDD VNW P12LL W=1.3u L=60.00n
MM0 N62 B1 N69 VNW P12LL W=520.00n L=60.00n
.ENDS AO22HSV4
****Sub-Circuit for AO31HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO31HSV0 A1 A2 A3 B Z VDD VSS
MM6 net2 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=300.00n L=60.00n
MM0 net2 B net1 VNW P12LL W=300.00n L=60.00n
.ENDS AO31HSV0
****Sub-Circuit for AO31HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO31HSV1 A1 A2 A3 B Z VDD VSS
MM6 net2 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=290.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=440.00n L=60.00n
MM0 net2 B net1 VNW P12LL W=300.00n L=60.00n
.ENDS AO31HSV1
****Sub-Circuit for AO31HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO31HSV2 A1 A2 A3 B Z VDD VSS
MM6 net2 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=430.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=650.00n L=60.00n
MM0 net2 B net1 VNW P12LL W=300.00n L=60.00n
.ENDS AO31HSV2
****Sub-Circuit for AO31HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO31HSV4 A1 A2 A3 B Z VDD VSS
MM6 net2 B VSS VPW N12LL W=350.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=350.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=860.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=350.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=520.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=520.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=1.3u L=60.00n
MM0 net2 B net1 VNW P12LL W=520.00n L=60.00n
.ENDS AO31HSV4
****Sub-Circuit for AO32HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO32HSV0 A1 A2 A3 B1 B2 Z VDD VSS
MM6 net2 B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=300.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AO32HSV0
****Sub-Circuit for AO32HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO32HSV1 A1 A2 A3 B1 B2 Z VDD VSS
MM6 net2 B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=290.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=440.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AO32HSV1
****Sub-Circuit for AO32HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO32HSV2 A1 A2 A3 B1 B2 Z VDD VSS
MM6 net2 B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=430.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=650.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AO32HSV2
****Sub-Circuit for AO32HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO32HSV4 A1 A2 A3 B1 B2 Z VDD VSS
MM6 net2 B1 net5 VPW N12LL W=350.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=350.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=860.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=350.00n L=60.00n
MM11 net5 B2 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=350.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=520.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=520.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=520.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=1.3u L=60.00n
MM0 net2 B1 net1 VNW P12LL W=520.00n L=60.00n
.ENDS AO32HSV4
****Sub-Circuit for AO33HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO33HSV0 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM12 net_69 B3 VSS VPW N12LL W=200.00n L=60.00n
MM6 net2 B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 net_69 VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=300.00n L=60.00n
MM13 net2 B3 net1 VNW P12LL W=300.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AO33HSV0
****Sub-Circuit for AO33HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO33HSV1 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM12 net_69 B3 VSS VPW N12LL W=200.00n L=60.00n
MM6 net2 B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=290.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 net_69 VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=440.00n L=60.00n
MM13 net2 B3 net1 VNW P12LL W=300.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AO33HSV1
****Sub-Circuit for AO33HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO33HSV2 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM12 net_69 B3 VSS VPW N12LL W=200.00n L=60.00n
MM6 net2 B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=430.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 net_69 VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=650.00n L=60.00n
MM13 net2 B3 net1 VNW P12LL W=300.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AO33HSV2
****Sub-Circuit for AO33HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AO33HSV4 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM12 net_69 B3 VSS VPW N12LL W=350.00n L=60.00n
MM6 net2 B1 net5 VPW N12LL W=350.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=350.00n L=60.00n
MM2 Z net2 VSS VPW N12LL W=860.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=350.00n L=60.00n
MM11 net5 B2 net_69 VPW N12LL W=350.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=350.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=520.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=520.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=520.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=520.00n L=60.00n
MM3 Z net2 VDD VNW P12LL W=1.3u L=60.00n
MM13 net2 B3 net1 VNW P12LL W=520.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=520.00n L=60.00n
.ENDS AO33HSV4
****Sub-Circuit for AOA211HSV0, Thu May 19 13:57:40 CST 2011****
.SUBCKT AOA211HSV0 A1 A2 B C Z VDD VSS
MMN1 net4 A2 VSS VPW N12LL W=180.00n L=60.00n
MM4 net_34 B VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net_38 VSS VPW N12LL W=200.00n L=60.00n
MM1 net_34 A1 net4 VPW N12LL W=180.00n L=60.00n
MM6 net_38 C net_34 VPW N12LL W=180.00n L=60.00n
MMP1 net_38 C VDD VNW P12LL W=200.00n L=60.00n
MM0 net_38 B net3 VNW P12LL W=200.00n L=60.00n
MM3 Z net_38 VDD VNW P12LL W=250.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=200.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=200.00n L=60.00n
.ENDS AOA211HSV0
****Sub-Circuit for AOA211HSV1, Thu May 19 13:57:40 CST 2011****
.SUBCKT AOA211HSV1 A1 A2 B C Z VDD VSS
MM0 net_42 B net3 VNW P12LL W=200.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=200.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=200.00n L=60.00n
MMP1 net_42 C VDD VNW P12LL W=200.00n L=60.00n
MM3 Z net_42 VDD VNW P12LL W=440.00n L=60.00n
MM1 net_26 A1 net4 VPW N12LL W=180.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=180.00n L=60.00n
MM4 net_26 B VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net_42 VSS VPW N12LL W=350.00n L=60.00n
MM6 net_42 C net_26 VPW N12LL W=180.00n L=60.00n
.ENDS AOA211HSV1
****Sub-Circuit for AOA211HSV2, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOA211HSV2 A1 A2 B C Z VDD VSS
MM0 net_42 B net3 VNW P12LL W=220.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=220.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=220.00n L=60.00n
MMP1 net_42 C VDD VNW P12LL W=220.00n L=60.00n
MM3 Z net_42 VDD VNW P12LL W=540.00n L=60.00n
MM1 net_26 A1 net4 VPW N12LL W=180.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=180.00n L=60.00n
MM4 net_26 B VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net_42 VSS VPW N12LL W=430.00n L=60.00n
MM6 net_42 C net_26 VPW N12LL W=180.00n L=60.00n
.ENDS AOA211HSV2
****Sub-Circuit for AOA211HSV4, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOA211HSV4 A1 A2 B C Z VDD VSS
MM0 net_42 B net3 VNW P12LL W=440.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=440.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 net_42 C VDD VNW P12LL W=440.00n L=60.00n
MM3 Z net_42 VDD VNW P12LL W=1.08u L=60.00n
MM1 net_26 A1 net4 VPW N12LL W=350.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=350.00n L=60.00n
MM4 net_26 B VSS VPW N12LL W=350.00n L=60.00n
MM2 Z net_42 VSS VPW N12LL W=860.00n L=60.00n
MM6 net_42 C net_26 VPW N12LL W=350.00n L=60.00n
.ENDS AOA211HSV4
****Sub-Circuit for AOAI211HSV0, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAI211HSV0 A1 A2 B C ZN VDD VSS
MM7 net3 A1 VDD VNW P12LL W=250.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=250.00n L=60.00n
MM0 ZN B net3 VNW P12LL W=250.00n L=60.00n
MMP1 ZN C VDD VNW P12LL W=250.00n L=60.00n
MM6 ZN C net_26 VPW N12LL W=200.00n L=60.00n
MM1 net_26 A1 net4 VPW N12LL W=200.00n L=60.00n
MM4 net_26 B VSS VPW N12LL W=200.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=200.00n L=60.00n
.ENDS AOAI211HSV0
****Sub-Circuit for AOAI211HSV1, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAI211HSV1 A1 A2 B C ZN VDD VSS
MMN1 net4 A2 VSS VPW N12LL W=350.00n L=60.00n
MM4 net_14 B VSS VPW N12LL W=350.00n L=60.00n
MM1 net_14 A1 net4 VPW N12LL W=350.00n L=60.00n
MM6 ZN C net_14 VPW N12LL W=350.00n L=60.00n
MMP1 ZN C VDD VNW P12LL W=440.00n L=60.00n
MM0 ZN B net3 VNW P12LL W=440.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=440.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=440.00n L=60.00n
.ENDS AOAI211HSV1
****Sub-Circuit for AOAI211HSV2, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAI211HSV2 A1 A2 B C ZN VDD VSS
MMN1 net4 A2 VSS VPW N12LL W=430.00n L=60.00n
MM4 net_14 B VSS VPW N12LL W=430.00n L=60.00n
MM1 net_14 A1 net4 VPW N12LL W=430.00n L=60.00n
MM6 ZN C net_14 VPW N12LL W=430.00n L=60.00n
MMP1 ZN C VDD VNW P12LL W=540.00n L=60.00n
MM0 ZN B net3 VNW P12LL W=540.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=540.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=540.00n L=60.00n
.ENDS AOAI211HSV2
****Sub-Circuit for AOAI211HSV4, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAI211HSV4 A1 A2 B C ZN VDD VSS
MMN1 net4 A2 VSS VPW N12LL W=860.00n L=60.00n
MM4 net_14 B VSS VPW N12LL W=860.00n L=60.00n
MM1 net_14 A1 net4 VPW N12LL W=860.00n L=60.00n
MM6 ZN C net_14 VPW N12LL W=860.00n L=60.00n
MMP1 ZN C VDD VNW P12LL W=1.08u L=60.00n
MM0 ZN B net3 VNW P12LL W=1.08u L=60.00n
MM5 net3 A2 VDD VNW P12LL W=1.08u L=60.00n
MM7 net3 A1 VDD VNW P12LL W=1.08u L=60.00n
.ENDS AOAI211HSV4
****Sub-Circuit for AOAOAOI211111HSV0, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAOAOI211111HSV0 A1 A2 B C D E F ZN VDD VSS
MM8 net_12 F VDD VNW P12LL W=250.00n L=60.00n
MM9 ZN E net_12 VNW P12LL W=250.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=250.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=250.00n L=60.00n
MM0 net_36 B net3 VNW P12LL W=250.00n L=60.00n
MMP1 net_36 C VDD VNW P12LL W=250.00n L=60.00n
MM2 net_12 D net_36 VNW P12LL W=250.00n L=60.00n
MM11 ZN E VSS VPW N12LL W=200.00n L=60.00n
MM10 ZN F net_45 VPW N12LL W=200.00n L=60.00n
MM6 net_45 C net_49 VPW N12LL W=200.00n L=60.00n
MM1 net_49 A1 net4 VPW N12LL W=200.00n L=60.00n
MM4 net_49 B VSS VPW N12LL W=200.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=200.00n L=60.00n
MM3 net_45 D VSS VPW N12LL W=200.00n L=60.00n
.ENDS AOAOAOI211111HSV0
****Sub-Circuit for AOAOAOI211111HSV1, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAOAOI211111HSV1 A1 A2 B C D E F ZN VDD VSS
MM3 net_25 D VSS VPW N12LL W=350.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=350.00n L=60.00n
MM4 net_21 B VSS VPW N12LL W=350.00n L=60.00n
MM1 net_21 A1 net4 VPW N12LL W=350.00n L=60.00n
MM6 net_25 C net_21 VPW N12LL W=350.00n L=60.00n
MM10 ZN F net_25 VPW N12LL W=350.00n L=60.00n
MM11 ZN E VSS VPW N12LL W=350.00n L=60.00n
MM2 net_64 D net_40 VNW P12LL W=440.00n L=60.00n
MMP1 net_40 C VDD VNW P12LL W=440.00n L=60.00n
MM0 net_40 B net3 VNW P12LL W=440.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=440.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=440.00n L=60.00n
MM8 net_64 F VDD VNW P12LL W=440.00n L=60.00n
MM9 ZN E net_64 VNW P12LL W=440.00n L=60.00n
.ENDS AOAOAOI211111HSV1
****Sub-Circuit for AOAOAOI211111HSV2, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAOAOI211111HSV2 A1 A2 B C D E F ZN VDD VSS
MM3 net_25 D VSS VPW N12LL W=430.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=430.00n L=60.00n
MM4 net_21 B VSS VPW N12LL W=430.00n L=60.00n
MM1 net_21 A1 net4 VPW N12LL W=430.00n L=60.00n
MM6 net_25 C net_21 VPW N12LL W=430.00n L=60.00n
MM10 ZN F net_25 VPW N12LL W=430.00n L=60.00n
MM11 ZN E VSS VPW N12LL W=430.00n L=60.00n
MM2 net_64 D net_40 VNW P12LL W=540.00n L=60.00n
MMP1 net_40 C VDD VNW P12LL W=540.00n L=60.00n
MM0 net_40 B net3 VNW P12LL W=540.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=540.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=540.00n L=60.00n
MM8 net_64 F VDD VNW P12LL W=540.00n L=60.00n
MM9 ZN E net_64 VNW P12LL W=540.00n L=60.00n
.ENDS AOAOAOI211111HSV2
****Sub-Circuit for AOAOAOI211111HSV4, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAOAOI211111HSV4 A1 A2 B C D E F ZN VDD VSS
MM3 net_25 D VSS VPW N12LL W=860.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=860.00n L=60.00n
MM4 net_21 B VSS VPW N12LL W=860.00n L=60.00n
MM1 net_21 A1 net4 VPW N12LL W=860.00n L=60.00n
MM6 net_25 C net_21 VPW N12LL W=860.00n L=60.00n
MM10 ZN F net_25 VPW N12LL W=860.00n L=60.00n
MM11 ZN E VSS VPW N12LL W=860.00n L=60.00n
MM2 net_64 D net_40 VNW P12LL W=1.08u L=60.00n
MMP1 net_40 C VDD VNW P12LL W=1.08u L=60.00n
MM0 net_40 B net3 VNW P12LL W=1.08u L=60.00n
MM5 net3 A2 VDD VNW P12LL W=1.08u L=60.00n
MM7 net3 A1 VDD VNW P12LL W=1.08u L=60.00n
MM8 net_64 F VDD VNW P12LL W=1.08u L=60.00n
MM9 ZN E net_64 VNW P12LL W=1.08u L=60.00n
.ENDS AOAOAOI211111HSV4
****Sub-Circuit for AOAOI2111HSV0, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAOI2111HSV0 A1 A2 B C D ZN VDD VSS
MM3 ZN D VSS VPW N12LL W=200.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 net_19 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net_19 A1 net4 VPW N12LL W=200.00n L=60.00n
MM6 ZN C net_19 VPW N12LL W=200.00n L=60.00n
MM2 ZN D net_30 VNW P12LL W=250.00n L=60.00n
MMP1 net_30 C VDD VNW P12LL W=250.00n L=60.00n
MM0 net_30 B net3 VNW P12LL W=250.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=250.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=250.00n L=60.00n
.ENDS AOAOI2111HSV0
****Sub-Circuit for AOAOI2111HSV1, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAOI2111HSV1 A1 A2 B C D ZN VDD VSS
MM7 net3 A1 VDD VNW P12LL W=440.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=440.00n L=60.00n
MM0 net_26 B net3 VNW P12LL W=440.00n L=60.00n
MMP1 net_26 C VDD VNW P12LL W=440.00n L=60.00n
MM2 ZN D net_26 VNW P12LL W=440.00n L=60.00n
MM6 ZN C net_31 VPW N12LL W=350.00n L=60.00n
MM1 net_31 A1 net4 VPW N12LL W=350.00n L=60.00n
MM4 net_31 B VSS VPW N12LL W=350.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=350.00n L=60.00n
MM3 ZN D VSS VPW N12LL W=350.00n L=60.00n
.ENDS AOAOI2111HSV1
****Sub-Circuit for AOAOI2111HSV2, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAOI2111HSV2 A1 A2 B C D ZN VDD VSS
MM7 net3 A1 VDD VNW P12LL W=540.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=540.00n L=60.00n
MM0 net_26 B net3 VNW P12LL W=540.00n L=60.00n
MMP1 net_26 C VDD VNW P12LL W=540.00n L=60.00n
MM2 ZN D net_26 VNW P12LL W=540.00n L=60.00n
MM6 ZN C net_31 VPW N12LL W=430.00n L=60.00n
MM1 net_31 A1 net4 VPW N12LL W=430.00n L=60.00n
MM4 net_31 B VSS VPW N12LL W=430.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=430.00n L=60.00n
MM3 ZN D VSS VPW N12LL W=430.00n L=60.00n
.ENDS AOAOI2111HSV2
****Sub-Circuit for AOAOI2111HSV4, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT AOAOI2111HSV4 A1 A2 B C D ZN VDD VSS
MM7 net3 A1 VDD VNW P12LL W=1.08u L=60.00n
MM5 net3 A2 VDD VNW P12LL W=1.08u L=60.00n
MM0 net_26 B net3 VNW P12LL W=1.08u L=60.00n
MMP1 net_26 C VDD VNW P12LL W=1.08u L=60.00n
MM2 ZN D net_26 VNW P12LL W=1.08u L=60.00n
MM6 ZN C net_31 VPW N12LL W=860.00n L=60.00n
MM1 net_31 A1 net4 VPW N12LL W=860.00n L=60.00n
MM4 net_31 B VSS VPW N12LL W=860.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=860.00n L=60.00n
MM3 ZN D VSS VPW N12LL W=860.00n L=60.00n
.ENDS AOAOI2111HSV4
****Sub-Circuit for AOI211HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI211HSV0 A1 A2 B C ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 net4 VPW N12LL W=200.00n L=60.00n
MM4 ZN C VSS VPW N12LL W=200.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=200.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=300.0n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=300.0n L=60.00n
MM0 net2 B net3 VNW P12LL W=300.0n L=60.00n
MMP1 ZN C net2 VNW P12LL W=300.0n L=60.00n
.ENDS AOI211HSV0
****Sub-Circuit for AOI211HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI211HSV1 A1 A2 B C ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 net4 VPW N12LL W=290.00n L=60.00n
MM4 ZN C VSS VPW N12LL W=290.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=290.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=440.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=440.00n L=60.00n
MM0 net2 B net3 VNW P12LL W=440.00n L=60.00n
MMP1 ZN C net2 VNW P12LL W=440.00n L=60.00n
.ENDS AOI211HSV1
****Sub-Circuit for AOI211HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI211HSV2 A1 A2 B C ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 net4 VPW N12LL W=430.00n L=60.00n
MM4 ZN C VSS VPW N12LL W=430.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=430.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=650.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=650.00n L=60.00n
MM0 net2 B net3 VNW P12LL W=650.00n L=60.00n
MMP1 ZN C net2 VNW P12LL W=650.00n L=60.00n
.ENDS AOI211HSV2
****Sub-Circuit for AOI211HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI211HSV4 A1 A2 B C ZN VDD VSS
MM8 net_51 net1 VSS VPW N12LL W=350.00n L=60.00n
MM6 net1 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net1 A1 net4 VPW N12LL W=200.00n L=60.00n
MM2 ZN net_51 VSS VPW N12LL W=860.00n L=60.00n
MM4 net1 C VSS VPW N12LL W=200.00n L=60.00n
MMN1 net4 A2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net_51 net1 VDD VNW P12LL W=530.00n L=60.00n
MM7 net3 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net3 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 ZN net_51 VDD VNW P12LL W=1.3u L=60.00n
MM0 net2 B net3 VNW P12LL W=300.00n L=60.00n
MMP1 net1 C net2 VNW P12LL W=300.00n L=60.00n
.ENDS AOI211HSV4
****Sub-Circuit for AOI21HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI21HSV0 A1 A2 B ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 N3 VPW N12LL W=200.00n L=60.00n
MMN1 N3 A2 VSS VPW N12LL W=200.00n L=60.00n
MM7 N13 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N13 A2 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B N13 VNW P12LL W=300.00n L=60.00n
.ENDS AOI21HSV0
****Sub-Circuit for AOI21HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI21HSV1 A1 A2 B ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 N3 VPW N12LL W=290.00n L=60.00n
MMN1 N3 A2 VSS VPW N12LL W=290.00n L=60.00n
MM7 N13 A1 VDD VNW P12LL W=440.00n L=60.00n
MM5 N13 A2 VDD VNW P12LL W=440.00n L=60.00n
MM0 ZN B N13 VNW P12LL W=440.00n L=60.00n
.ENDS AOI21HSV1
****Sub-Circuit for AOI21HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI21HSV2 A1 A2 B ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 N3 VPW N12LL W=430.00n L=60.00n
MMN1 N3 A2 VSS VPW N12LL W=430.00n L=60.00n
MM7 N13 A1 VDD VNW P12LL W=650.00n L=60.00n
MM5 N13 A2 VDD VNW P12LL W=650.00n L=60.00n
MM0 ZN B N13 VNW P12LL W=650.00n L=60.00n
.ENDS AOI21HSV2
****Sub-Circuit for AOI21HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI21HSV4 A1 A2 B ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=860.00n L=60.00n
MM1 ZN A1 N3 VPW N12LL W=860.00n L=60.00n
MMN1 N3 A2 VSS VPW N12LL W=860.00n L=60.00n
MM7 N13 A1 VDD VNW P12LL W=1.3u L=60.00n
MM5 N13 A2 VDD VNW P12LL W=1.3u L=60.00n
MM0 ZN B N13 VNW P12LL W=1.3u L=60.00n
.ENDS AOI21HSV4
****Sub-Circuit for AOI221HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI221HSV0 A1 A2 B1 B2 C ZN VDD VSS
MM6 ZN C VSS VPW N12LL W=200.00n L=60.00n
MM9 N3 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 N14 VPW N12LL W=200.00n L=60.00n
MM4 ZN B1 N3 VPW N12LL W=200.00n L=60.00n
MMN1 N14 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 N9 B1 N11 VNW P12LL W=300.0n L=60.00n
MM7 N11 A1 VDD VNW P12LL W=300.0n L=60.00n
MM5 N11 A2 VDD VNW P12LL W=300.0n L=60.00n
MM0 N9 B2 N11 VNW P12LL W=300.0n L=60.00n
MMP1 ZN C N9 VNW P12LL W=300.0n L=60.00n
.ENDS AOI221HSV0
****Sub-Circuit for AOI221HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI221HSV1 A1 A2 B1 B2 C ZN VDD VSS
MM6 ZN C VSS VPW N12LL W=290.00n L=60.00n
MM9 N3 B2 VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 N14 VPW N12LL W=290.00n L=60.00n
MM4 ZN B1 N3 VPW N12LL W=290.00n L=60.00n
MMN1 N14 A2 VSS VPW N12LL W=290.00n L=60.00n
MM8 N9 B1 N11 VNW P12LL W=440.00n L=60.00n
MM7 N11 A1 VDD VNW P12LL W=440.00n L=60.00n
MM5 N11 A2 VDD VNW P12LL W=440.00n L=60.00n
MM0 N9 B2 N11 VNW P12LL W=440.00n L=60.00n
MMP1 ZN C N9 VNW P12LL W=440.00n L=60.00n
.ENDS AOI221HSV1
****Sub-Circuit for AOI221HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI221HSV2 A1 A2 B1 B2 C ZN VDD VSS
MM6 ZN C VSS VPW N12LL W=430.00n L=60.00n
MM9 N3 B2 VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 N14 VPW N12LL W=430.00n L=60.00n
MM4 ZN B1 N3 VPW N12LL W=430.00n L=60.00n
MMN1 N14 A2 VSS VPW N12LL W=430.00n L=60.00n
MM8 N9 B1 N11 VNW P12LL W=650.00n L=60.00n
MM7 N11 A1 VDD VNW P12LL W=650.00n L=60.00n
MM5 N11 A2 VDD VNW P12LL W=650.00n L=60.00n
MM0 N9 B2 N11 VNW P12LL W=650.00n L=60.00n
MMP1 ZN C N9 VNW P12LL W=650.00n L=60.00n
.ENDS AOI221HSV2
****Sub-Circuit for AOI221HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI221HSV4 A1 A2 B1 B2 C ZN VDD VSS
MM10 net61 net77 VSS VPW N12LL W=350.00n L=60.00n
MM6 net77 C VSS VPW N12LL W=200.00n L=60.00n
MM9 N3 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 net77 A1 N14 VPW N12LL W=200.00n L=60.00n
MM2 ZN net61 VSS VPW N12LL W=860.00n L=60.00n
MM4 net77 B1 N3 VPW N12LL W=200.00n L=60.00n
MMN1 N14 A2 VSS VPW N12LL W=200.00n L=60.00n
MM11 net61 net77 VDD VNW P12LL W=530.00n L=60.00n
MM8 N9 B1 N11 VNW P12LL W=300.00n L=60.00n
MM7 N11 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 N11 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 ZN net61 VDD VNW P12LL W=1.3u L=60.00n
MM0 N9 B2 N11 VNW P12LL W=300.00n L=60.00n
MMP1 net77 C N9 VNW P12LL W=300.00n L=60.00n
.ENDS AOI221HSV4
****Sub-Circuit for AOI222HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI222HSV0 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM6 ZN C1 net4 VPW N12LL W=200.00n L=60.00n
MM10 net4 C2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 net6 VPW N12LL W=200.00n L=60.00n
MM4 ZN B1 net5 VPW N12LL W=200.00n L=60.00n
MMN1 net6 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 net2 B2 net1 VNW P12LL W=300.0n L=60.00n
MM11 ZN A2 net2 VNW P12LL W=300.0n L=60.00n
MM7 net1 C1 VDD VNW P12LL W=300.0n L=60.00n
MM5 net1 C2 VDD VNW P12LL W=300.0n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.0n L=60.00n
MMP1 ZN A1 net2 VNW P12LL W=300.0n L=60.00n
.ENDS AOI222HSV0
****Sub-Circuit for AOI222HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI222HSV1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM6 ZN C1 net4 VPW N12LL W=290.00n L=60.00n
MM10 net4 C2 VSS VPW N12LL W=290.00n L=60.00n
MM9 net5 B2 VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 net6 VPW N12LL W=290.00n L=60.00n
MM4 ZN B1 net5 VPW N12LL W=290.00n L=60.00n
MMN1 net6 A2 VSS VPW N12LL W=290.00n L=60.00n
MM8 net2 B2 net1 VNW P12LL W=440.0n L=60.00n
MM11 ZN A2 net2 VNW P12LL W=440.0n L=60.00n
MM7 net1 C1 VDD VNW P12LL W=440.0n L=60.00n
MM5 net1 C2 VDD VNW P12LL W=440.0n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=440.0n L=60.00n
MMP1 ZN A1 net2 VNW P12LL W=440.0n L=60.00n
.ENDS AOI222HSV1
****Sub-Circuit for AOI222HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI222HSV2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM6 ZN C1 net4 VPW N12LL W=430.00n L=60.00n
MM10 net4 C2 VSS VPW N12LL W=430.00n L=60.00n
MM9 net5 B2 VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 net6 VPW N12LL W=430.00n L=60.00n
MM4 ZN B1 net5 VPW N12LL W=430.00n L=60.00n
MMN1 net6 A2 VSS VPW N12LL W=430.00n L=60.00n
MM8 net2 B2 net1 VNW P12LL W=650.0n L=60.00n
MM11 ZN A2 net2 VNW P12LL W=650.0n L=60.00n
MM7 net1 C1 VDD VNW P12LL W=650.0n L=60.00n
MM5 net1 C2 VDD VNW P12LL W=650.0n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=650.0n L=60.00n
MMP1 ZN A1 net2 VNW P12LL W=650.0n L=60.00n
.ENDS AOI222HSV2
****Sub-Circuit for AOI222HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI222HSV4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM12 net_42 net3 VSS VPW N12LL W=350.00n L=60.00n
MM6 net3 C1 net4 VPW N12LL W=200.00n L=60.00n
MM10 net4 C2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 net3 A1 net6 VPW N12LL W=200.00n L=60.00n
MM2 ZN net_42 VSS VPW N12LL W=860.00n L=60.00n
MM4 net3 B1 net5 VPW N12LL W=200.00n L=60.00n
MMN1 net6 A2 VSS VPW N12LL W=200.00n L=60.00n
MM13 net_42 net3 VDD VNW P12LL W=530.00n L=60.00n
MM8 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM11 net3 C2 net2 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 ZN net_42 VDD VNW P12LL W=1.3u L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
MMP1 net3 C1 net2 VNW P12LL W=300.00n L=60.00n
.ENDS AOI222HSV4
****Sub-Circuit for AOI22HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI22HSV0 A1 A2 B1 B2 ZN VDD VSS
MM9 N64 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 N49 VPW N12LL W=200.00n L=60.00n
MM4 ZN B1 N64 VPW N12LL W=200.00n L=60.00n
MMN1 N49 A2 VSS VPW N12LL W=200.00n L=60.00n
MM8 ZN B2 N69 VNW P12LL W=300.00n L=60.00n
MM7 N69 A2 VDD VNW P12LL W=300.00n L=60.00n
MM5 N69 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 N69 VNW P12LL W=300.00n L=60.00n
.ENDS AOI22HSV0
****Sub-Circuit for AOI22HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI22HSV1 A1 A2 B1 B2 ZN VDD VSS
MM9 N64 B2 VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 N49 VPW N12LL W=290.00n L=60.00n
MM4 ZN B1 N64 VPW N12LL W=290.00n L=60.00n
MMN1 N49 A2 VSS VPW N12LL W=290.00n L=60.00n
MM8 ZN B2 N69 VNW P12LL W=440.00n L=60.00n
MM7 N69 A2 VDD VNW P12LL W=440.00n L=60.00n
MM5 N69 A1 VDD VNW P12LL W=440.00n L=60.00n
MM0 ZN B1 N69 VNW P12LL W=440.00n L=60.00n
.ENDS AOI22HSV1
****Sub-Circuit for AOI22HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI22HSV2 A1 A2 B1 B2 ZN VDD VSS
MM9 N64 B2 VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 N49 VPW N12LL W=430.00n L=60.00n
MM4 ZN B1 N64 VPW N12LL W=430.00n L=60.00n
MMN1 N49 A2 VSS VPW N12LL W=430.00n L=60.00n
MM8 ZN B2 N69 VNW P12LL W=650.00n L=60.00n
MM7 N69 A2 VDD VNW P12LL W=650.00n L=60.00n
MM5 N69 A1 VDD VNW P12LL W=650.00n L=60.00n
MM0 ZN B1 N69 VNW P12LL W=650.00n L=60.00n
.ENDS AOI22HSV2
****Sub-Circuit for AOI22HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI22HSV4 A1 A2 B1 B2 ZN VDD VSS
MM9 N64 B2 VSS VPW N12LL W=860.00n L=60.00n
MM1 ZN A1 N49 VPW N12LL W=860.00n L=60.00n
MM4 ZN B1 N64 VPW N12LL W=860.00n L=60.00n
MMN1 N49 A2 VSS VPW N12LL W=860.00n L=60.00n
MM8 ZN B2 N69 VNW P12LL W=1.3u L=60.00n
MM7 N69 A2 VDD VNW P12LL W=1.3u L=60.00n
MM5 N69 A1 VDD VNW P12LL W=1.3u L=60.00n
MM0 ZN B1 N69 VNW P12LL W=1.3u L=60.00n
.ENDS AOI22HSV4
****Sub-Circuit for AOI31HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI31HSV0 A1 A2 A3 B ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 net3 VPW N12LL W=200.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B net1 VNW P12LL W=300.00n L=60.00n
.ENDS AOI31HSV0
****Sub-Circuit for AOI31HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI31HSV1 A1 A2 A3 B ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 net3 VPW N12LL W=290.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=290.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=440.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=440.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=440.00n L=60.00n
MM0 ZN B net1 VNW P12LL W=440.00n L=60.00n
.ENDS AOI31HSV1
****Sub-Circuit for AOI31HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI31HSV2 A1 A2 A3 B ZN VDD VSS
MM6 ZN B VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 net3 VPW N12LL W=430.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=430.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=650.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=650.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=650.00n L=60.00n
MM0 ZN B net1 VNW P12LL W=650.00n L=60.00n
.ENDS AOI31HSV2
****Sub-Circuit for AOI31HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI31HSV4 A1 A2 A3 B ZN VDD VSS
MM10 net_49 net2 VSS VPW N12LL W=350.00n L=60.00n
MM6 net2 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 ZN net_49 VSS VPW N12LL W=860.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM11 net_49 net2 VDD VNW P12LL W=530.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 ZN net_49 VDD VNW P12LL W=1.3u L=60.00n
MM0 net2 B net1 VNW P12LL W=300.00n L=60.00n
.ENDS AOI31HSV4
****Sub-Circuit for AOI32HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI32HSV0 A1 A2 A3 B1 B2 ZN VDD VSS
MM6 ZN B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 net3 VPW N12LL W=200.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 ZN B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AOI32HSV0
****Sub-Circuit for AOI32HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI32HSV1 A1 A2 A3 B1 B2 ZN VDD VSS
MM6 ZN B1 net5 VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 net3 VPW N12LL W=290.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=290.00n L=60.00n
MM11 net5 B2 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=290.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=440.00n L=60.00n
MM10 ZN B2 net1 VNW P12LL W=440.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=440.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=440.00n L=60.00n
MM0 ZN B1 net1 VNW P12LL W=440.00n L=60.00n
.ENDS AOI32HSV1
****Sub-Circuit for AOI32HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI32HSV2 A1 A2 A3 B1 B2 ZN VDD VSS
MM6 ZN B1 net5 VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 net3 VPW N12LL W=430.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=430.00n L=60.00n
MM11 net5 B2 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=430.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=650.00n L=60.00n
MM10 ZN B2 net1 VNW P12LL W=650.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=650.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=650.00n L=60.00n
MM0 ZN B1 net1 VNW P12LL W=650.00n L=60.00n
.ENDS AOI32HSV2
****Sub-Circuit for AOI32HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI32HSV4 A1 A2 A3 B1 B2 ZN VDD VSS
MM12 net_56 net2 VSS VPW N12LL W=350.00n L=60.00n
MM6 net2 B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 ZN net_56 VSS VPW N12LL W=860.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM13 net_56 net2 VDD VNW P12LL W=530.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 ZN net_56 VDD VNW P12LL W=1.3u L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AOI32HSV4
****Sub-Circuit for AOI33HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI33HSV0 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM12 net_69 B3 VSS VPW N12LL W=200.00n L=60.00n
MM6 ZN B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 net3 VPW N12LL W=200.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 net_69 VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 ZN B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM13 ZN B3 net1 VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AOI33HSV0
****Sub-Circuit for AOI33HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI33HSV1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM12 net_69 B3 VSS VPW N12LL W=290.00n L=60.00n
MM6 ZN B1 net5 VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 net3 VPW N12LL W=290.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=290.00n L=60.00n
MM11 net5 B2 net_69 VPW N12LL W=290.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=290.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=440.00n L=60.00n
MM10 ZN B2 net1 VNW P12LL W=440.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=440.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=440.00n L=60.00n
MM13 ZN B3 net1 VNW P12LL W=440.00n L=60.00n
MM0 ZN B1 net1 VNW P12LL W=440.00n L=60.00n
.ENDS AOI33HSV1
****Sub-Circuit for AOI33HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI33HSV2 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM12 net_69 B3 VSS VPW N12LL W=430.00n L=60.00n
MM6 ZN B1 net5 VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 net3 VPW N12LL W=430.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=430.00n L=60.00n
MM11 net5 B2 net_69 VPW N12LL W=430.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=430.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=650.00n L=60.00n
MM10 ZN B2 net1 VNW P12LL W=650.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=650.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=650.00n L=60.00n
MM13 ZN B3 net1 VNW P12LL W=650.00n L=60.00n
MM0 ZN B1 net1 VNW P12LL W=650.00n L=60.00n
.ENDS AOI33HSV2
****Sub-Circuit for AOI33HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT AOI33HSV4 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM14 net_068 net2 VSS VPW N12LL W=350.00n L=60.00n
MM12 net_69 B3 VSS VPW N12LL W=200.00n L=60.00n
MM6 net2 B1 net5 VPW N12LL W=200.00n L=60.00n
MM1 net2 A1 net3 VPW N12LL W=200.00n L=60.00n
MM2 ZN net_068 VSS VPW N12LL W=860.00n L=60.00n
MM9 net4 A3 VSS VPW N12LL W=200.00n L=60.00n
MM11 net5 B2 net_69 VPW N12LL W=200.00n L=60.00n
MMN1 net3 A2 net4 VPW N12LL W=200.00n L=60.00n
MM15 net_068 net2 VDD VNW P12LL W=530.00n L=60.00n
MM8 net1 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net2 B2 net1 VNW P12LL W=300.00n L=60.00n
MM7 net1 A1 VDD VNW P12LL W=300.00n L=60.00n
MM5 net1 A2 VDD VNW P12LL W=300.00n L=60.00n
MM3 ZN net_068 VDD VNW P12LL W=1.3u L=60.00n
MM13 net2 B3 net1 VNW P12LL W=300.00n L=60.00n
MM0 net2 B1 net1 VNW P12LL W=300.00n L=60.00n
.ENDS AOI33HSV4
****Sub-Circuit for BENCHSV1, Thu May 19 13:57:40 CST 2011****
.SUBCKT BENCHSV1 A MI0 MI1 MI2 S X2 VDD VSS
MM21 X2 net112 VSS VPW N12LL W=350n L=60.0n
MM17 S net102 VSS VPW N12LL W=350n L=60.0n
MM19 A net104 VSS VPW N12LL W=350n L=60.0n
MM15 net106 MI1 net93 VPW N12LL W=180n L=60.0n
MM23 net100 MI2 VSS VPW N12LL W=220n L=60.0n
MM8 net60 MI2 net78 VPW N12LL W=180n L=60.0n
MM9 net78 net110 VSS VPW N12LL W=250n L=60.0n
MM10 net78 net108 VSS VPW N12LL W=250n L=60.0n
MM25 net102 net60 VSS VPW N12LL W=180n L=60.0n
MM11 net63 net100 net87 VPW N12LL W=180n L=60.0n
MM27 net104 net63 VSS VPW N12LL W=180n L=60.0n
MM29 net106 net110 VSS VPW N12LL W=180n L=60.0n
MM31 net108 MI1 VSS VPW N12LL W=280n L=60.0n
MM33 net110 MI0 VSS VPW N12LL W=280n L=60.0n
MM35 net112 net93 VSS VPW N12LL W=180n L=60.0n
MM12 net87 MI0 VSS VPW N12LL W=250n L=60.0n
MM13 net87 MI1 VSS VPW N12LL W=250n L=60.0n
MM14 net110 net108 net93 VPW N12LL W=180n L=60.0n
MM0 net_0272 net108 VDD VNW P12LL W=200n L=60.0n
MM1 net60 net110 net_0272 VNW P12LL W=200n L=60.0n
MM3 net63 MI0 net_0236 VNW P12LL W=200n L=60.0n
MM4 net60 MI2 VDD VNW P12LL W=200n L=60.0n
MM18 A net104 VDD VNW P12LL W=440n L=60.0n
MM5 net63 net100 VDD VNW P12LL W=200n L=60.0n
MM6 net110 MI1 net93 VNW P12LL W=220n L=60.0n
MM16 S net102 VDD VNW P12LL W=440n L=60.0n
MM7 net106 net108 net93 VNW P12LL W=220n L=60.0n
MM22 net100 MI2 VDD VNW P12LL W=270n L=60.0n
MM2 net_0236 MI1 VDD VNW P12LL W=200n L=60.0n
MM24 net102 net60 VDD VNW P12LL W=220n L=60.0n
MM26 net104 net63 VDD VNW P12LL W=220n L=60.0n
MM20 X2 net112 VDD VNW P12LL W=440n L=60.0n
MM28 net106 net110 VDD VNW P12LL W=220n L=60.0n
MM30 net108 MI1 VDD VNW P12LL W=350n L=60.0n
MM32 net110 MI0 VDD VNW P12LL W=350n L=60.0n
MM34 net112 net93 VDD VNW P12LL W=220n L=60.0n
.ENDS BENCHSV1
****Sub-Circuit for BENCHSV2, Wed Feb 16 10:30:57 CST 2011****
.SUBCKT BENCHSV2 A MI0 MI1 MI2 S X2 VDD VSS
MM21 X2 net112 VSS VPW N12LL W=430n L=60.0n
MM17 S net102 VSS VPW N12LL W=430n L=60.0n
MM19 A net104 VSS VPW N12LL W=430n L=60.0n
MM15 net106 MI1 net93 VPW N12LL W=220n L=60.0n
MM23 net100 MI2 VSS VPW N12LL W=280n L=60.0n
MM8 net60 MI2 net78 VPW N12LL W=180n L=60.0n
MM9 net78 net110 VSS VPW N12LL W=320n L=60.0n
MM10 net78 net108 VSS VPW N12LL W=320n L=60.0n
MM25 net102 net60 VSS VPW N12LL W=220n L=60.0n
MM11 net63 net100 net87 VPW N12LL W=180n L=60.0n
MM27 net104 net63 VSS VPW N12LL W=220n L=60.0n
MM29 net106 net110 VSS VPW N12LL W=220n L=60.0n
MM31 net108 MI1 VSS VPW N12LL W=350n L=60.0n
MM33 net110 MI0 VSS VPW N12LL W=350n L=60.0n
MM35 net112 net93 VSS VPW N12LL W=220n L=60.0n
MM12 net87 MI0 VSS VPW N12LL W=320n L=60.0n
MM13 net87 MI1 VSS VPW N12LL W=320n L=60.0n
MM14 net110 net108 net93 VPW N12LL W=220n L=60.0n
MM0 net_0216 net108 VDD VNW P12LL W=220n L=60.0n
MM1 net60 net110 net_0216 VNW P12LL W=220n L=60.0n
MM3 net63 MI0 net_0220 VNW P12LL W=220n L=60.0n
MM4 net60 MI2 VDD VNW P12LL W=220n L=60.0n
MM18 A net104 VDD VNW P12LL W=540n L=60.0n
MM5 net63 net100 VDD VNW P12LL W=220n L=60.0n
MM6 net110 MI1 net93 VNW P12LL W=270n L=60.0n
MM16 S net102 VDD VNW P12LL W=540n L=60.0n
MM7 net106 net108 net93 VNW P12LL W=270n L=60.0n
MM22 net100 MI2 VDD VNW P12LL W=350n L=60.0n
MM2 net_0220 MI1 VDD VNW P12LL W=220n L=60.0n
MM24 net102 net60 VDD VNW P12LL W=270n L=60.0n
MM26 net104 net63 VDD VNW P12LL W=270n L=60.0n
MM20 X2 net112 VDD VNW P12LL W=540n L=60.0n
MM28 net106 net110 VDD VNW P12LL W=270n L=60.0n
MM30 net108 MI1 VDD VNW P12LL W=440n L=60.0n
MM32 net110 MI0 VDD VNW P12LL W=440n L=60.0n
MM34 net112 net93 VDD VNW P12LL W=270n L=60.0n
.ENDS BENCHSV2
****Sub-Circuit for BENCHSV4, Wed Feb 16 10:30:57 CST 2011****
.SUBCKT BENCHSV4 A MI0 MI1 MI2 S X2 VDD VSS
MM21 X2 net112 VSS VPW N12LL W=860n L=60.0n
MM17 S net102 VSS VPW N12LL W=860n L=60.0n
MM19 A net104 VSS VPW N12LL W=860n L=60.0n
MM15 net106 MI1 net93 VPW N12LL W=350n L=60.0n
MM23 net100 MI2 VSS VPW N12LL W=350n L=60.0n
MM8 net60 MI2 net78 VPW N12LL W=350n L=60.0n
MM9 net78 net110 VSS VPW N12LL W=430n L=60.0n
MM10 net78 net108 VSS VPW N12LL W=430n L=60.0n
MM25 net102 net60 VSS VPW N12LL W=430n L=60.0n
MM11 net63 net100 net87 VPW N12LL W=350n L=60.0n
MM27 net104 net63 VSS VPW N12LL W=430n L=60.0n
MM29 net106 net110 VSS VPW N12LL W=350n L=60.0n
MM31 net108 MI1 VSS VPW N12LL W=430n L=60.0n
MM33 net110 MI0 VSS VPW N12LL W=430n L=60.0n
MM35 net112 net93 VSS VPW N12LL W=430n L=60.0n
MM12 net87 MI0 VSS VPW N12LL W=430n L=60.0n
MM13 net87 MI1 VSS VPW N12LL W=430n L=60.0n
MM14 net110 net108 net93 VPW N12LL W=350n L=60.0n
MM0 net_0216 net108 VDD VNW P12LL W=440n L=60.0n
MM1 net60 net110 net_0216 VNW P12LL W=440n L=60.0n
MM3 net63 MI0 net_0220 VNW P12LL W=440n L=60.0n
MM4 net60 MI2 VDD VNW P12LL W=440n L=60.0n
MM18 A net104 VDD VNW P12LL W=1.08u L=60.0n
MM5 net63 net100 VDD VNW P12LL W=440n L=60.0n
MM6 net110 MI1 net93 VNW P12LL W=440n L=60.0n
MM16 S net102 VDD VNW P12LL W=1.08u L=60.0n
MM7 net106 net108 net93 VNW P12LL W=440n L=60.0n
MM22 net100 MI2 VDD VNW P12LL W=440n L=60.0n
MM2 net_0220 MI1 VDD VNW P12LL W=440n L=60.0n
MM24 net102 net60 VDD VNW P12LL W=540n L=60.0n
MM26 net104 net63 VDD VNW P12LL W=540n L=60.0n
MM20 X2 net112 VDD VNW P12LL W=1.08u L=60.0n
MM28 net106 net110 VDD VNW P12LL W=440n L=60.0n
MM30 net108 MI1 VDD VNW P12LL W=540n L=60.0n
MM32 net110 MI0 VDD VNW P12LL W=540n L=60.0n
MM34 net112 net93 VDD VNW P12LL W=540n L=60.0n
.ENDS BENCHSV4
****Sub-Circuit for BMUXHSV1, Wed Mar  9 14:52:41 CST 2011****
.SUBCKT BMUXHSV1 A MI0 MI1 PP S X2 VDD VSS
MM7 net64 MI0 VSS VPW N12LL W=180n L=60.0n
MM9 net66 A VSS VPW N12LL W=290n L=60.0n
MM11 net68 S VSS VPW N12LL W=290n L=60.0n
MM1 net58 net103 VSS VPW N12LL W=180n L=60.0n
MM13 PP net109 VSS VPW N12LL W=350n L=60.0n
MM5 net62 MI1 VSS VPW N12LL W=180n L=60.0n
MM22 net68 net62 net97 VPW N12LL W=220n L=60.0n
MM23 net66 MI1 net97 VPW N12LL W=220n L=60.0n
MM24 net68 net64 net103 VPW N12LL W=220n L=60.0n
MM15 net89 X2 VSS VPW N12LL W=180n L=60.0n
MM25 net66 MI0 net103 VPW N12LL W=220n L=60.0n
MM26 net60 net89 net109 VPW N12LL W=180n L=60.0n
MM27 net58 X2 net109 VPW N12LL W=180n L=60.0n
MM3 net60 net97 VSS VPW N12LL W=180n L=60.0n
MM6 net64 MI0 VDD VNW P12LL W=220n L=60.0n
MM8 net66 A VDD VNW P12LL W=360n L=60.0n
MM2 net60 net97 VDD VNW P12LL W=220n L=60.0n
MM10 net68 S VDD VNW P12LL W=360n L=60.0n
MM19 net66 net64 net103 VNW P12LL W=270n L=60.0n
MM12 PP net109 VDD VNW P12LL W=440n L=60.0n
MM20 net60 X2 net109 VNW P12LL W=220n L=60.0n
MM14 net89 X2 VDD VNW P12LL W=220n L=60.0n
MM21 net58 net89 net109 VNW P12LL W=220n L=60.0n
MM0 net58 net103 VDD VNW P12LL W=220n L=60.0n
MM4 net62 MI1 VDD VNW P12LL W=220n L=60.0n
MM16 net68 MI1 net97 VNW P12LL W=270n L=60.0n
MM17 net66 net62 net97 VNW P12LL W=270n L=60.0n
MM18 net68 MI0 net103 VNW P12LL W=270n L=60.0n
.ENDS BMUXHSV1
****Sub-Circuit for BMUXHSV2, Wed Mar  9 14:52:41 CST 2011****
.SUBCKT BMUXHSV2 A MI0 MI1 PP S X2 VDD VSS
MM7 net64 MI0 VSS VPW N12LL W=220n L=60.0n
MM9 net66 A VSS VPW N12LL W=350n L=60.0n
MM11 net68 S VSS VPW N12LL W=350n L=60.0n
MM1 net58 net103 VSS VPW N12LL W=220n L=60.0n
MM13 PP net109 VSS VPW N12LL W=430n L=60.0n
MM5 net62 MI1 VSS VPW N12LL W=220n L=60.0n
MM22 net68 net62 net97 VPW N12LL W=290n L=60.0n
MM23 net66 MI1 net97 VPW N12LL W=290n L=60.0n
MM24 net68 net64 net103 VPW N12LL W=290n L=60.0n
MM15 net89 X2 VSS VPW N12LL W=220n L=60.0n
MM25 net66 MI0 net103 VPW N12LL W=290n L=60.0n
MM26 net60 net89 net109 VPW N12LL W=220n L=60.0n
MM27 net58 X2 net109 VPW N12LL W=220n L=60.0n
MM3 net60 net97 VSS VPW N12LL W=220n L=60.0n
MM6 net64 MI0 VDD VNW P12LL W=270n L=60.0n
MM8 net66 A VDD VNW P12LL W=440n L=60.0n
MM2 net60 net97 VDD VNW P12LL W=270n L=60.0n
MM10 net68 S VDD VNW P12LL W=440n L=60.0n
MM19 net66 net64 net103 VNW P12LL W=360n L=60.0n
MM12 PP net109 VDD VNW P12LL W=540n L=60.0n
MM20 net60 X2 net109 VNW P12LL W=270n L=60.0n
MM14 net89 X2 VDD VNW P12LL W=270n L=60.0n
MM21 net58 net89 net109 VNW P12LL W=270n L=60.0n
MM0 net58 net103 VDD VNW P12LL W=270n L=60.0n
MM4 net62 MI1 VDD VNW P12LL W=270n L=60.0n
MM16 net68 MI1 net97 VNW P12LL W=360n L=60.0n
MM17 net66 net62 net97 VNW P12LL W=360n L=60.0n
MM18 net68 MI0 net103 VNW P12LL W=360n L=60.0n
.ENDS BMUXHSV2
****Sub-Circuit for BMUXHSV4, Wed Mar  9 14:52:41 CST 2011****
.SUBCKT BMUXHSV4 A MI0 MI1 PP S X2 VDD VSS
MM7 net64 MI0 VSS VPW N12LL W=220n L=60.0n
MM9 net66 A VSS VPW N12LL W=430n L=60.0n
MM11 net68 S VSS VPW N12LL W=430n L=60.0n
MM1 net58 net103 VSS VPW N12LL W=350n L=60.0n
MM13 PP net109 VSS VPW N12LL W=860n L=60.0n
MM5 net62 MI1 VSS VPW N12LL W=220n L=60.0n
MM22 net68 net62 net97 VPW N12LL W=430n L=60.0n
MM23 net66 MI1 net97 VPW N12LL W=430n L=60.0n
MM24 net68 net64 net103 VPW N12LL W=430n L=60.0n
MM15 net89 X2 VSS VPW N12LL W=220n L=60.0n
MM25 net66 MI0 net103 VPW N12LL W=430n L=60.0n
MM26 net60 net89 net109 VPW N12LL W=350n L=60.0n
MM27 net58 X2 net109 VPW N12LL W=350n L=60.0n
MM3 net60 net97 VSS VPW N12LL W=350n L=60.0n
MM6 net64 MI0 VDD VNW P12LL W=270n L=60.0n
MM8 net66 A VDD VNW P12LL W=540n L=60.0n
MM2 net60 net97 VDD VNW P12LL W=440n L=60.0n
MM10 net68 S VDD VNW P12LL W=540n L=60.0n
MM19 net66 net64 net103 VNW P12LL W=540n L=60.0n
MM12 PP net109 VDD VNW P12LL W=1.08u L=60.0n
MM20 net60 X2 net109 VNW P12LL W=440n L=60.0n
MM14 net89 X2 VDD VNW P12LL W=270n L=60.0n
MM21 net58 net89 net109 VNW P12LL W=440n L=60.0n
MM0 net58 net103 VDD VNW P12LL W=440n L=60.0n
MM4 net62 MI1 VDD VNW P12LL W=270n L=60.0n
MM16 net68 MI1 net97 VNW P12LL W=540n L=60.0n
MM17 net66 net62 net97 VNW P12LL W=540n L=60.0n
MM18 net68 MI0 net103 VNW P12LL W=540n L=60.0n
.ENDS BMUXHSV4
****Sub-Circuit for BUFHSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV0 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=200.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=300.00n L=60.00n
.ENDS BUFHSV0
****Sub-Circuit for BUFHSV0RT, Thu May 19 13:57:40 CST 2011****
.SUBCKT BUFHSV0RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=250.00n L=60.00n
MM3 net11 I VDD VNW P12LL W=200.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=180.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=200.00n L=60.00n
.ENDS BUFHSV0RT
****Sub-Circuit for BUFHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV1 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=290.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=440.00n L=60.00n
.ENDS BUFHSV1
****Sub-Circuit for BUFHSV12, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV12 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=1.02u L=60.00n
MM2 Z net13 VSS VPW N12LL W=2.58u L=60.00n
MM1 net13 I VDD VNW P12LL W=1.53u L=60.00n
MM3 Z net13 VDD VNW P12LL W=3.9u L=60.00n
.ENDS BUFHSV12
****Sub-Circuit for BUFHSV12RO, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV12RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=2.58u L=60.00n
MM2 net7 I VSS VPW N12LL W=320.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=400.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=3.24u L=60.00n
.ENDS BUFHSV12RO
****Sub-Circuit for BUFHSV12RQ, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV12RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=2.58u L=60.00n
MM2 net7 I VSS VPW N12LL W=640.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=800.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=3.24u L=60.00n
.ENDS BUFHSV12RQ
****Sub-Circuit for BUFHSV12RT, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV12RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=3.24u L=60.00n
MM3 net11 I VDD VNW P12LL W=1.08u L=60.00n
MM2 net11 I VSS VPW N12LL W=860.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=2.58u L=60.00n
.ENDS BUFHSV12RT
****Sub-Circuit for BUFHSV16, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV16 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=1.29u L=60.00n
MM2 Z net13 VSS VPW N12LL W=3.44u L=60.00n
MM1 net13 I VDD VNW P12LL W=1.95u L=60.00n
MM3 Z net13 VDD VNW P12LL W=5.2u L=60.00n
.ENDS BUFHSV16
****Sub-Circuit for BUFHSV16RO, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV16RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=3.44u L=60.00n
MM2 net7 I VSS VPW N12LL W=430.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=540.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=4.32u L=60.00n
.ENDS BUFHSV16RO
****Sub-Circuit for BUFHSV16RQ, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV16RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=3.44u L=60.00n
MM2 net7 I VSS VPW N12LL W=860.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=1.08u L=60.00n
MM0 Z net7 VDD VNW P12LL W=4.32u L=60.00n
.ENDS BUFHSV16RQ
****Sub-Circuit for BUFHSV16RT, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV16RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=4.32u L=60.00n
MM3 net11 I VDD VNW P12LL W=1.44u L=60.00n
MM2 net11 I VSS VPW N12LL W=1.14u L=60.00n
MM1 Z net11 VSS VPW N12LL W=3.44u L=60.00n
.ENDS BUFHSV16RT
****Sub-Circuit for BUFHSV1RT, Thu May 19 13:57:40 CST 2011****
.SUBCKT BUFHSV1RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=440.00n L=60.00n
MM3 net11 I VDD VNW P12LL W=200.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=180.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=350.00n L=60.00n
.ENDS BUFHSV1RT
****Sub-Circuit for BUFHSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV2 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=430.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=300.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=650.00n L=60.00n
.ENDS BUFHSV2
****Sub-Circuit for BUFHSV20, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV20 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=1.72u L=60.00n
MM2 Z net13 VSS VPW N12LL W=4.3u L=60.00n
MM1 net13 I VDD VNW P12LL W=2.6u L=60.00n
MM3 Z net13 VDD VNW P12LL W=6.5u L=60.00n
.ENDS BUFHSV20
****Sub-Circuit for BUFHSV20RO, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV20RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=4.3u L=60.00n
MM2 net7 I VSS VPW N12LL W=540.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=680.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=5.4u L=60.00n
.ENDS BUFHSV20RO
****Sub-Circuit for BUFHSV20RQ, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV20RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=4.3u L=60.00n
MM2 net7 I VSS VPW N12LL W=1.07u L=60.00n
MM3 net7 I VDD VNW P12LL W=1.34u L=60.00n
MM0 Z net7 VDD VNW P12LL W=5.4u L=60.00n
.ENDS BUFHSV20RQ
****Sub-Circuit for BUFHSV20RT, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV20RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=5.4u L=60.00n
MM3 net11 I VDD VNW P12LL W=1.8u L=60.00n
MM2 net11 I VSS VPW N12LL W=1.43u L=60.00n
MM1 Z net11 VSS VPW N12LL W=4.3u L=60.00n
.ENDS BUFHSV20RT
****Sub-Circuit for BUFHSV24, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV24 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=2.05u L=60.00n
MM2 Z net13 VSS VPW N12LL W=5.16u L=60.00n
MM1 net13 I VDD VNW P12LL W=3.05u L=60.00n
MM3 Z net13 VDD VNW P12LL W=7.8u L=60.00n
.ENDS BUFHSV24
****Sub-Circuit for BUFHSV24RO, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV24RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=5.16u L=60.00n
MM2 net7 I VSS VPW N12LL W=640.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=800.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=6.48u L=60.00n
.ENDS BUFHSV24RO
****Sub-Circuit for BUFHSV24RQ, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV24RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=5.16u L=60.00n
MM2 net7 I VSS VPW N12LL W=1.29u L=60.00n
MM3 net7 I VDD VNW P12LL W=1.62u L=60.00n
MM0 Z net7 VDD VNW P12LL W=6.48u L=60.00n
.ENDS BUFHSV24RQ
****Sub-Circuit for BUFHSV24RT, Wed Dec  8 16:10:26 CST 2010****
.SUBCKT BUFHSV24RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=6.48u L=60.00n
MM3 net11 I VDD VNW P12LL W=2.16u L=60.00n
MM2 net11 I VSS VPW N12LL W=1.72u L=60.00n
MM1 Z net11 VSS VPW N12LL W=5.16u L=60.00n
.ENDS BUFHSV24RT
****Sub-Circuit for BUFHSV2RQ, Thu May 19 13:57:40 CST 2011****
.SUBCKT BUFHSV2RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=430.00n L=60.00n
MM2 net7 I VSS VPW N12LL W=180.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=200.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=540.00n L=60.00n
.ENDS BUFHSV2RQ
****Sub-Circuit for BUFHSV2RT, Thu May 19 13:57:40 CST 2011****
.SUBCKT BUFHSV2RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=540.00n L=60.00n
MM3 net11 I VDD VNW P12LL W=200.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=180.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=430.00n L=60.00n
.ENDS BUFHSV2RT
****Sub-Circuit for BUFHSV3, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV3 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=260.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=650.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=390.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=980.00n L=60.00n
.ENDS BUFHSV3
****Sub-Circuit for BUFHSV32, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV32 I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=8.64u L=60.00n
MM3 net11 I VDD VNW P12LL W=4.32u L=60.00n
MM2 net11 I VSS VPW N12LL W=3.44u L=60.00n
MM1 Z net11 VSS VPW N12LL W=6.88u L=60.00n
.ENDS BUFHSV32
****Sub-Circuit for BUFHSV32RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV32RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=6.88u L=60.00n
MM2 net7 I VSS VPW N12LL W=860.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=1.08u L=60.00n
MM0 Z net7 VDD VNW P12LL W=8.64u L=60.00n
.ENDS BUFHSV32RO
****Sub-Circuit for BUFHSV32RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV32RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=6.88u L=60.00n
MM2 net7 I VSS VPW N12LL W=1.72u L=60.00n
MM3 net7 I VDD VNW P12LL W=2.16u L=60.00n
MM0 Z net7 VDD VNW P12LL W=8.64u L=60.00n
.ENDS BUFHSV32RQ
****Sub-Circuit for BUFHSV32RT, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV32RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=8.64u L=60.00n
MM3 net11 I VDD VNW P12LL W=2.88u L=60.00n
MM2 net11 I VSS VPW N12LL W=2.29u L=60.00n
MM1 Z net11 VSS VPW N12LL W=6.88u L=60.00n
.ENDS BUFHSV32RT
****Sub-Circuit for BUFHSV3RQ, Thu May 19 13:57:40 CST 2011****
.SUBCKT BUFHSV3RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=650.00n L=60.00n
MM2 net7 I VSS VPW N12LL W=180.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=200.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=810.00n L=60.00n
.ENDS BUFHSV3RQ
****Sub-Circuit for BUFHSV3RT, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV3RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=810.00n L=60.00n
MM3 net11 I VDD VNW P12LL W=270.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=220.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=650.00n L=60.00n
.ENDS BUFHSV3RT
****Sub-Circuit for BUFHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV4 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=340.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=860.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=520.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=1.3u L=60.00n
.ENDS BUFHSV4
****Sub-Circuit for BUFHSV40, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV40 I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=10.8u L=60.00n
MM3 net11 I VDD VNW P12LL W=5.4u L=60.00n
MM2 net11 I VSS VPW N12LL W=4.3u L=60.00n
MM1 Z net11 VSS VPW N12LL W=8.6u L=60.00n
.ENDS BUFHSV40
****Sub-Circuit for BUFHSV40RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV40RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=8.6u L=60.00n
MM2 net7 I VSS VPW N12LL W=1.07u L=60.00n
MM3 net7 I VDD VNW P12LL W=1.34u L=60.00n
MM0 Z net7 VDD VNW P12LL W=10.8u L=60.00n
.ENDS BUFHSV40RO
****Sub-Circuit for BUFHSV40RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV40RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=8.6u L=60.00n
MM2 net7 I VSS VPW N12LL W=2.15u L=60.00n
MM3 net7 I VDD VNW P12LL W=2.7u L=60.00n
MM0 Z net7 VDD VNW P12LL W=10.8u L=60.00n
.ENDS BUFHSV40RQ
****Sub-Circuit for BUFHSV40RT, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV40RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=10.8u L=60.00n
MM3 net11 I VDD VNW P12LL W=3.6u L=60.00n
MM2 net11 I VSS VPW N12LL W=2.87u L=60.00n
MM1 Z net11 VSS VPW N12LL W=8.6u L=60.00n
.ENDS BUFHSV40RT
****Sub-Circuit for BUFHSV48, Thu Feb 17 14:51:05 CST 2011****
.SUBCKT BUFHSV48 I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=12.96u L=60.00n
MM3 net11 I VDD VNW P12LL W=6.48u L=60.00n
MM2 net11 I VSS VPW N12LL W=5.16u L=60.00n
MM1 Z net11 VSS VPW N12LL W=10.32u L=60.00n
.ENDS BUFHSV48
****Sub-Circuit for BUFHSV48RO, Thu Feb 17 14:51:05 CST 2011****
.SUBCKT BUFHSV48RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=10.32u L=60.00n
MM2 net7 I VSS VPW N12LL W=1.29u L=60.00n
MM3 net7 I VDD VNW P12LL W=1.62u L=60.00n
MM0 Z net7 VDD VNW P12LL W=12.96u L=60.00n
.ENDS BUFHSV48RO
****Sub-Circuit for BUFHSV48RQ, Thu Feb 17 14:51:05 CST 2011****
.SUBCKT BUFHSV48RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=10.32u L=60.00n
MM2 net7 I VSS VPW N12LL W=2.58u L=60.00n
MM3 net7 I VDD VNW P12LL W=3.24u L=60.00n
MM0 Z net7 VDD VNW P12LL W=12.96u L=60.00n
.ENDS BUFHSV48RQ
****Sub-Circuit for BUFHSV4RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV4RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=860.00n L=60.00n
MM2 net7 I VSS VPW N12LL W=210.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=270.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=1.08u L=60.00n
.ENDS BUFHSV4RQ
****Sub-Circuit for BUFHSV4RT, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV4RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=1.08u L=60.00n
MM3 net11 I VDD VNW P12LL W=360.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=290.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=860.00n L=60.00n
.ENDS BUFHSV4RT
****Sub-Circuit for BUFHSV6, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV6 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=430.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=1.29u L=60.00n
MM1 net13 I VDD VNW P12LL W=650.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=1.95u L=60.00n
.ENDS BUFHSV6
****Sub-Circuit for BUFHSV6RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV6RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=1.29u L=60.00n
MM2 net7 I VSS VPW N12LL W=320.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=400.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=1.62u L=60.00n
.ENDS BUFHSV6RQ
****Sub-Circuit for BUFHSV6RT, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV6RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=1.62u L=60.00n
MM3 net11 I VDD VNW P12LL W=540.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=430.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=1.29u L=60.00n
.ENDS BUFHSV6RT
****Sub-Circuit for BUFHSV8, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT BUFHSV8 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=680.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=1.72u L=60.00n
MM1 net13 I VDD VNW P12LL W=1.02u L=60.00n
MM3 Z net13 VDD VNW P12LL W=2.6u L=60.00n
.ENDS BUFHSV8
****Sub-Circuit for BUFHSV8RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV8RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=1.72u L=60.00n
MM2 net7 I VSS VPW N12LL W=210.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=270.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=2.16u L=60.00n
.ENDS BUFHSV8RO
****Sub-Circuit for BUFHSV8RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV8RQ I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=1.72u L=60.00n
MM2 net7 I VSS VPW N12LL W=430.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=540.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=2.16u L=60.00n
.ENDS BUFHSV8RQ
****Sub-Circuit for BUFHSV8RT, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT BUFHSV8RT I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=2.16u L=60.00n
MM3 net11 I VDD VNW P12LL W=720.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=570.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=1.72u L=60.00n
.ENDS BUFHSV8RT
****Sub-Circuit for CKMUX2HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CKMUX2HSV0 I0 I1 S Z VDD VSS
MM47 net41 S net27 VPW N12LL W=180.00n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=180.00n L=60.00n
MM31 net43 S VSS VPW N12LL W=180.00n L=60.00n
MM30 Z net27 VSS VPW N12LL W=200.00n L=60.00n
MM27 net41 I1 VSS VPW N12LL W=180.00n L=60.00n
MM36 net39 net43 net27 VPW N12LL W=180.00n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=350.00n L=60.00n
MM48 net41 net43 net27 VNW P12LL W=350.00n L=60.00n
MM32 net43 S VDD VNW P12LL W=350.00n L=60.00n
MM29 Z net27 VDD VNW P12LL W=400.00n L=60.00n
MM28 net41 I1 VDD VNW P12LL W=350.00n L=60.00n
MM39 net39 S net27 VNW P12LL W=350.00n L=60.00n
.ENDS CKMUX2HSV0
****Sub-Circuit for CKMUX2HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CKMUX2HSV1 I0 I1 S Z VDD VSS
MM47 net41 S net27 VPW N12LL W=200.00n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=200.00n L=60.00n
MM31 net43 S VSS VPW N12LL W=200.00n L=60.00n
MM30 Z net27 VSS VPW N12LL W=260.00n L=60.00n
MM27 net41 I1 VSS VPW N12LL W=200.00n L=60.00n
MM36 net39 net43 net27 VPW N12LL W=200.00n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=360.00n L=60.00n
MM48 net41 net43 net27 VNW P12LL W=330.00n L=60.00n
MM32 net43 S VDD VNW P12LL W=330.00n L=60.00n
MM29 Z net27 VDD VNW P12LL W=450.00n L=60.00n
MM28 net41 I1 VDD VNW P12LL W=360.00n L=60.00n
MM39 net39 S net27 VNW P12LL W=330.00n L=60.00n
.ENDS CKMUX2HSV1
****Sub-Circuit for CKMUX2HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CKMUX2HSV2 I0 I1 S Z VDD VSS
MM47 net41 S net27 VPW N12LL W=260.00n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=260.00n L=60.00n
MM31 net43 S VSS VPW N12LL W=280.00n L=60.00n
MM30 Z net27 VSS VPW N12LL W=360.00n L=60.00n
MM27 net41 I1 VSS VPW N12LL W=260.00n L=60.00n
MM36 net39 net43 net27 VPW N12LL W=260.00n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=450.00n L=60.00n
MM48 net41 net43 net27 VNW P12LL W=450.00n L=60.00n
MM32 net43 S VDD VNW P12LL W=450.00n L=60.00n
MM29 Z net27 VDD VNW P12LL W=650.00n L=60.00n
MM28 net41 I1 VDD VNW P12LL W=450.00n L=60.00n
MM39 net39 S net27 VNW P12LL W=450.00n L=60.00n
.ENDS CKMUX2HSV2
****Sub-Circuit for CKMUX2HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CKMUX2HSV4 I0 I1 S Z VDD VSS
MM47 net41 S net27 VPW N12LL W=350.00n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=360.00n L=60.00n
MM31 net43 S VSS VPW N12LL W=430.00n L=60.00n
MM30 Z net27 VSS VPW N12LL W=710.00n L=60.00n
MM27 net41 I1 VSS VPW N12LL W=350.00n L=60.00n
MM36 net39 net43 net27 VPW N12LL W=360.00n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=650.00n L=60.00n
MM48 net41 net43 net27 VNW P12LL W=650.00n L=60.00n
MM32 net43 S VDD VNW P12LL W=650.00n L=60.00n
MM29 Z net27 VDD VNW P12LL W=1.3u L=60.00n
MM28 net41 I1 VDD VNW P12LL W=650.00n L=60.00n
MM39 net39 S net27 VNW P12LL W=650.00n L=60.00n
.ENDS CKMUX2HSV4
****Sub-Circuit for CLKAND2HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKAND2HSV0 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=280.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=280.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=330.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=280.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=280.00n L=60.00n
.ENDS CLKAND2HSV0
****Sub-Circuit for CLKAND2HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKAND2HSV1 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=300.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=260.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=300.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=450.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS CLKAND2HSV1
****Sub-Circuit for CLKAND2HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKAND2HSV2 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=410.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=360.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=410.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=650.00n L=60.00n
MM0 net11 A2 VDD VNW P12LL W=420.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=420.00n L=60.00n
.ENDS CLKAND2HSV2
****Sub-Circuit for CLKAND2HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKAND2HSV4 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=640.00n L=60.00n
MM2 Z net11 VSS VPW N12LL W=710.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=640.00n L=60.00n
MM3 Z net11 VDD VNW P12LL W=1.3u L=60.00n
MM0 net11 A2 VDD VNW P12LL W=640.00n L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=640.00n L=60.00n
.ENDS CLKAND2HSV4
****Sub-Circuit for CLKAND2HSV8, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKAND2HSV8 A1 A2 Z VDD VSS
MM1 net11 A1 net18 VPW N12LL W=1.2u L=60.00n
MM2 Z net11 VSS VPW N12LL W=1.3u L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=1.2u L=60.00n
MM3 Z net11 VDD VNW P12LL W=2.6u L=60.00n
MM0 net11 A2 VDD VNW P12LL W=1.28u L=60.00n
MMP1 net11 A1 VDD VNW P12LL W=1.28u L=60.00n
.ENDS CLKAND2HSV8
****Sub-Circuit for CLKBUFHSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV0 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=200.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=330.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=330.0n L=60.00n
.ENDS CLKBUFHSV0
****Sub-Circuit for CLKBUFHSV0P5, Thu May 19 13:57:40 CST 2011****
.SUBCKT CLKBUFHSV0P5 I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=220.00n L=60.00n
MM2 net7 I VSS VPW N12LL W=180.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=360.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=450.00n L=60.00n
.ENDS CLKBUFHSV0P5
****Sub-Circuit for CLKBUFHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV1 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=260.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=350.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=450.0n L=60.00n
.ENDS CLKBUFHSV1
****Sub-Circuit for CLKBUFHSV12, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV12 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=640.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=1.86u L=60.00n
MM1 net13 I VDD VNW P12LL W=1.3u L=60.00n
MM3 Z net13 VDD VNW P12LL W=3.9u L=60.00n
.ENDS CLKBUFHSV12
****Sub-Circuit for CLKBUFHSV12RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV12RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=1.92u L=60.00n
MM2 net7 I VSS VPW N12LL W=240.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=480.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=3.9u L=60.00n
.ENDS CLKBUFHSV12RO
****Sub-Circuit for CLKBUFHSV12RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV12RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=3.9u L=60.00n
MM3 net11 I VDD VNW P12LL W=970.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=480.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=1.92u L=60.00n
.ENDS CLKBUFHSV12RQ
****Sub-Circuit for CLKBUFHSV16, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV16 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=840.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=2.56u L=60.00n
MM1 net13 I VDD VNW P12LL W=1.74u L=60.00n
MM3 Z net13 VDD VNW P12LL W=5.2u L=60.00n
.ENDS CLKBUFHSV16
****Sub-Circuit for CLKBUFHSV16RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV16RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=2.56u L=60.00n
MM2 net7 I VSS VPW N12LL W=320.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=650.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=5.2u L=60.00n
.ENDS CLKBUFHSV16RO
****Sub-Circuit for CLKBUFHSV16RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV16RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=5.2u L=60.00n
MM3 net11 I VDD VNW P12LL W=1.3u L=60.00n
MM2 net11 I VSS VPW N12LL W=640.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=2.56u L=60.00n
.ENDS CLKBUFHSV16RQ
****Sub-Circuit for CLKBUFHSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV2 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=360.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=340.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=640.0n L=60.00n
.ENDS CLKBUFHSV2
****Sub-Circuit for CLKBUFHSV20, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV20 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=1.08u L=60.00n
MM2 Z net13 VSS VPW N12LL W=3.25u L=60.00n
MM1 net13 I VDD VNW P12LL W=2.28u L=60.00n
MM3 Z net13 VDD VNW P12LL W=6.5u L=60.00n
.ENDS CLKBUFHSV20
****Sub-Circuit for CLKBUFHSV20RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV20RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=3.2u L=60.00n
MM2 net7 I VSS VPW N12LL W=400.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=810.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=6.5u L=60.00n
.ENDS CLKBUFHSV20RO
****Sub-Circuit for CLKBUFHSV20RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV20RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=6.5u L=60.00n
MM3 net11 I VDD VNW P12LL W=1.62u L=60.00n
MM2 net11 I VSS VPW N12LL W=800.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=3.2u L=60.00n
.ENDS CLKBUFHSV20RQ
****Sub-Circuit for CLKBUFHSV24, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV24 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=1.24u L=60.00n
MM2 Z net13 VSS VPW N12LL W=3.84u L=60.00n
MM1 net13 I VDD VNW P12LL W=2.6u L=60.00n
MM3 Z net13 VDD VNW P12LL W=7.8u L=60.00n
.ENDS CLKBUFHSV24
****Sub-Circuit for CLKBUFHSV24RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV24RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=3.84u L=60.00n
MM2 net7 I VSS VPW N12LL W=480.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=970.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=7.8u L=60.00n
.ENDS CLKBUFHSV24RO
****Sub-Circuit for CLKBUFHSV24RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV24RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=7.8u L=60.00n
MM3 net11 I VDD VNW P12LL W=1.95u L=60.00n
MM2 net11 I VSS VPW N12LL W=960.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=3.84u L=60.00n
.ENDS CLKBUFHSV24RQ
****Sub-Circuit for CLKBUFHSV2RQ, Thu May 19 13:57:40 CST 2011****
.SUBCKT CLKBUFHSV2RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=650.00n L=60.00n
MM3 net11 I VDD VNW P12LL W=360.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=180.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=320.00n L=60.00n
.ENDS CLKBUFHSV2RQ
****Sub-Circuit for CLKBUFHSV3, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV3 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=270.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=530.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=500.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=980.00n L=60.00n
.ENDS CLKBUFHSV3
****Sub-Circuit for CLKBUFHSV32, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV32 I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=5.12u L=60.00n
MM2 net7 I VSS VPW N12LL W=2.56u L=60.00n
MM3 net7 I VDD VNW P12LL W=5.2u L=60.00n
MM0 Z net7 VDD VNW P12LL W=10.4u L=60.00n
.ENDS CLKBUFHSV32
****Sub-Circuit for CLKBUFHSV32RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV32RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=5.12u L=60.00n
MM2 net7 I VSS VPW N12LL W=640.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=1.3u L=60.00n
MM0 Z net7 VDD VNW P12LL W=10.4u L=60.00n
.ENDS CLKBUFHSV32RO
****Sub-Circuit for CLKBUFHSV32RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV32RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=10.4u L=60.00n
MM3 net11 I VDD VNW P12LL W=2.6u L=60.00n
MM2 net11 I VSS VPW N12LL W=1.28u L=60.00n
MM1 Z net11 VSS VPW N12LL W=5.12u L=60.00n
.ENDS CLKBUFHSV32RQ
****Sub-Circuit for CLKBUFHSV3RQ, Thu May 19 13:57:40 CST 2011****
.SUBCKT CLKBUFHSV3RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=970.00n L=60.00n
MM3 net11 I VDD VNW P12LL W=360.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=180.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=480.00n L=60.00n
.ENDS CLKBUFHSV3RQ
****Sub-Circuit for CLKBUFHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV4 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=360.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=710.00n L=60.00n
MM1 net13 I VDD VNW P12LL W=630.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=1.3u L=60.00n
.ENDS CLKBUFHSV4
****Sub-Circuit for CLKBUFHSV40, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV40 I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=6.4u L=60.00n
MM2 net7 I VSS VPW N12LL W=3.2u L=60.00n
MM3 net7 I VDD VNW P12LL W=6.5u L=60.00n
MM0 Z net7 VDD VNW P12LL W=13.00u L=60.00n
.ENDS CLKBUFHSV40
****Sub-Circuit for CLKBUFHSV40RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV40RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=6.4u L=60.00n
MM2 net7 I VSS VPW N12LL W=800.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=1.62u L=60.00n
MM0 Z net7 VDD VNW P12LL W=13.00u L=60.00n
.ENDS CLKBUFHSV40RO
****Sub-Circuit for CLKBUFHSV40RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV40RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=13.00u L=60.00n
MM3 net11 I VDD VNW P12LL W=3.25u L=60.00n
MM2 net11 I VSS VPW N12LL W=1.6u L=60.00n
MM1 Z net11 VSS VPW N12LL W=6.4u L=60.00n
.ENDS CLKBUFHSV40RQ
****Sub-Circuit for CLKBUFHSV48, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV48 I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=7.68u L=60.00n
MM2 net7 I VSS VPW N12LL W=3.84u L=60.00n
MM3 net7 I VDD VNW P12LL W=7.8u L=60.00n
MM0 Z net7 VDD VNW P12LL W=15.6u L=60.00n
.ENDS CLKBUFHSV48
****Sub-Circuit for CLKBUFHSV48RO, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV48RO I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=7.68u L=60.00n
MM2 net7 I VSS VPW N12LL W=960.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=1.95u L=60.00n
MM0 Z net7 VDD VNW P12LL W=15.6u L=60.00n
.ENDS CLKBUFHSV48RO
****Sub-Circuit for CLKBUFHSV48RQ, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV48RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=15.6u L=60.00n
MM3 net11 I VDD VNW P12LL W=3.9u L=60.00n
MM2 net11 I VSS VPW N12LL W=1.92u L=60.00n
MM1 Z net11 VSS VPW N12LL W=7.68u L=60.00n
.ENDS CLKBUFHSV48RQ
****Sub-Circuit for CLKBUFHSV4RQ, Thu May 19 13:57:40 CST 2011****
.SUBCKT CLKBUFHSV4RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=1.3u L=60.00n
MM3 net11 I VDD VNW P12LL W=360.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=180.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=640.00n L=60.00n
.ENDS CLKBUFHSV4RQ
****Sub-Circuit for CLKBUFHSV5, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKBUFHSV5 I Z VDD VSS
MM1 Z net7 VSS VPW N12LL W=800.00n L=60.00n
MM2 net7 I VSS VPW N12LL W=400.00n L=60.00n
MM3 net7 I VDD VNW P12LL W=810.00n L=60.00n
MM0 Z net7 VDD VNW P12LL W=1.62u L=60.00n
.ENDS CLKBUFHSV5
****Sub-Circuit for CLKBUFHSV5RQ, Thu Feb 17 17:27:06 CST 2011****
.SUBCKT CLKBUFHSV5RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=1.62u L=60.00n
MM3 net11 I VDD VNW P12LL W=400.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=200.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=800.00n L=60.00n
.ENDS CLKBUFHSV5RQ
****Sub-Circuit for CLKBUFHSV6, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV6 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=350.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=1.02u L=60.00n
MM1 net13 I VDD VNW P12LL W=650.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=1.95u L=60.00n
.ENDS CLKBUFHSV6
****Sub-Circuit for CLKBUFHSV6RQ, Thu Feb 17 17:27:06 CST 2011****
.SUBCKT CLKBUFHSV6RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=1.95u L=60.00n
MM3 net11 I VDD VNW P12LL W=480.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=240.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=960.00n L=60.00n
.ENDS CLKBUFHSV6RQ
****Sub-Circuit for CLKBUFHSV8, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKBUFHSV8 I Z VDD VSS
MM0 net13 I VSS VPW N12LL W=430.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=1.3u L=60.00n
MM1 net13 I VDD VNW P12LL W=850.00n L=60.00n
MM3 Z net13 VDD VNW P12LL W=2.6u L=60.00n
.ENDS CLKBUFHSV8
****Sub-Circuit for CLKBUFHSV8RO, Thu May 19 13:57:40 CST 2011****
.SUBCKT CLKBUFHSV8RO I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=2.6u L=60.00n
MM3 net11 I VDD VNW P12LL W=360.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=180.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=1.28u L=60.00n
.ENDS CLKBUFHSV8RO
****Sub-Circuit for CLKBUFHSV8RQ, Thu Feb 17 17:27:06 CST 2011****
.SUBCKT CLKBUFHSV8RQ I Z VDD VSS
MM0 Z net11 VDD VNW P12LL W=2.6u L=60.00n
MM3 net11 I VDD VNW P12LL W=650.00n L=60.00n
MM2 net11 I VSS VPW N12LL W=320.00n L=60.00n
MM1 Z net11 VSS VPW N12LL W=1.28u L=60.00n
.ENDS CLKBUFHSV8RQ
****Sub-Circuit for CLKLAHAQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHAQHSV1 CK E Q TE VDD VSS
MM51 s c VSS VPW N12LL W=200.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=200.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=260.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=200.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM0 ten TE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=220.00n L=60.00n
MM22 Q s VSS VPW N12LL W=320.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=260.00n L=60.00n
MM45 s c nt21 VNW P12LL W=540.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=540.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=500.00n L=60.00n
MM1 ten TE VDD VNW P12LL W=300.00n L=60.00n
MM54 nt21 pm VDD VNW P12LL W=540.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=330.00n L=60.00n
MM21 Q s VDD VNW P12LL W=460.00n L=60.00n
MM39 pm cn nt11 VNW P12LL W=500.00n L=60.00n
.ENDS CLKLAHAQHSV1
****Sub-Circuit for CLKLAHAQHSV2, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHAQHSV2 CK E Q TE VDD VSS
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM39 pm cn nt11 VNW P12LL W=440.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=250.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=540.00n L=60.00n
MM45 s c nt21 VNW P12LL W=440.00n L=60.00n
MM54 nt21 pm VDD VNW P12LL W=540.00n L=60.00n
MM21 Q s VDD VNW P12LL W=540.00n L=60.00n
MM1 ten TE VDD VNW P12LL W=340.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=440.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=350.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=350.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=350.00n L=60.00n
MM51 s c VSS VPW N12LL W=350.00n L=60.00n
MM22 Q s VSS VPW N12LL W=430.00n L=60.00n
MM0 ten TE VSS VPW N12LL W=270.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=350.00n L=60.00n
.ENDS CLKLAHAQHSV2
****Sub-Circuit for CLKLAHAQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHAQHSV4 CK E Q TE VDD VSS
MM51 s c VSS VPW N12LL W=300.00n L=60.00n
MM49 m pm VSS VPW N12LL W=300.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=300.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=260.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=300.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM0 ten TE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=220.00n L=60.00n
MM22 Q s VSS VPW N12LL W=860.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=260.00n L=60.00n
MM45 s c nt21 VNW P12LL W=600.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=600.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=600.00n L=60.00n
MM1 ten TE VDD VNW P12LL W=300.00n L=60.00n
MM54 nt21 pm VDD VNW P12LL W=590.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=330.00n L=60.00n
MM21 Q s VDD VNW P12LL W=1.2u L=60.00n
MM39 pm cn nt11 VNW P12LL W=600.00n L=60.00n
.ENDS CLKLAHAQHSV4
****Sub-Circuit for CLKLAHAQHSV8, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHAQHSV8 CK E Q TE VDD VSS
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM39 pm cn nt11 VNW P12LL W=540.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM14 nt13 c pm VNW P12LL W=250.00n L=60.00n
MM46 nt21 ten VDD VNW P12LL W=1.3u L=60.00n
MM45 s c nt21 VNW P12LL W=1.08u L=60.00n
MM54 nt21 pm VDD VNW P12LL W=1.3u L=60.00n
MM21 Q s VDD VNW P12LL W=2.16u L=60.00n
MM1 ten TE VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=540.00n L=60.00n
MM51 s c VSS VPW N12LL W=860.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=430.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 cn pm VPW N12LL W=200.00n L=60.00n
MM43 s pm nt22 VPW N12LL W=860.00n L=60.00n
MM44 nt22 ten VSS VPW N12LL W=860.00n L=60.00n
MM22 Q s VSS VPW N12LL W=1.72u L=60.00n
MM0 ten TE VSS VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM36 pm c nt12 VPW N12LL W=430.00n L=60.00n
.ENDS CLKLAHAQHSV8
****Sub-Circuit for CLKLAHQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHQHSV1 CK E Q TE VDD VSS
MM51 hnet12 TE VSS VPW N12LL W=300.00n L=60.00n
MM49 m pm VSS VPW N12LL W=300.00n L=60.00n
MM43 s pm VSS VPW N12LL W=230.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=300.00n L=60.00n
MM44 s c VSS VPW N12LL W=230.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=270n L=60.00n
MM27 cn CK VSS VPW N12LL W=220n L=60.00n
MM22 Q s VSS VPW N12LL W=340.00n L=60.00n
MM36 pm c hnet12 VPW N12LL W=300.00n L=60.00n
MM45 s c hnet31 VNW P12LL W=550.00n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=550.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=590.0n L=60.00n
MM54 hnet13 TE VDD VNW P12LL W=590.0n L=60.00n
MM14 hnet21 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400n L=60.00n
MM28 cn CK VDD VNW P12LL W=330n L=60.00n
MM21 Q s VDD VNW P12LL W=440.00n L=60.00n
MM39 pm cn hnet11 VNW P12LL W=590.0n L=60.00n
.ENDS CLKLAHQHSV1
****Sub-Circuit for CLKLAHQHSV2, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHQHSV2 CK E Q TE VDD VSS
MM22 Q s VSS VPW N12LL W=430.00n L=60.00n
MM44 s c VSS VPW N12LL W=270.00n L=60.00n
MM43 s pm VSS VPW N12LL W=270.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM51 hnet12 TE VSS VPW N12LL W=350.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=350.00n L=60.00n
MM36 pm c hnet12 VPW N12LL W=350.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270n L=60.00n
MM30 c cn VSS VPW N12LL W=350n L=60.00n
MM21 Q s VDD VNW P12LL W=540.00n L=60.00n
MM45 s c hnet31 VNW P12LL W=500.00n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=500.00n L=60.00n
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM14 hnet21 c pm VNW P12LL W=250.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=250.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=440.0n L=60.00n
MM39 pm cn hnet11 VNW P12LL W=440.0n L=60.00n
MM54 hnet13 TE VDD VNW P12LL W=440.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=340n L=60.00n
MM29 c cn VDD VNW P12LL W=440n L=60.00n
.ENDS CLKLAHQHSV2
****Sub-Circuit for CLKLAHQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLAHQHSV4 CK E Q TE VDD VSS
MM51 hnet12 TE VSS VPW N12LL W=340.00n L=60.00n
MM49 m pm VSS VPW N12LL W=400.00n L=60.00n
MM43 s pm VSS VPW N12LL W=280.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=340.00n L=60.00n
MM44 s c VSS VPW N12LL W=280.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=270n L=60.00n
MM27 cn CK VSS VPW N12LL W=220n L=60.00n
MM22 Q s VSS VPW N12LL W=860n L=60.00n
MM36 pm c hnet12 VPW N12LL W=340.00n L=60.00n
MM45 s c hnet31 VNW P12LL W=640.00n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=640.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=650.0n L=60.00n
MM54 hnet13 TE VDD VNW P12LL W=650.0n L=60.00n
MM14 hnet21 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400n L=60.00n
MM28 cn CK VDD VNW P12LL W=330n L=60.00n
MM21 Q s VDD VNW P12LL W=1.2u L=60.00n
MM39 pm cn hnet11 VNW P12LL W=650.0n L=60.00n
.ENDS CLKLAHQHSV4
****Sub-Circuit for CLKLAHQHSV8, Wed Apr  6 20:02:58 CST 2011****
.SUBCKT CLKLAHQHSV8 CK E Q TE VDD VSS
MM22 Q s VSS VPW N12LL W=1.72u L=60.00n
MM44 s c VSS VPW N12LL W=580.00n L=60.00n
MM43 s pm VSS VPW N12LL W=580.00n L=60.00n
MM11 VSS m hnet22 VPW N12LL W=200.00n L=60.00n
MM12 hnet22 cn pm VPW N12LL W=200.00n L=60.00n
MM51 hnet12 TE VSS VPW N12LL W=430.00n L=60.00n
MM52 hnet12 E VSS VPW N12LL W=430.00n L=60.00n
MM36 pm c hnet12 VPW N12LL W=430.00n L=60.00n
MM49 m pm VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270n L=60.00n
MM30 c cn VSS VPW N12LL W=430n L=60.00n
MM21 Q s VDD VNW P12LL W=2.16u L=60.00n
MM45 s c hnet31 VNW P12LL W=1080n L=60.00n
MM46 hnet31 pm VDD VNW P12LL W=1080n L=60.00n
MM50 m pm VDD VNW P12LL W=250.00n L=60.00n
MM14 hnet21 c pm VNW P12LL W=250.00n L=60.00n
MM13 VDD m hnet21 VNW P12LL W=250.00n L=60.00n
MM53 hnet11 E hnet13 VNW P12LL W=540.00n L=60.00n
MM39 pm cn hnet11 VNW P12LL W=540.00n L=60.00n
MM54 hnet13 TE VDD VNW P12LL W=540.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340n L=60.00n
MM29 c cn VDD VNW P12LL W=540n L=60.00n
.ENDS CLKLAHQHSV8
****Sub-Circuit for CLKLANAQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANAQHSV1 CK E Q TE VDD VSS
MM51 nt22 TE VSS VPW N12LL W=300.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c nt22 VPW N12LL W=300.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=260.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=300.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM22 Q s VSS VPW N12LL W=290.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=260.00n L=60.00n
MM45 s m nt21 VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=400.00n L=60.00n
MM54 nt21 TE VDD VNW P12LL W=300.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=360.00n L=60.00n
MM21 Q s VDD VNW P12LL W=460.00n L=60.00n
MM39 pm c nt11 VNW P12LL W=400.00n L=60.00n
.ENDS CLKLANAQHSV1
****Sub-Circuit for CLKLANAQHSV2, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT CLKLANAQHSV2 CK E Q TE VDD VSS
MM39 pm c nt11 VNW P12LL W=440.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=440.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=250.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM50 m pm VDD VNW P12LL W=350.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM29 c cn VDD VNW P12LL W=430.00n L=60.00n
MM54 nt21 TE VDD VNW P12LL W=350.00n L=60.00n
MM45 s m nt21 VNW P12LL W=350.00n L=60.00n
MM46 s c VDD VNW P12LL W=350.00n L=60.00n
MM21 Q s VDD VNW P12LL W=540.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=350.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=350.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM49 m pm VSS VPW N12LL W=280.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=350.00n L=60.00n
MM51 nt22 TE VSS VPW N12LL W=350.00n L=60.00n
MM43 s c nt22 VPW N12LL W=350.00n L=60.00n
MM22 Q s VSS VPW N12LL W=430.00n L=60.00n
.ENDS CLKLANAQHSV2
****Sub-Circuit for CLKLANAQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANAQHSV4 CK E Q TE VDD VSS
MM51 nt22 TE VSS VPW N12LL W=430.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c nt22 VPW N12LL W=430.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=320.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=270.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM22 Q s VSS VPW N12LL W=800.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=320.00n L=60.00n
MM45 s m nt21 VNW P12LL W=430.00n L=60.00n
MM46 s c VDD VNW P12LL W=430.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=450.00n L=60.00n
MM54 nt21 TE VDD VNW P12LL W=430.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=360.00n L=60.00n
MM21 Q s VDD VNW P12LL W=1.3u L=60.00n
MM39 pm c nt11 VNW P12LL W=450.00n L=60.00n
.ENDS CLKLANAQHSV4
****Sub-Circuit for CLKLANAQHSV8, Fri Jan 28 15:34:45 CST 2011****
.SUBCKT CLKLANAQHSV8 CK E Q TE VDD VSS
MM21 Q s VDD VNW P12LL W=2.16u L=60.00n
MM46 s c VDD VNW P12LL W=860.00n L=60.00n
MM45 s m nt21 VNW P12LL W=860.00n L=60.00n
MM54 nt21 TE VDD VNW P12LL W=860.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=340.00n L=60.00n
MM50 m pm VDD VNW P12LL W=540.00n L=60.00n
MM13 VDD m nt13 VNW P12LL W=250.00n L=60.00n
MM14 nt13 cn pm VNW P12LL W=250.00n L=60.00n
MM53 nt11 E VDD VNW P12LL W=540.00n L=60.00n
MM39 pm c nt11 VNW P12LL W=540.00n L=60.00n
MM43 s c nt22 VPW N12LL W=860.00n L=60.00n
MM22 Q s VSS VPW N12LL W=1.72u L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM51 nt22 TE VSS VPW N12LL W=860.00n L=60.00n
MM44 nt22 m VSS VPW N12LL W=860.00n L=60.00n
MM12 nt14 c pm VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=270.00n L=60.00n
MM49 m pm VSS VPW N12LL W=430.00n L=60.00n
MM52 nt12 E VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m nt14 VPW N12LL W=200.00n L=60.00n
MM36 pm cn nt12 VPW N12LL W=430.00n L=60.00n
.ENDS CLKLANAQHSV8
****Sub-Circuit for CLKLANQHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV1 CK E Q TE VDD VSS
MM51 hnet22 TE VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 Q s VSS VPW N12LL W=290.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 Q s VDD VNW P12LL W=460.00n L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV1
****Sub-Circuit for CLKLANQHSV12, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV12 CK E Q TE VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 TE VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=860.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 Q pq VSS VPW N12LL W=2.46u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.2u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 Q pq VDD VNW P12LL W=3.9u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV12
****Sub-Circuit for CLKLANQHSV16, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV16 CK E Q TE VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 TE VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=860.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 Q pq VSS VPW N12LL W=3.42u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.2u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 Q pq VDD VNW P12LL W=5.2u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV16
****Sub-Circuit for CLKLANQHSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV2 CK E Q TE VDD VSS
MM51 hnet22 TE VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 Q s VSS VPW N12LL W=420.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 Q s VDD VNW P12LL W=650.00n L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV2
****Sub-Circuit for CLKLANQHSV20, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV20 CK E Q TE VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 TE VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=1.29u L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 Q pq VSS VPW N12LL W=4.2u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.74u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 Q pq VDD VNW P12LL W=6.5u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV20
****Sub-Circuit for CLKLANQHSV24, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV24 CK E Q TE VDD VSS
MM55 ps s VSS VPW N12LL W=420.00n L=60.00n
MM51 hnet22 TE VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=280.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=280.00n L=60.00n
MM57 pq ps VSS VPW N12LL W=1.29u L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 Q pq VSS VPW N12LL W=5.16u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM56 ps s VDD VNW P12LL W=650.00n L=60.00n
MM45 s m VDD VNW P12LL W=300.00n L=60.00n
MM46 s c VDD VNW P12LL W=300.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=400.0n L=60.00n
MM58 pq ps VDD VNW P12LL W=1.74u L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 Q pq VDD VNW P12LL W=7.8u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV24
****Sub-Circuit for CLKLANQHSV3, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV3 CK E Q TE VDD VSS
MM51 hnet22 TE VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=360.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=360.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 Q s VSS VPW N12LL W=620.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=400.00n L=60.00n
MM46 s c VDD VNW P12LL W=400.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 Q s VDD VNW P12LL W=960.00n L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV3
****Sub-Circuit for CLKLANQHSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV4 CK E Q TE VDD VSS
MM51 hnet22 TE VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=260.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=430.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=260n L=60.00n
MM27 cn CK VSS VPW N12LL W=240n L=60.00n
MM22 Q s VSS VPW N12LL W=800.00n L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=500.00n L=60.00n
MM46 s c VDD VNW P12LL W=500.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=400n L=60.00n
MM28 cn CK VDD VNW P12LL W=360n L=60.00n
MM21 Q s VDD VNW P12LL W=1.3u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV4
****Sub-Circuit for CLKLANQHSV6, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV6 CK E Q TE VDD VSS
MM51 hnet22 TE VSS VPW N12LL W=340.00n L=60.00n
MM49 m pm VSS VPW N12LL W=380.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=430.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=340.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=430.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=360n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM22 Q s VSS VPW N12LL W=1.14u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=340.00n L=60.00n
MM45 s m VDD VNW P12LL W=440.00n L=60.00n
MM46 s c VDD VNW P12LL W=440.00n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=600.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=600.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540n L=60.00n
MM28 cn CK VDD VNW P12LL W=450n L=60.00n
MM21 Q s VDD VNW P12LL W=1.95u L=60.00n
MM39 pm c hnet24 VNW P12LL W=600.0n L=60.00n
.ENDS CLKLANQHSV6
****Sub-Circuit for CLKLANQHSV8, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKLANQHSV8 CK E Q TE VDD VSS
MM51 hnet22 TE VSS VPW N12LL W=320.00n L=60.00n
MM49 m pm VSS VPW N12LL W=360.00n L=60.00n
MM43 s c hnet36 VPW N12LL W=740.00n L=60.00n
MM52 hnet22 E VSS VPW N12LL W=320.00n L=60.00n
MM44 hnet36 m VSS VPW N12LL W=740.00n L=60.00n
MM11 VSS m hnet38 VPW N12LL W=200.00n L=60.00n
MM12 hnet38 c pm VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=360n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM22 Q s VSS VPW N12LL W=1.6u L=60.00n
MM36 pm cn hnet22 VPW N12LL W=320.00n L=60.00n
MM45 s m VDD VNW P12LL W=800.0n L=60.00n
MM46 s c VDD VNW P12LL W=800.0n L=60.00n
MM53 hnet24 E hnet26 VNW P12LL W=400.0n L=60.00n
MM54 hnet26 TE VDD VNW P12LL W=400.0n L=60.00n
MM14 hnet40 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m hnet40 VNW P12LL W=300.00n L=60.00n
MM50 m pm VDD VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=540n L=60.00n
MM28 cn CK VDD VNW P12LL W=450n L=60.00n
MM21 Q s VDD VNW P12LL W=2.6u L=60.00n
MM39 pm c hnet24 VNW P12LL W=400.0n L=60.00n
.ENDS CLKLANQHSV8
****Sub-Circuit for CLKNAND2HSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNAND2HSV0 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=300.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=300.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=330.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=330.00n L=60.00n
.ENDS CLKNAND2HSV0
****Sub-Circuit for CLKNAND2HSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNAND2HSV1 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=400.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=400.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=450.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=450.00n L=60.00n
.ENDS CLKNAND2HSV1
****Sub-Circuit for CLKNAND2HSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNAND2HSV2 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=540.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=540.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=650.00n L=60.00n
.ENDS CLKNAND2HSV2
****Sub-Circuit for CLKNAND2HSV3, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNAND2HSV3 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=740.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=740.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=980.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=980.00n L=60.00n
.ENDS CLKNAND2HSV3
****Sub-Circuit for CLKNAND2HSV4, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNAND2HSV4 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=1.00u L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=1.00u L=60.00n
MM0 ZN A2 VDD VNW P12LL W=1.3u L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=1.3u L=60.00n
.ENDS CLKNAND2HSV4
****Sub-Circuit for CLKNAND2HSV8, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNAND2HSV8 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=2.00u L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=2.00u L=60.00n
MM0 ZN A2 VDD VNW P12LL W=2.6u L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=2.6u L=60.00n
.ENDS CLKNAND2HSV8
****Sub-Circuit for CLKNHSV0, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNHSV0 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=200.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=330.0n L=60.00n
.ENDS CLKNHSV0
****Sub-Circuit for CLKNHSV0P5, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKNHSV0P5 I ZN VDD VSS
MM1 ZN I VSS VPW N12LL W=220.00n L=60.00n
MM0 ZN I VDD VNW P12LL W=450.00n L=60.00n
.ENDS CLKNHSV0P5
****Sub-Circuit for CLKNHSV1, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNHSV1 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=260.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=450.00n L=60.00n
.ENDS CLKNHSV1
****Sub-Circuit for CLKNHSV10, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKNHSV10 I ZN VDD VSS
MM1 ZN I VSS VPW N12LL W=1.6u L=60.00n
MM0 ZN I VDD VNW P12LL W=3.25u L=60.00n
.ENDS CLKNHSV10
****Sub-Circuit for CLKNHSV12, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNHSV12 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=1.86u L=60.00n
MMP1 ZN I VDD VNW P12LL W=3.9u L=60.00n
.ENDS CLKNHSV12
****Sub-Circuit for CLKNHSV16, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNHSV16 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=2.56u L=60.00n
MMP1 ZN I VDD VNW P12LL W=5.2u L=60.00n
.ENDS CLKNHSV16
****Sub-Circuit for CLKNHSV2, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNHSV2 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=360.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=650.00n L=60.00n
.ENDS CLKNHSV2
****Sub-Circuit for CLKNHSV20, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNHSV20 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=3.25u L=60.00n
MMP1 ZN I VDD VNW P12LL W=6.5u L=60.00n
.ENDS CLKNHSV20
****Sub-Circuit for CLKNHSV24, Wed Dec  8 11:21:14 CST 2010****
.SUBCKT CLKNHSV24 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=3.84u L=60.00n
MMP1 ZN I VDD VNW P12LL W=7.8u L=60.00n
.ENDS CLKNHSV24
****Sub-Circuit for CLKNHSV2P5, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKNHSV2P5 I ZN VDD VSS
MM1 ZN I VSS VPW N12LL W=400.00n L=60.00n
MM0 ZN I VDD VNW P12LL W=810.00n L=60.00n
.ENDS CLKNHSV2P5
****Sub-Circuit for CLKNHSV3, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT CLKNHSV3 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=530.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=980.00n L=60.00n
.ENDS CLKNHSV3
****Sub-Circuit for CLKNHSV32, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKNHSV32 I ZN VDD VSS
MM1 ZN I VSS VPW N12LL W=5.12u L=60.00n
MM0 ZN I VDD VNW P12LL W=10.4u L=60.00n
.ENDS CLKNHSV32
****Sub-Circuit for CLKNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT CLKNHSV4 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=710.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=1.3u L=60.00n
.ENDS CLKNHSV4
****Sub-Circuit for CLKNHSV48, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKNHSV48 I ZN VDD VSS
MM1 ZN I VSS VPW N12LL W=7.68u L=60.00n
MM0 ZN I VDD VNW P12LL W=15.6u L=60.00n
.ENDS CLKNHSV48
****Sub-Circuit for CLKNHSV5, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKNHSV5 I ZN VDD VSS
MM1 ZN I VSS VPW N12LL W=800.00n L=60.00n
MM0 ZN I VDD VNW P12LL W=1.62u L=60.00n
.ENDS CLKNHSV5
****Sub-Circuit for CLKNHSV6, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT CLKNHSV6 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=1.02u L=60.00n
MMP1 ZN I VDD VNW P12LL W=1.95u L=60.00n
.ENDS CLKNHSV6
****Sub-Circuit for CLKNHSV64, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT CLKNHSV64 I ZN VDD VSS
MM1 ZN I VSS VPW N12LL W=10.24u L=60.00n
MM0 ZN I VDD VNW P12LL W=20.8u L=60.00n
.ENDS CLKNHSV64
****Sub-Circuit for CLKNHSV8, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT CLKNHSV8 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=1.3u L=60.00n
MMP1 ZN I VDD VNW P12LL W=2.6u L=60.00n
.ENDS CLKNHSV8
****Sub-Circuit for CLKXOR2HSV0, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT CLKXOR2HSV0 A1 A2 Z VDD VSS
MM47 a2n a1n xna1a2 VPW N12LL W=200.00n L=60.00n
MM51 Z xna1a2 VSS VPW N12LL W=200.00n L=60.00n
MM49 a2n A2 VSS VPW N12LL W=200.00n L=60.00n
MM31 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM27 a2nn a2n VSS VPW N12LL W=200.00n L=60.00n
MM36 a2nn A1 xna1a2 VPW N12LL W=200.00n L=60.00n
MM50 a2n A2 VDD VNW P12LL W=350.00n L=60.00n
MM52 Z xna1a2 VDD VNW P12LL W=330.00n L=60.00n
MM48 a2n A1 xna1a2 VNW P12LL W=330.00n L=60.00n
MM32 a1n A1 VDD VNW P12LL W=330.00n L=60.00n
MM28 a2nn a2n VDD VNW P12LL W=350.00n L=60.00n
MM39 a2nn a1n xna1a2 VNW P12LL W=330.00n L=60.00n
.ENDS CLKXOR2HSV0
****Sub-Circuit for CLKXOR2HSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT CLKXOR2HSV1 A1 A2 Z VDD VSS
MM47 a2n a1n xna1a2 VPW N12LL W=200.00n L=60.00n
MM51 Z xna1a2 VSS VPW N12LL W=260.00n L=60.00n
MM49 a2n A2 VSS VPW N12LL W=200.00n L=60.00n
MM31 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM27 a2nn a2n VSS VPW N12LL W=200.00n L=60.00n
MM36 a2nn A1 xna1a2 VPW N12LL W=200.00n L=60.00n
MM50 a2n A2 VDD VNW P12LL W=340.00n L=60.00n
MM52 Z xna1a2 VDD VNW P12LL W=450.00n L=60.00n
MM48 a2n A1 xna1a2 VNW P12LL W=330.00n L=60.00n
MM32 a1n A1 VDD VNW P12LL W=330.00n L=60.00n
MM28 a2nn a2n VDD VNW P12LL W=350.00n L=60.00n
MM39 a2nn a1n xna1a2 VNW P12LL W=330.00n L=60.00n
.ENDS CLKXOR2HSV1
****Sub-Circuit for CLKXOR2HSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT CLKXOR2HSV2 A1 A2 Z VDD VSS
MM47 a2n a1n xna1a2 VPW N12LL W=250.00n L=60.00n
MM51 Z xna1a2 VSS VPW N12LL W=360.00n L=60.00n
MM49 a2n A2 VSS VPW N12LL W=250.00n L=60.00n
MM31 a1n A1 VSS VPW N12LL W=250.00n L=60.00n
MM27 a2nn a2n VSS VPW N12LL W=250.00n L=60.00n
MM36 a2nn A1 xna1a2 VPW N12LL W=250.00n L=60.00n
MM50 a2n A2 VDD VNW P12LL W=460.00n L=60.00n
MM52 Z xna1a2 VDD VNW P12LL W=650.00n L=60.00n
MM48 a2n A1 xna1a2 VNW P12LL W=460.00n L=60.00n
MM32 a1n A1 VDD VNW P12LL W=460.00n L=60.00n
MM28 a2nn a2n VDD VNW P12LL W=460.00n L=60.00n
MM39 a2nn a1n xna1a2 VNW P12LL W=460.00n L=60.00n
.ENDS CLKXOR2HSV2
****Sub-Circuit for CLKXOR2HSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT CLKXOR2HSV4 A1 A2 Z VDD VSS
MM47 a2n a1n xna1a2 VPW N12LL W=300.00n L=60.00n
MM51 Z xna1a2 VSS VPW N12LL W=710.00n L=60.00n
MM49 a2n A2 VSS VPW N12LL W=320.00n L=60.00n
MM31 a1n A1 VSS VPW N12LL W=300.00n L=60.00n
MM27 a2nn a2n VSS VPW N12LL W=320.00n L=60.00n
MM36 a2nn A1 xna1a2 VPW N12LL W=300.00n L=60.00n
MM50 a2n A2 VDD VNW P12LL W=630.00n L=60.00n
MM52 Z xna1a2 VDD VNW P12LL W=1.3u L=60.00n
MM48 a2n A1 xna1a2 VNW P12LL W=450.00n L=60.00n
MM32 a1n A1 VDD VNW P12LL W=450.00n L=60.00n
MM28 a2nn a2n VDD VNW P12LL W=630.00n L=60.00n
MM39 a2nn a1n xna1a2 VNW P12LL W=450.00n L=60.00n
.ENDS CLKXOR2HSV4
****Sub-Circuit for DELHS0, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DELHS0 I Z VDD VSS
MM4 net026 I VSS VPW N12LL W=200.00n L=60.00n
MM5 net022 net026 VSS VPW N12LL W=200.00n L=60.00n
MM0 net13 net022 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=200.00n L=60.00n
MM6 net026 I VDD VNW P12LL W=300.0n L=60.00n
MM7 net022 net026 VDD VNW P12LL W=300.0n L=60.00n
MM1 net13 net022 VDD VNW P12LL W=300.0n L=60.00n
MM3 Z net13 VDD VNW P12LL W=300.00n L=60.00n
.ENDS DELHS0
****Sub-Circuit for DELHS1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DELHS1 I Z VDD VSS
MM4 net026 I VSS VPW N12LL W=200.00n L=60.00n
MM5 net022 net026 VSS VPW N12LL W=200.00n L=60.00n
MM0 net13 net022 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net13 VSS VPW N12LL W=300.00n L=60.00n
MM6 net026 I VDD VNW P12LL W=300.0n L=60.00n
MM7 net022 net026 VDD VNW P12LL W=300.0n L=60.00n
MM1 net13 net022 VDD VNW P12LL W=300.0n L=60.00n
MM3 Z net13 VDD VNW P12LL W=450.00n L=60.00n
.ENDS DELHS1
****Sub-Circuit for DELHS2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DELHS2 I Z VDD VSS
MM4 net026 I VSS VPW N12LL W=200.00n L=60.00n
MM5 net022 net026 VSS VPW N12LL W=200.00n L=120.00n
MM0 net13 net022 VSS VPW N12LL W=200.00n L=120.00n
MM2 Z net13 VSS VPW N12LL W=300.00n L=60.00n
MM6 net026 I VDD VNW P12LL W=300.0n L=60.00n
MM7 net022 net026 VDD VNW P12LL W=300.0n L=120.00n
MM1 net13 net022 VDD VNW P12LL W=300.0n L=120.00n
MM3 Z net13 VDD VNW P12LL W=450.00n L=60.00n
.ENDS DELHS2
****Sub-Circuit for DELHS3, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DELHS3 I Z VDD VSS
MM4 net026 I VSS VPW N12LL W=200.00n L=60.00n
MM5 net022 net026 VSS VPW N12LL W=200.00n L=180.00n
MM0 net13 net022 VSS VPW N12LL W=200.00n L=180.00n
MM2 Z net13 VSS VPW N12LL W=300.00n L=60.00n
MM6 net026 I VDD VNW P12LL W=300.0n L=60.00n
MM7 net022 net026 VDD VNW P12LL W=300.0n L=180.00n
MM1 net13 net022 VDD VNW P12LL W=300.0n L=180.00n
MM3 Z net13 VDD VNW P12LL W=450.00n L=60.00n
.ENDS DELHS3
****Sub-Circuit for DELHS4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DELHS4 I Z VDD VSS
MM4 net026 I VSS VPW N12LL W=200.00n L=60.00n
MM5 net022 net026 VSS VPW N12LL W=200.00n L=240.00n
MM0 net13 net022 VSS VPW N12LL W=200.00n L=240.00n
MM2 Z net13 VSS VPW N12LL W=300.00n L=60.00n
MM6 net026 I VDD VNW P12LL W=300.0n L=60.00n
MM7 net022 net026 VDD VNW P12LL W=300.0n L=240.00n
MM1 net13 net022 VDD VNW P12LL W=300.0n L=240.00n
MM3 Z net13 VDD VNW P12LL W=450.00n L=60.00n
.ENDS DELHS4
****Sub-Circuit for DGRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNHSV1 CK D Q QN RN VDD VSS
MM39 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM3 m c net43 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=250.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=250.00n L=60.00n
MM0 m pm VSS VPW N12LL W=340.00n L=60.00n
MM40 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM4 m cn net43 VNW P12LL W=500.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=330.00n L=60.00n
MM1 m pm VDD VNW P12LL W=500.00n L=60.00n
.ENDS DGRNHSV1
****Sub-Circuit for DGRNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNHSV2 CK D Q QN RN VDD VSS
MM39 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM3 m c net43 VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM40 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM4 m cn net43 VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=450.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS DGRNHSV2
****Sub-Circuit for DGRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNHSV4 CK D Q QN RN VDD VSS
MM39 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM3 m c net43 VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=360.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 m pm VSS VPW N12LL W=390.00n L=60.00n
MM40 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM4 m cn net43 VNW P12LL W=580.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=540.0n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=580.00n L=60.00n
.ENDS DGRNHSV4
****Sub-Circuit for DGRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNQHSV1 CK D Q RN VDD VSS
MM3 m c net43 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=250.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=250.00n L=60.00n
MM0 m pm VSS VPW N12LL W=340.00n L=60.00n
MM4 m cn net43 VNW P12LL W=500.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=330.00n L=60.00n
MM1 m pm VDD VNW P12LL W=500.00n L=60.00n
.ENDS DGRNQHSV1
****Sub-Circuit for DGRNQHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT DGRNQHSV2 CK D Q RN VDD VSS
MM3 m c net43 VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=270.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=270.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM4 m cn net43 VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=450.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=350.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS DGRNQHSV2
****Sub-Circuit for DGRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRNQHSV4 CK D Q RN VDD VSS
MM3 m c net43 VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=340.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=270.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=270.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM4 m cn net43 VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.0n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM10 pm c net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=350.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS DGRNQHSV4
****Sub-Circuit for DGRSNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRSNHSV1 CK D Q QN RN SN VDD VSS
MM43 snn SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN net073 VSS VPW N12LL W=290.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=340.00n L=60.00n
MM42 net69 snn net_0162 VPW N12LL W=250.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=250.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=290.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=250.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=340.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=450.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=380.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=440.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=500.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=440.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=380.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=380.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=500.00n L=60.00n
.ENDS DGRSNHSV1
****Sub-Circuit for DGRSNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRSNHSV2 CK D Q QN RN SN VDD VSS
MM43 snn SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN net073 VSS VPW N12LL W=430.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=360.00n L=60.00n
MM42 net69 snn net_0162 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=430.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=360.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=450.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=650.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=650.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGRSNHSV2
****Sub-Circuit for DGRSNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGRSNHSV4 CK D Q QN RN SN VDD VSS
MM43 snn SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN net073 VSS VPW N12LL W=860.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=360.00n L=60.00n
MM42 net69 snn net_0162 VPW N12LL W=340.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=340.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=860.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=340.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=360.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=450.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=1.3u L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM37 net128 RN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=1.3u L=60.00n
MM18 net063 net073 VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGRSNHSV4
****Sub-Circuit for DGSNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGSNHSV1 CK D Q QN SN VDD VSS
MM39 QN net073 VSS VPW N12LL W=290.00n L=60.00n
MM43 snn SN VSS VPW N12LL W=200.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=270.00n L=60.00n
MM42 net69 snn VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=290.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=250.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=270.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=440.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=440.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=300.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=440.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=440.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=400.00n L=60.00n
.ENDS DGSNHSV1
****Sub-Circuit for DGSNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGSNHSV2 CK D Q QN SN VDD VSS
MM39 QN net073 VSS VPW N12LL W=430.00n L=60.00n
MM43 snn SN VSS VPW N12LL W=200.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=350.00n L=60.00n
MM42 net69 snn VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=380.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=430.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=260.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=260.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=350.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=650.00n L=60.00n
MM44 snn SN VDD VNW P12LL W=300.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=570.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=650.00n L=60.00n
MM18 net063 net073 VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGSNHSV2
****Sub-Circuit for DGSNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DGSNHSV4 CK D Q QN SN VDD VSS
MM39 QN net073 VSS VPW N12LL W=860.00n L=60.00n
MM43 snn SN VSS VPW N12LL W=200.00n L=60.00n
MM3 net049 c net073 VPW N12LL W=340.00n L=60.00n
MM42 net69 snn VSS VPW N12LL W=250.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net073 VPW N12LL W=200.00n L=60.00n
MM23 VSS net063 net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net063 VSS VPW N12LL W=860.00n L=60.00n
MM17 net063 net073 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net051 VPW N12LL W=200.00n L=60.00n
MM11 VSS net049 net52 VPW N12LL W=200.00n L=60.00n
MM9 net051 cn net69 VPW N12LL W=270.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=270.00n L=60.00n
MM0 net049 net051 VSS VPW N12LL W=340.00n L=60.00n
MM41 net_0231 snn VDD VNW P12LL W=510.00n L=60.00n
MM40 QN net073 VDD VNW P12LL W=1.3u L=60.00n
MM44 snn SN VDD VNW P12LL W=300.00n L=60.00n
MM4 net049 cn net073 VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM26 VDD net063 net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net073 VNW P12LL W=300.00n L=60.00n
MM20 Q net063 VDD VNW P12LL W=1.3u L=60.00n
MM18 net063 net073 VDD VNW P12LL W=490.00n L=60.00n
MM14 net117 cn net051 VNW P12LL W=300.00n L=60.00n
MM13 VDD net049 net117 VNW P12LL W=300.00n L=60.00n
MM10 net051 c net128 VNW P12LL W=510.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=510.00n L=60.00n
MM1 net049 net051 VDD VNW P12LL W=510.00n L=60.00n
.ENDS DGSNHSV4
****Sub-Circuit for DHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DHSV1 CK D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=290.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM43 QN s VDD VNW P12LL W=440.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DHSV1
****Sub-Circuit for DHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DHSV2 CK D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=430.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=640.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=640.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DHSV2
****Sub-Circuit for DHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DHSV4 CK D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 net43 c net_099 VPW N12LL W=300.00n L=60.00n m=2
MM40 net_099 m VSS VPW N12LL W=300.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM17 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 net43 cn net_0158 VNW P12LL W=450.00n L=60.00n m=2
MM41 net_0158 m VDD VNW P12LL W=450.00n L=60.00n m=2
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM18 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DHSV4
****Sub-Circuit for DQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DQHSV1 CK D Q VDD VSS
MM39 net43 c net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS DQHSV1
****Sub-Circuit for DQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DQHSV2 CK D Q VDD VSS
MM39 net43 c net_099 VPW N12LL W=430.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=290.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=290.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=440.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=440.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DQHSV2
****Sub-Circuit for DQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DQHSV4 CK D Q VDD VSS
MM39 net43 c net_099 VPW N12LL W=600.0n L=60.00n
MM40 net_099 m VSS VPW N12LL W=600.0n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=290.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=290.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 m pm VSS VPW N12LL W=290.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=910.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=910.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=440.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=440.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DQHSV4
****Sub-Circuit for DRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNHSV1 CK D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DRNHSV1
****Sub-Circuit for DRNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNHSV2 CK D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNHSV2
****Sub-Circuit for DRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNHSV4 CK D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=330.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=330.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNHSV4
****Sub-Circuit for DRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNQHSV1 CK D Q RDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DRNQHSV1
****Sub-Circuit for DRNQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNQHSV2 CK D Q RDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNQHSV2
****Sub-Circuit for DRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DRNQHSV4 CK D Q RDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=330.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=330.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=340.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS DRNQHSV4
****Sub-Circuit for DRSNHSV1, Mon May 30 16:01:10 CST 2011****
.SUBCKT DRSNHSV1 CK D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=290.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=220.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=220.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=360.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=440.00n L=60.00n
.ENDS DRSNHSV1
****Sub-Circuit for DRSNHSV2, Mon May 30 19:07:49 CST 2011****
.SUBCKT DRSNHSV2 CK D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=360.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=380.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=400.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=390.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=220.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=220.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=400.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=600.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=600.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=600.00n L=60.00n
.ENDS DRSNHSV2
****Sub-Circuit for DRSNHSV4, Mon May 30 19:07:49 CST 2011****
.SUBCKT DRSNHSV4 CK D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=360.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=410.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n m=2
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=320.00n L=60.00n m=2
MM40 net43 R net_0132 VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=220.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=220.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 s net43 VDD VNW P12LL W=600.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=650.00n L=60.00n m=2
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=650.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=290.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=290.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=630.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=650.00n L=60.00n
.ENDS DRSNHSV4
****Sub-Circuit for DSNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DSNHSV1 CK D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=400.00n L=60.00n
.ENDS DSNHSV1
****Sub-Circuit for DSNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DSNHSV2 CK D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=300.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=390.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS DSNHSV2
****Sub-Circuit for DSNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DSNHSV4 CK D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=780.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=780.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM38 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=570.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=910.00n L=60.00n
.ENDS DSNHSV4
****Sub-Circuit for DXHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DXHSV1 CK DA DB Q QN SA VDD VSS
MM33 m c net43 VPW N12LL W=350.00n L=60.00n
MM16 net_0144 DB VSS VPW N12LL W=350.00n L=60.00n
MM31 san SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=350.00n L=60.00n
MM19 QN s VSS VPW N12LL W=350.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=310.00n L=60.00n
MM3 net_0148 SA n43 VPW N12LL W=240.00n L=60.00n
MM7 net69 n43 VSS VPW N12LL W=310.00n L=60.00n
MM5 net_0144 san n43 VPW N12LL W=240.00n L=60.00n
MM2 net_0148 DA VSS VPW N12LL W=350.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM38 m cn net43 VNW P12LL W=440.00n L=60.00n
MM37 net_0144 DB VDD VNW P12LL W=440.00n L=60.00n
MM15 net_0148 DA VDD VNW P12LL W=440.00n L=60.00n
MM32 san SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM20 QN s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 n43 VDD VNW P12LL W=390.00n L=60.00n
MM4 net_0148 san n43 VNW P12LL W=300.00n L=60.00n
MM6 net_0144 SA n43 VNW P12LL W=300.00n L=60.00n
MM1 m pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS DXHSV1
****Sub-Circuit for DXHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DXHSV2 CK DA DB Q QN SA VDD VSS
MM5 net_0150 san n43 VPW N12LL W=240.00n L=60.00n
MM2 net_0138 DA VSS VPW N12LL W=350.00n L=60.00n
MM31 san SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM19 QN s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM33 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=310.00n L=60.00n
MM16 net_0150 DB VSS VPW N12LL W=350.00n L=60.00n
MM7 net69 n43 VSS VPW N12LL W=430.00n L=60.00n
MM3 net_0138 SA n43 VPW N12LL W=240.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM15 net_0138 DA VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0150 DB VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0138 san n43 VNW P12LL W=300.00n L=60.00n
MM6 net_0150 SA n43 VNW P12LL W=300.00n L=60.00n
MM32 san SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=550.00n L=60.00n
MM20 QN s VDD VNW P12LL W=550.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 m cn net43 VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 n43 VDD VNW P12LL W=550.00n L=60.00n
MM1 m pm VDD VNW P12LL W=550.00n L=60.00n
.ENDS DXHSV2
****Sub-Circuit for DXHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT DXHSV4 CK DA DB Q QN SA VDD VSS
MM2 net_0156 DA VSS VPW N12LL W=350.00n L=60.00n
MM5 net_0144 san n43 VPW N12LL W=240.00n L=60.00n
MM3 net_0156 SA n43 VPW N12LL W=240.00n L=60.00n
MM16 net_0144 DB VSS VPW N12LL W=350.00n L=60.00n
MM31 san SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM19 QN s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM33 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=260.00n L=60.00n
MM7 net69 n43 VSS VPW N12LL W=260.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM6 net_0144 SA n43 VNW P12LL W=300.00n L=60.00n
MM4 net_0156 san n43 VNW P12LL W=300.00n L=60.00n
MM15 net_0156 DA VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0144 DB VDD VNW P12LL W=440.00n L=60.00n
MM32 san SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.1u L=60.00n
MM20 QN s VDD VNW P12LL W=1.1u L=60.00n
MM18 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM38 m cn net43 VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM10 pm c net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 n43 VDD VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=550.00n L=60.00n
.ENDS DXHSV4
****Sub-Circuit for EDGRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNHSV1 CK D E Q QN RN VDD VSS
MM43 QN s VSS VPW N12LL W=290.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=280.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=280.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM44 QN s VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNHSV1
****Sub-Circuit for EDGRNHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNHSV2 CK D E Q QN RN VDD VSS
MM43 QN s VSS VPW N12LL W=390.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=390.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM44 QN s VDD VNW P12LL W=610.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=610.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=440.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNHSV2
****Sub-Circuit for EDGRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNHSV4 CK D E Q QN RN VDD VSS
MM43 QN s VSS VPW N12LL W=860.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=260.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=260.00n L=60.00n
MM44 QN s VDD VNW P12LL W=1.3u L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=500.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=400.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=400.00n L=60.00n
.ENDS EDGRNHSV4
****Sub-Circuit for EDGRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNQHSV1 CK D E Q RN VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=300.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=280.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=280.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=415.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNQHSV1
****Sub-Circuit for EDGRNQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNQHSV2 CK D E Q RN VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=420.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=420.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=440.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNQHSV2
****Sub-Circuit for EDGRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDGRNQHSV4 CK D E Q RN VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=340.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=340.00n L=60.00n
MM42 net_0164 RN VSS VPW N12LL W=385.00n L=60.00n
MM31 en E VSS VPW N12LL W=300.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.0n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=185.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=185.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=340.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=355.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=340.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=360.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=360.00n L=60.00n
MM39 net_0157 RN VDD VNW P12LL W=200.00n L=60.00n
MM32 en E VDD VNW P12LL W=450.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.0n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=440.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=360.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=360.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=555.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDGRNQHSV4
****Sub-Circuit for EDHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDHSV1 CK D E Q QN VDD VSS
MM43 QN s VSS VPW N12LL W=290.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=395.00n L=60.00n
MM42 QN s VDD VNW P12LL W=440.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=495.00n L=60.00n
.ENDS EDHSV1
****Sub-Circuit for EDHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT EDHSV2 CK D E Q QN VDD VSS
MM43 QN s VSS VPW N12LL W=430.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=340.00n L=60.00n
MM42 QN s VDD VNW P12LL W=650.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=400.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=400.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=550.00n L=60.00n
.ENDS EDHSV2
****Sub-Circuit for EDHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDHSV4 CK D E Q QN VDD VSS
MM43 QN s VSS VPW N12LL W=860.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 QN s VDD VNW P12LL W=1.3u L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDHSV4
****Sub-Circuit for EDQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDQHSV1 CK D E Q VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=395.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=300.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=495.00n L=60.00n
.ENDS EDQHSV1
****Sub-Circuit for EDQHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT EDQHSV2 CK D E Q VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=340.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=400.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=400.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=550.00n L=60.00n
.ENDS EDQHSV2
****Sub-Circuit for EDQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDQHSV4 CK D E Q VDD VSS
MM40 net_0157 s net_0149 VPW N12LL W=290.00n L=60.00n
MM41 net_0149 en VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=430.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=430.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=290.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=390.00n L=60.00n
MM7 net69 E VSS VPW N12LL W=290.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDQHSV4
****Sub-Circuit for EDRNHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNHSV1 CK D E Q QN RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM47 QN s VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM48 QN s VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=320.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=320.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNHSV1
****Sub-Circuit for EDRNHSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT EDRNHSV2 CK D E Q QN RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM47 QN s VSS VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM48 QN s VDD VNW P12LL W=650.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=430.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=430.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNHSV2
****Sub-Circuit for EDRNHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNHSV4 CK D E Q QN RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM47 QN s VSS VPW N12LL W=860.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM48 QN s VDD VNW P12LL W=1.3u L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=420.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNHSV4
****Sub-Circuit for EDRNQHSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNQHSV1 CK D E Q RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=300.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=320.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=320.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNQHSV1
****Sub-Circuit for EDRNQHSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNQHSV2 CK D E Q RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=430.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=430.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNQHSV2
****Sub-Circuit for EDRNQHSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT EDRNQHSV4 CK D E Q RDN VDD VSS
MM45 VSS RDN net_0134 VPW N12LL W=300.00n L=60.00n
MM40 net_0157 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0213 VPW N12LL W=420.00n L=60.00n
MM31 en E VSS VPW N12LL W=240.00n L=60.00n
MM33 net43 c net_0136 VPW N12LL W=400.00n L=60.00n
MM34 net_0136 m VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM44 VSS RDN net_0138 VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=300.00n L=60.00n
MM23 net_0138 s net48 VPW N12LL W=300.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net_0144 VPW N12LL W=300.00n L=60.00n
MM11 net_0134 m net52 VPW N12LL W=300.00n L=60.00n
MM9 net_0157 D net69 VPW N12LL W=420.00n L=60.00n
MM3 net_0157 cn net_0144 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0213 VPW N12LL W=420.00n L=60.00n
MM46 net_0213 RDN VSS VPW N12LL W=420.00n L=60.00n
MM0 m net_0144 VSS VPW N12LL W=400.00n L=60.00n
MM42 VDD RDN net_0144 VNW P12LL W=300.00n L=60.00n
MM43 VDD RDN net43 VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=440.00n L=60.00n
MM38 net_0228 E VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=360.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.3u L=60.00n
MM18 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM35 net43 cn net_0211 VNW P12LL W=460.00n L=60.00n
MM36 net_0211 m VDD VNW P12LL W=460.00n L=60.00n
MM14 net117 cn net_0144 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 en VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0157 c net_0144 VNW P12LL W=600.00n L=60.00n
MM1 m net_0144 VDD VNW P12LL W=600.00n L=60.00n
.ENDS EDRNQHSV4
****Sub-Circuit for FDCAPHS16, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT FDCAPHS16 VDD VSS
MMN1 VSS net13 net14 VPW N12LL W=330.00n L=2.63u
MMP1 net13 net14 VDD VNW P12LL W=550.00n L=2.63u
.ENDS FDCAPHS16
****Sub-Circuit for FDCAPHS32, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT FDCAPHS32 VDD VSS
MMN1 VSS net13 net14 VPW N12LL W=330.00n L=5.83u
MMP1 net13 net14 VDD VNW P12LL W=550.00n L=5.83u
.ENDS FDCAPHS32
****Sub-Circuit for FDCAPHS4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT FDCAPHS4 VDD VSS
MMN1 VSS net13 net14 VPW N12LL W=360.00n L=230.00n
MMP1 net13 net14 VDD VNW P12LL W=580.00n L=230.00n
.ENDS FDCAPHS4
****Sub-Circuit for FDCAPHS64, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT FDCAPHS64 VDD VSS
MMN1 VSS net13 net14 VPW N12LL W=330.00n L=12.23u
MMP1 net13 net14 VDD VNW P12LL W=550.00n L=12.23u
.ENDS FDCAPHS64
****Sub-Circuit for FDCAPHS8, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT FDCAPHS8 VDD VSS
MMN1 VSS net13 net14 VPW N12LL W=330.00n L=1.03u
MMP1 net13 net14 VDD VNW P12LL W=550.00n L=1.03u
.ENDS FDCAPHS8
****Sub-Circuit for FILLTIEHS, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT FILLTIEHS VDD VSS
.ENDS FILLTIEHS
****Sub-Circuit for F_FILLHS1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT F_FILLHS1 VDD VSS
.ENDS F_FILLHS1
****Sub-Circuit for F_FILLHS16, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT F_FILLHS16 VDD VSS
.ENDS F_FILLHS16
****Sub-Circuit for F_FILLHS2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT F_FILLHS2 VDD VSS
.ENDS F_FILLHS2
****Sub-Circuit for F_FILLHS4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT F_FILLHS4 VDD VSS
.ENDS F_FILLHS4
****Sub-Circuit for F_FILLHS8, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT F_FILLHS8 VDD VSS
.ENDS F_FILLHS8
****Sub-Circuit for I2NAND4HSV0, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT I2NAND4HSV0 A1 A2 B1 B2 ZN VDD VSS
MM9 a2n A2 VSS VPW N12LL W=200.00n L=60.00n
MM6 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM3 net031 B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN a1n net18 VPW N12LL W=200.00n L=60.00n
MM2 net039 B1 net031 VPW N12LL W=200.00n L=60.00n
MMN1 net18 a2n net039 VPW N12LL W=200.00n L=60.00n
MM8 a2n A2 VDD VNW P12LL W=300.00n L=60.00n
MM7 a1n A1 VDD VNW P12LL W=300.00n L=60.00n
MM4 ZN B2 VDD VNW P12LL W=300.00n L=60.00n
MM5 ZN B1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN a2n VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN a1n VDD VNW P12LL W=300.00n L=60.00n
.ENDS I2NAND4HSV0
****Sub-Circuit for I2NAND4HSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT I2NAND4HSV1 A1 A2 B1 B2 ZN VDD VSS
MM9 a2n A2 VSS VPW N12LL W=200.00n L=60.00n
MM6 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM3 net031 B2 VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN a1n net18 VPW N12LL W=290.00n L=60.00n
MM2 net039 B1 net031 VPW N12LL W=290.00n L=60.00n
MMN1 net18 a2n net039 VPW N12LL W=290.00n L=60.00n
MM8 a2n A2 VDD VNW P12LL W=300.00n L=60.00n
MM7 a1n A1 VDD VNW P12LL W=300.00n L=60.00n
MM4 ZN B2 VDD VNW P12LL W=440.00n L=60.00n
MM5 ZN B1 VDD VNW P12LL W=440.00n L=60.00n
MM0 ZN a2n VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN a1n VDD VNW P12LL W=440.00n L=60.00n
.ENDS I2NAND4HSV1
****Sub-Circuit for I2NAND4HSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT I2NAND4HSV2 A1 A2 B1 B2 ZN VDD VSS
MM9 a2n A2 VSS VPW N12LL W=200.00n L=60.00n
MM6 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM3 net031 B2 VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN a1n net18 VPW N12LL W=430.00n L=60.00n
MM2 net039 B1 net031 VPW N12LL W=430.00n L=60.00n
MMN1 net18 a2n net039 VPW N12LL W=430.00n L=60.00n
MM8 a2n A2 VDD VNW P12LL W=300.00n L=60.00n
MM7 a1n A1 VDD VNW P12LL W=300.00n L=60.00n
MM4 ZN B2 VDD VNW P12LL W=650.00n L=60.00n
MM5 ZN B1 VDD VNW P12LL W=650.00n L=60.00n
MM0 ZN a2n VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN a1n VDD VNW P12LL W=650.00n L=60.00n
.ENDS I2NAND4HSV2
****Sub-Circuit for I2NAND4HSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT I2NAND4HSV4 A1 A2 B1 B2 ZN VDD VSS
MM9 a2n A2 VSS VPW N12LL W=350.00n L=60.00n
MM6 a1n A1 VSS VPW N12LL W=350.00n L=60.00n
MM3 net031 B2 VSS VPW N12LL W=860.00n L=60.00n
MM1 ZN a1n net18 VPW N12LL W=860.00n L=60.00n
MM2 net039 B1 net031 VPW N12LL W=860.00n L=60.00n
MMN1 net18 a2n net039 VPW N12LL W=860.00n L=60.00n
MM8 a2n A2 VDD VNW P12LL W=520.00n L=60.00n
MM7 a1n A1 VDD VNW P12LL W=520.00n L=60.00n
MM4 ZN B2 VDD VNW P12LL W=1.29u L=60.00n
MM5 ZN B1 VDD VNW P12LL W=1.29u L=60.00n
MM0 ZN a2n VDD VNW P12LL W=1.29u L=60.00n
MMP1 ZN a1n VDD VNW P12LL W=1.29u L=60.00n
.ENDS I2NAND4HSV4
****Sub-Circuit for I2NOR4HSV0, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT I2NOR4HSV0 A1 A2 B1 B2 ZN VDD VSS
MM9 a2n A2 VSS VPW N12LL W=200.00n L=60.00n
MM6 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM3 ZN B2 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN a1n VSS VPW N12LL W=200.00n L=60.00n
MM2 ZN B1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 ZN a2n VSS VPW N12LL W=200.00n L=60.00n
MM8 a2n A2 VDD VNW P12LL W=300.0n L=60.00n
MM7 a1n A1 VDD VNW P12LL W=300.0n L=60.00n
MM4 net0139 B1 net0143 VNW P12LL W=300.0n L=60.00n
MM5 ZN B2 net0139 VNW P12LL W=300.0n L=60.00n
MM0 net0147 a1n VDD VNW P12LL W=300.0n L=60.00n
MMP1 net0143 a2n net0147 VNW P12LL W=300.0n L=60.00n
.ENDS I2NOR4HSV0
****Sub-Circuit for I2NOR4HSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT I2NOR4HSV1 A1 A2 B1 B2 ZN VDD VSS
MM9 a2n A2 VSS VPW N12LL W=200.00n L=60.00n
MM6 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM3 ZN B2 VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN a1n VSS VPW N12LL W=290.00n L=60.00n
MM2 ZN B1 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN a2n VSS VPW N12LL W=290.00n L=60.00n
MM8 a2n A2 VDD VNW P12LL W=300.00n L=60.00n
MM7 a1n A1 VDD VNW P12LL W=300.00n L=60.00n
MM4 net0139 B1 net0143 VNW P12LL W=440.00n L=60.00n
MM5 ZN B2 net0139 VNW P12LL W=440.00n L=60.00n
MM0 net0147 a1n VDD VNW P12LL W=440.00n L=60.00n
MMP1 net0143 a2n net0147 VNW P12LL W=440.00n L=60.00n
.ENDS I2NOR4HSV1
****Sub-Circuit for I2NOR4HSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT I2NOR4HSV2 A1 A2 B1 B2 ZN VDD VSS
MM9 a2n A2 VSS VPW N12LL W=200.00n L=60.00n
MM6 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM3 ZN B2 VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN a1n VSS VPW N12LL W=430.00n L=60.00n
MM2 ZN B1 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN a2n VSS VPW N12LL W=430.00n L=60.00n
MM8 a2n A2 VDD VNW P12LL W=300.00n L=60.00n
MM7 a1n A1 VDD VNW P12LL W=300.00n L=60.00n
MM4 net0139 B1 net0143 VNW P12LL W=650.00n L=60.00n
MM5 ZN B2 net0139 VNW P12LL W=650.00n L=60.00n
MM0 net0147 a1n VDD VNW P12LL W=650.00n L=60.00n
MMP1 net0143 a2n net0147 VNW P12LL W=650.00n L=60.00n
.ENDS I2NOR4HSV2
****Sub-Circuit for I2NOR4HSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT I2NOR4HSV4 A1 A2 B1 B2 ZN VDD VSS
MM9 a2n A2 VSS VPW N12LL W=350.00n L=60.00n
MM6 a1n A1 VSS VPW N12LL W=350.00n L=60.00n
MM3 ZN B2 VSS VPW N12LL W=860.00n L=60.00n
MM1 ZN a1n VSS VPW N12LL W=860.00n L=60.00n
MM2 ZN B1 VSS VPW N12LL W=860.00n L=60.00n
MMN1 ZN a2n VSS VPW N12LL W=860.00n L=60.00n
MM8 a2n A2 VDD VNW P12LL W=520.00n L=60.00n
MM7 a1n A1 VDD VNW P12LL W=520.00n L=60.00n
MM4 net0139 B1 net0143 VNW P12LL W=1.3u L=60.00n
MM5 ZN B2 net0139 VNW P12LL W=1.3u L=60.00n
MM0 net0147 a1n VDD VNW P12LL W=1.3u L=60.00n
MMP1 net0143 a2n net0147 VNW P12LL W=1.3u L=60.00n
.ENDS I2NOR4HSV4
****Sub-Circuit for IAO21HSV0, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT IAO21HSV0 A1 A2 B ZN VDD VSS
MM3 net24 A1 VSS VPW N12LL W=200.00n L=60.00n
MM2 net24 A2 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN B VSS VPW N12LL W=200.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=200.00n L=60.00n
MM4 net24 A1 net056 VNW P12LL W=300.00n L=60.00n
MM5 net056 A2 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net24 net064 VNW P12LL W=300.00n L=60.00n
MMP1 net064 B VDD VNW P12LL W=300.00n L=60.00n
.ENDS IAO21HSV0
****Sub-Circuit for IAO21HSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT IAO21HSV1 A1 A2 B ZN VDD VSS
MM3 net24 A1 VSS VPW N12LL W=200.00n L=60.00n
MM2 net24 A2 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN B VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=290.00n L=60.00n
MM4 net24 A1 net056 VNW P12LL W=300.00n L=60.00n
MM5 net056 A2 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net24 net064 VNW P12LL W=440.00n L=60.00n
MMP1 net064 B VDD VNW P12LL W=440.00n L=60.00n
.ENDS IAO21HSV1
****Sub-Circuit for IAO21HSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT IAO21HSV2 A1 A2 B ZN VDD VSS
MM3 net24 A1 VSS VPW N12LL W=200.00n L=60.00n
MM2 net24 A2 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN B VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=430.00n L=60.00n
MM4 net24 A1 net056 VNW P12LL W=300.00n L=60.00n
MM5 net056 A2 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net24 net064 VNW P12LL W=650.00n L=60.00n
MMP1 net064 B VDD VNW P12LL W=650.00n L=60.00n
.ENDS IAO21HSV2
****Sub-Circuit for IAO21HSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT IAO21HSV4 A1 A2 B ZN VDD VSS
MM3 net24 A1 VSS VPW N12LL W=350.00n L=60.00n
MM2 net24 A2 VSS VPW N12LL W=350.00n L=60.00n
MM0 ZN B VSS VPW N12LL W=720.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=720.00n L=60.00n
MM4 net24 A1 net056 VNW P12LL W=520.00n L=60.00n
MM5 net056 A2 VDD VNW P12LL W=520.00n L=60.00n
MM1 ZN net24 net064 VNW P12LL W=1.2u L=60.00n
MMP1 net064 B VDD VNW P12LL W=1.2u L=60.00n
.ENDS IAO21HSV4
****Sub-Circuit for IAO22HSV0, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT IAO22HSV0 A1 A2 B1 B2 ZN VDD VSS
MM3 net24 A1 VSS VPW N12LL W=200.00n L=60.00n
MM2 net24 A2 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN B1 net050 VPW N12LL W=200.00n L=60.00n
MM7 net050 B2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=200.00n L=60.00n
MM6 net061 B2 VDD VNW P12LL W=300.00n L=60.00n
MM4 net24 A1 net074 VNW P12LL W=300.00n L=60.00n
MM5 net074 A2 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net24 net061 VNW P12LL W=300.00n L=60.00n
MMP1 net061 B1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS IAO22HSV0
****Sub-Circuit for IAO22HSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT IAO22HSV1 A1 A2 B1 B2 ZN VDD VSS
MM3 net24 A1 VSS VPW N12LL W=200.00n L=60.00n
MM2 net24 A2 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN B1 net050 VPW N12LL W=290.00n L=60.00n
MM7 net050 B2 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=290.00n L=60.00n
MM6 net061 B2 VDD VNW P12LL W=440.00n L=60.00n
MM4 net24 A1 net074 VNW P12LL W=300.00n L=60.00n
MM5 net074 A2 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net24 net061 VNW P12LL W=440.00n L=60.00n
MMP1 net061 B1 VDD VNW P12LL W=440.00n L=60.00n
.ENDS IAO22HSV1
****Sub-Circuit for IAO22HSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT IAO22HSV2 A1 A2 B1 B2 ZN VDD VSS
MM3 net24 A1 VSS VPW N12LL W=200.00n L=60.00n
MM2 net24 A2 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN B1 net050 VPW N12LL W=430.00n L=60.00n
MM7 net050 B2 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=430.00n L=60.00n
MM6 net061 B2 VDD VNW P12LL W=650.00n L=60.00n
MM4 net24 A1 net074 VNW P12LL W=300.00n L=60.00n
MM5 net074 A2 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net24 net061 VNW P12LL W=650.00n L=60.00n
MMP1 net061 B1 VDD VNW P12LL W=650.00n L=60.00n
.ENDS IAO22HSV2
****Sub-Circuit for IAO22HSV4, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT IAO22HSV4 A1 A2 B1 B2 ZN VDD VSS
MM3 net24 A1 VSS VPW N12LL W=350.00n L=60.00n
MM2 net24 A2 VSS VPW N12LL W=350.00n L=60.00n
MM0 ZN B1 net050 VPW N12LL W=860.00n L=60.00n
MM7 net050 B2 VSS VPW N12LL W=860.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=860.00n L=60.00n
MM6 net061 B2 VDD VNW P12LL W=1.24u L=60.00n
MM4 net24 A1 net074 VNW P12LL W=520.00n L=60.00n
MM5 net074 A2 VDD VNW P12LL W=520.00n L=60.00n
MM1 ZN net24 net061 VNW P12LL W=1.3u L=60.00n
MMP1 net061 B1 VDD VNW P12LL W=1.24u L=60.00n
.ENDS IAO22HSV4
****Sub-Circuit for INAND2HSV0, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT INAND2HSV0 A1 B1 ZN VDD VSS
MM3 net021 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 B1 VSS VPW N12LL W=200.00n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=300.00n L=60.00n
.ENDS INAND2HSV0
****Sub-Circuit for INAND2HSV1, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT INAND2HSV1 A1 B1 ZN VDD VSS
MM3 net021 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=290.0n L=60.00n
MMN1 net18 B1 VSS VPW N12LL W=290.0n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=440.0n L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=440.0n L=60.00n
.ENDS INAND2HSV1
****Sub-Circuit for INAND2HSV2, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT INAND2HSV2 A1 B1 ZN VDD VSS
MM3 net021 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=430.00n L=60.00n
MMN1 net18 B1 VSS VPW N12LL W=430.00n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=650.00n L=60.00n
.ENDS INAND2HSV2
****Sub-Circuit for INAND2HSV4, Wed Dec  8 11:21:15 CST 2010****
.SUBCKT INAND2HSV4 A1 B1 ZN VDD VSS
MM3 net021 A1 VSS VPW N12LL W=340.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=820.00n L=60.00n
MMN1 net18 B1 VSS VPW N12LL W=820.00n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=510.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=1.26u L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=1.26u L=60.00n
.ENDS INAND2HSV4
****Sub-Circuit for INAND3HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INAND3HSV0 A1 B1 B2 ZN VDD VSS
MM5 net029 B2 VSS VPW N12LL W=200.00n L=60.00n
MM3 net021 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 B1 net029 VPW N12LL W=200.00n L=60.00n
MM6 ZN B2 VDD VNW P12LL W=300.00n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=300.00n L=60.00n
.ENDS INAND3HSV0
****Sub-Circuit for INAND3HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INAND3HSV1 A1 B1 B2 ZN VDD VSS
MM5 net029 B2 VSS VPW N12LL W=290.00n L=60.00n
MM3 net021 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=290.00n L=60.00n
MMN1 net18 B1 net029 VPW N12LL W=290.00n L=60.00n
MM6 ZN B2 VDD VNW P12LL W=440.00n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=440.00n L=60.00n
.ENDS INAND3HSV1
****Sub-Circuit for INAND3HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INAND3HSV2 A1 B1 B2 ZN VDD VSS
MM5 net029 B2 VSS VPW N12LL W=430.00n L=60.00n
MM3 net021 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=430.00n L=60.00n
MMN1 net18 B1 net029 VPW N12LL W=430.00n L=60.00n
MM6 ZN B2 VDD VNW P12LL W=650.00n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=650.00n L=60.00n
.ENDS INAND3HSV2
****Sub-Circuit for INAND3HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INAND3HSV4 A1 B1 B2 ZN VDD VSS
MM5 net029 B2 VSS VPW N12LL W=860.00n L=60.00n
MM3 net021 A1 VSS VPW N12LL W=340.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=860.00n L=60.00n
MMN1 net18 B1 net029 VPW N12LL W=860.00n L=60.00n
MM6 ZN B2 VDD VNW P12LL W=1.29u L=60.00n
MM4 net021 A1 VDD VNW P12LL W=510.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=1.29u L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=1.29u L=60.00n
.ENDS INAND3HSV4
****Sub-Circuit for INAND4HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INAND4HSV0 A1 B1 B2 B3 ZN VDD VSS
MM8 net040 B3 VSS VPW N12LL W=200.00n L=60.00n
MM5 net029 B2 net040 VPW N12LL W=200.00n L=60.00n
MM3 net021 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 B1 net029 VPW N12LL W=200.00n L=60.00n
MM7 ZN B3 VDD VNW P12LL W=300.00n L=60.00n
MM6 ZN B2 VDD VNW P12LL W=300.00n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=300.00n L=60.00n
.ENDS INAND4HSV0
****Sub-Circuit for INAND4HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INAND4HSV1 A1 B1 B2 B3 ZN VDD VSS
MM8 net040 B3 VSS VPW N12LL W=290.00n L=60.00n
MM5 net029 B2 net040 VPW N12LL W=290.00n L=60.00n
MM3 net021 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=290.00n L=60.00n
MMN1 net18 B1 net029 VPW N12LL W=290.00n L=60.00n
MM7 ZN B3 VDD VNW P12LL W=440.00n L=60.00n
MM6 ZN B2 VDD VNW P12LL W=440.00n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=440.00n L=60.00n
.ENDS INAND4HSV1
****Sub-Circuit for INAND4HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INAND4HSV2 A1 B1 B2 B3 ZN VDD VSS
MM8 net040 B3 VSS VPW N12LL W=430.00n L=60.00n
MM5 net029 B2 net040 VPW N12LL W=430.00n L=60.00n
MM3 net021 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=430.00n L=60.00n
MMN1 net18 B1 net029 VPW N12LL W=430.00n L=60.00n
MM7 ZN B3 VDD VNW P12LL W=650.00n L=60.00n
MM6 ZN B2 VDD VNW P12LL W=650.00n L=60.00n
MM4 net021 A1 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=650.00n L=60.00n
.ENDS INAND4HSV2
****Sub-Circuit for INAND4HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INAND4HSV4 A1 B1 B2 B3 ZN VDD VSS
MM8 net040 B3 VSS VPW N12LL W=860.00n L=60.00n
MM5 net029 B2 net040 VPW N12LL W=860.00n L=60.00n
MM3 net021 A1 VSS VPW N12LL W=340.00n L=60.00n
MM1 ZN net021 net18 VPW N12LL W=860.00n L=60.00n
MMN1 net18 B1 net029 VPW N12LL W=860.00n L=60.00n
MM7 ZN B3 VDD VNW P12LL W=1.29u L=60.00n
MM6 ZN B2 VDD VNW P12LL W=1.29u L=60.00n
MM4 net021 A1 VDD VNW P12LL W=510.00n L=60.00n
MM0 ZN B1 VDD VNW P12LL W=1.29u L=60.00n
MMP1 ZN net021 VDD VNW P12LL W=1.29u L=60.00n
.ENDS INAND4HSV4
****Sub-Circuit for INHSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV0 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=200.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=300.00n L=60.00n
.ENDS INHSV0
****Sub-Circuit for INHSV0P5, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT INHSV0P5 I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=370.00n L=60.00n
MM1 ZN I VSS VPW N12LL W=240.00n L=60.00n
.ENDS INHSV0P5
****Sub-Circuit for INHSV0P5SR, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT INHSV0P5SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=350.00n L=60.00n
MM1 ZN I VSS VPW N12LL W=280.00n L=60.00n
.ENDS INHSV0P5SR
****Sub-Circuit for INHSV0SR, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT INHSV0SR I ZN VDD VSS
MM1 ZN I VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN I VDD VNW P12LL W=250.00n L=60.00n
.ENDS INHSV0SR
****Sub-Circuit for INHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV1 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=290.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=440.00n L=60.00n
.ENDS INHSV1
****Sub-Circuit for INHSV10, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT INHSV10 I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=3.25u L=60.00n
MM1 ZN I VSS VPW N12LL W=2.15u L=60.00n
.ENDS INHSV10
****Sub-Circuit for INHSV10SR, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT INHSV10SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=2.7u L=60.00n
MM1 ZN I VSS VPW N12LL W=2.15u L=60.00n
.ENDS INHSV10SR
****Sub-Circuit for INHSV12, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV12 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=2.58u L=60.00n
MMP1 ZN I VDD VNW P12LL W=3.9u L=60.00n
.ENDS INHSV12
****Sub-Circuit for INHSV12SR, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT INHSV12SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=3.24u L=60.00n
MM1 ZN I VSS VPW N12LL W=2.58u L=60.00n
.ENDS INHSV12SR
****Sub-Circuit for INHSV16, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV16 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=3.44u L=60.00n
MMP1 ZN I VDD VNW P12LL W=5.20u L=60.00n
.ENDS INHSV16
****Sub-Circuit for INHSV16SR, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT INHSV16SR I ZN VDD VSS
MM1 ZN I VSS VPW N12LL W=3.44u L=60.00n
MM0 ZN I VDD VNW P12LL W=4.32u L=60.00n
.ENDS INHSV16SR
****Sub-Circuit for INHSV1SR, Wed Dec  8 16:10:27 CST 2010****
.SUBCKT INHSV1SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=440.00n L=60.00n
MM1 ZN I VSS VPW N12LL W=350.00n L=60.00n
.ENDS INHSV1SR
****Sub-Circuit for INHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV2 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=430.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=650.00n L=60.00n
.ENDS INHSV2
****Sub-Circuit for INHSV20, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV20 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=4.3u L=60.00n
MMP1 ZN I VDD VNW P12LL W=6.50u L=60.00n
.ENDS INHSV20
****Sub-Circuit for INHSV20SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV20SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=5.4u L=60.00n
MM1 ZN I VSS VPW N12LL W=4.3u L=60.00n
.ENDS INHSV20SR
****Sub-Circuit for INHSV24, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV24 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=5.16u L=60.00n
MMP1 ZN I VDD VNW P12LL W=7.80u L=60.00n
.ENDS INHSV24
****Sub-Circuit for INHSV24SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV24SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=6.48u L=60.00n
MM1 ZN I VSS VPW N12LL W=5.16u L=60.00n
.ENDS INHSV24SR
****Sub-Circuit for INHSV2P5, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV2P5 I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=810.00n L=60.00n
MM1 ZN I VSS VPW N12LL W=540.00n L=60.00n
.ENDS INHSV2P5
****Sub-Circuit for INHSV2SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV2SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=540.00n L=60.00n
MM1 ZN I VSS VPW N12LL W=430.00n L=60.00n
.ENDS INHSV2SR
****Sub-Circuit for INHSV3, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV3 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=650.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=980.00n L=60.00n
.ENDS INHSV3
****Sub-Circuit for INHSV32, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV32 I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=10.4u L=60.00n
MM1 ZN I VSS VPW N12LL W=6.88u L=60.00n
.ENDS INHSV32
****Sub-Circuit for INHSV32SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV32SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=8.64u L=60.00n
MM1 ZN I VSS VPW N12LL W=6.88u L=60.00n
.ENDS INHSV32SR
****Sub-Circuit for INHSV3SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV3SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=810.00n L=60.00n
MM1 ZN I VSS VPW N12LL W=650.00n L=60.00n
.ENDS INHSV3SR
****Sub-Circuit for INHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV4 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=860.00n L=60.00n
MMP1 ZN I VDD VNW P12LL W=1.3u L=60.00n
.ENDS INHSV4
****Sub-Circuit for INHSV48, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV48 I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=15.6u L=60.00n
MM1 ZN I VSS VPW N12LL W=10.32u L=60.00n
.ENDS INHSV48
****Sub-Circuit for INHSV48SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV48SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=12.96u L=60.00n
MM1 ZN I VSS VPW N12LL W=10.32u L=60.00n
.ENDS INHSV48SR
****Sub-Circuit for INHSV4SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV4SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=1.08u L=60.00n
MM1 ZN I VSS VPW N12LL W=860.00n L=60.00n
.ENDS INHSV4SR
****Sub-Circuit for INHSV5, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV5 I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=1.62u L=60.00n
MM1 ZN I VSS VPW N12LL W=1.07u L=60.00n
.ENDS INHSV5
****Sub-Circuit for INHSV5SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV5SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=1.35u L=60.00n
MM1 ZN I VSS VPW N12LL W=1.08u L=60.00n
.ENDS INHSV5SR
****Sub-Circuit for INHSV6, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV6 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=1.29u L=60.00n
MMP1 ZN I VDD VNW P12LL W=1.95u L=60.00n
.ENDS INHSV6
****Sub-Circuit for INHSV64, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV64 I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=20.8u L=60.00n
MM1 ZN I VSS VPW N12LL W=13.76u L=60.00n
.ENDS INHSV64
****Sub-Circuit for INHSV64SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV64SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=17.28u L=60.00n
MM1 ZN I VSS VPW N12LL W=13.76u L=60.00n
.ENDS INHSV64SR
****Sub-Circuit for INHSV6SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV6SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=1.62u L=60.00n
MM1 ZN I VSS VPW N12LL W=1.29u L=60.00n
.ENDS INHSV6SR
****Sub-Circuit for INHSV8, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INHSV8 I ZN VDD VSS
MMN1 ZN I VSS VPW N12LL W=1.72u L=60.00n
MMP1 ZN I VDD VNW P12LL W=2.6u L=60.00n
.ENDS INHSV8
****Sub-Circuit for INHSV8SR, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT INHSV8SR I ZN VDD VSS
MM0 ZN I VDD VNW P12LL W=2.16u L=60.00n
MM1 ZN I VSS VPW N12LL W=1.72u L=60.00n
.ENDS INHSV8SR
****Sub-Circuit for INOR2HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR2HSV0 A1 B1 ZN VDD VSS
MM2 net27 A1 VSS VPW N12LL W=200.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=200.0n L=60.00n
MMN1 ZN net27 VSS VPW N12LL W=200.0n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=300.00n L=60.00n
MM3 net27 A1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 B1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS INOR2HSV0
****Sub-Circuit for INOR2HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR2HSV1 A1 B1 ZN VDD VSS
MM2 net27 A1 VSS VPW N12LL W=200.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN net27 VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=440.00n L=60.00n
MM3 net27 A1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 B1 VDD VNW P12LL W=440.00n L=60.00n
.ENDS INOR2HSV1
****Sub-Circuit for INOR2HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR2HSV2 A1 B1 ZN VDD VSS
MM2 net27 A1 VSS VPW N12LL W=200.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN net27 VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=650.00n L=60.00n
MM3 net27 A1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 B1 VDD VNW P12LL W=650.00n L=60.00n
.ENDS INOR2HSV2
****Sub-Circuit for INOR2HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR2HSV4 A1 B1 ZN VDD VSS
MM2 net27 A1 VSS VPW N12LL W=350.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=860.00n L=60.00n
MMN1 ZN net27 VSS VPW N12LL W=860.00n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=1.3u L=60.00n
MM3 net27 A1 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net42 B1 VDD VNW P12LL W=1.3u L=60.00n
.ENDS INOR2HSV4
****Sub-Circuit for INOR3HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR3HSV0 A1 B1 B2 ZN VDD VSS
MM5 ZN net27 VSS VPW N12LL W=200.0n L=60.00n
MM2 net27 A1 VSS VPW N12LL W=200.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=200.0n L=60.00n
MMN1 ZN B2 VSS VPW N12LL W=200.0n L=60.00n
MM4 net061 B2 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=300.00n L=60.00n
MM3 net27 A1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 B1 net061 VNW P12LL W=300.00n L=60.00n
.ENDS INOR3HSV0
****Sub-Circuit for INOR3HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR3HSV1 A1 B1 B2 ZN VDD VSS
MM5 ZN net27 VSS VPW N12LL W=290.00n L=60.00n
MM2 net27 A1 VSS VPW N12LL W=200.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN B2 VSS VPW N12LL W=290.00n L=60.00n
MM4 net061 B2 VDD VNW P12LL W=440.00n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=440.00n L=60.00n
MM3 net27 A1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 B1 net061 VNW P12LL W=440.00n L=60.00n
.ENDS INOR3HSV1
****Sub-Circuit for INOR3HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR3HSV2 A1 B1 B2 ZN VDD VSS
MM5 ZN net27 VSS VPW N12LL W=430.00n L=60.00n
MM2 net27 A1 VSS VPW N12LL W=200.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN B2 VSS VPW N12LL W=430.00n L=60.00n
MM4 net061 B2 VDD VNW P12LL W=650.00n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=650.00n L=60.00n
MM3 net27 A1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 B1 net061 VNW P12LL W=650.00n L=60.00n
.ENDS INOR3HSV2
****Sub-Circuit for INOR3HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR3HSV4 A1 B1 B2 ZN VDD VSS
MM5 ZN net27 VSS VPW N12LL W=860.00n L=60.00n
MM2 net27 A1 VSS VPW N12LL W=350.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=860.00n L=60.00n
MMN1 ZN B2 VSS VPW N12LL W=860.00n L=60.00n
MM4 net061 B2 VDD VNW P12LL W=1.3u L=60.00n
MM1 ZN net27 net42 VNW P12LL W=1.3u L=60.00n
MM3 net27 A1 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net42 B1 net061 VNW P12LL W=1.3u L=60.00n
.ENDS INOR3HSV4
****Sub-Circuit for INOR4HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR4HSV0 A1 B1 B2 B3 ZN VDD VSS
MM7 ZN B3 VSS VPW N12LL W=200.0n L=60.00n
MM5 ZN net27 VSS VPW N12LL W=200.0n L=60.00n
MM2 net27 A1 VSS VPW N12LL W=200.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=200.0n L=60.00n
MMN1 ZN B2 VSS VPW N12LL W=200.0n L=60.00n
MM4 net061 B2 net070 VNW P12LL W=300.0n L=60.00n
MM6 net070 B3 VDD VNW P12LL W=300.0n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=300.0n L=60.00n
MM3 net27 A1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 B1 net061 VNW P12LL W=300.0n L=60.00n
.ENDS INOR4HSV0
****Sub-Circuit for INOR4HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR4HSV1 A1 B1 B2 B3 ZN VDD VSS
MM7 ZN B3 VSS VPW N12LL W=290.00n L=60.00n
MM5 ZN net27 VSS VPW N12LL W=290.00n L=60.00n
MM2 net27 A1 VSS VPW N12LL W=200.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN B2 VSS VPW N12LL W=290.00n L=60.00n
MM4 net061 B2 net070 VNW P12LL W=440.00n L=60.00n
MM6 net070 B3 VDD VNW P12LL W=440.00n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=440.00n L=60.00n
MM3 net27 A1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 B1 net061 VNW P12LL W=440.00n L=60.00n
.ENDS INOR4HSV1
****Sub-Circuit for INOR4HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR4HSV2 A1 B1 B2 B3 ZN VDD VSS
MM7 ZN B3 VSS VPW N12LL W=430.00n L=60.00n
MM5 ZN net27 VSS VPW N12LL W=430.00n L=60.00n
MM2 net27 A1 VSS VPW N12LL W=200.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN B2 VSS VPW N12LL W=430.00n L=60.00n
MM4 net061 B2 net070 VNW P12LL W=650.00n L=60.00n
MM6 net070 B3 VDD VNW P12LL W=650.00n L=60.00n
MM1 ZN net27 net42 VNW P12LL W=650.00n L=60.00n
MM3 net27 A1 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 B1 net061 VNW P12LL W=650.00n L=60.00n
.ENDS INOR4HSV2
****Sub-Circuit for INOR4HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT INOR4HSV4 A1 B1 B2 B3 ZN VDD VSS
MM7 ZN B3 VSS VPW N12LL W=860.00n L=60.00n
MM5 ZN net27 VSS VPW N12LL W=860.00n L=60.00n
MM2 net27 A1 VSS VPW N12LL W=350.0n L=60.00n
MM0 ZN B1 VSS VPW N12LL W=860.00n L=60.00n
MMN1 ZN B2 VSS VPW N12LL W=860.00n L=60.00n
MM4 net061 B2 net070 VNW P12LL W=1.3u L=60.00n
MM6 net070 B3 VDD VNW P12LL W=1.3u L=60.00n
MM1 ZN net27 net42 VNW P12LL W=1.3u L=60.00n
MM3 net27 A1 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net42 B1 net061 VNW P12LL W=1.3u L=60.00n
.ENDS INOR4HSV4
****Sub-Circuit for IOA21HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT IOA21HSV0 A1 A2 B ZN VDD VSS
MM2 ZN net038 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 B VSS VPW N12LL W=200.00n L=60.00n
MM1 net038 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=300.00n L=60.00n
MM5 ZN net038 VDD VNW P12LL W=300.00n L=60.00n
MM0 net038 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net038 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS IOA21HSV0
****Sub-Circuit for IOA21HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT IOA21HSV1 A1 A2 B ZN VDD VSS
MM2 ZN net038 net030 VPW N12LL W=290.00n L=60.00n
MM3 net030 B VSS VPW N12LL W=290.00n L=60.00n
MM1 net038 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=440.00n L=60.00n
MM5 ZN net038 VDD VNW P12LL W=440.00n L=60.00n
MM0 net038 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net038 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS IOA21HSV1
****Sub-Circuit for IOA21HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT IOA21HSV2 A1 A2 B ZN VDD VSS
MM2 ZN net038 net030 VPW N12LL W=430.00n L=60.00n
MM3 net030 B VSS VPW N12LL W=430.00n L=60.00n
MM1 net038 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=650.00n L=60.00n
MM5 ZN net038 VDD VNW P12LL W=650.00n L=60.00n
MM0 net038 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net038 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS IOA21HSV2
****Sub-Circuit for IOA21HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT IOA21HSV4 A1 A2 B ZN VDD VSS
MM2 ZN net038 net030 VPW N12LL W=860.00n L=60.00n
MM3 net030 B VSS VPW N12LL W=860.00n L=60.00n
MM1 net038 A1 net18 VPW N12LL W=350.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=350.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=1.3u L=60.00n
MM5 ZN net038 VDD VNW P12LL W=1.3u L=60.00n
MM0 net038 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net038 A1 VDD VNW P12LL W=520.00n L=60.00n
.ENDS IOA21HSV4
****Sub-Circuit for IOA22HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT IOA22HSV0 A1 A2 B1 B2 ZN VDD VSS
MM6 net030 B2 VSS VPW N12LL W=200.00n L=60.00n
MM2 ZN net038 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net038 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN B1 net063 VNW P12LL W=300.00n L=60.00n
MM5 ZN net038 VDD VNW P12LL W=300.00n L=60.00n
MM7 net063 B2 VDD VNW P12LL W=300.00n L=60.00n
MM0 net038 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net038 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS IOA22HSV0
****Sub-Circuit for IOA22HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT IOA22HSV1 A1 A2 B1 B2 ZN VDD VSS
MM6 net030 B2 VSS VPW N12LL W=290.00n L=60.00n
MM2 ZN net038 net030 VPW N12LL W=290.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=290.00n L=60.00n
MM1 net038 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN B1 net063 VNW P12LL W=440.00n L=60.00n
MM5 ZN net038 VDD VNW P12LL W=440.00n L=60.00n
MM7 net063 B2 VDD VNW P12LL W=440.00n L=60.00n
MM0 net038 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net038 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS IOA22HSV1
****Sub-Circuit for IOA22HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT IOA22HSV2 A1 A2 B1 B2 ZN VDD VSS
MM6 net030 B2 VSS VPW N12LL W=430.00n L=60.00n
MM2 ZN net038 net030 VPW N12LL W=430.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=430.00n L=60.00n
MM1 net038 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN B1 net063 VNW P12LL W=650.00n L=60.00n
MM5 ZN net038 VDD VNW P12LL W=650.00n L=60.00n
MM7 net063 B2 VDD VNW P12LL W=650.00n L=60.00n
MM0 net038 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net038 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS IOA22HSV2
****Sub-Circuit for IOA22HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT IOA22HSV4 A1 A2 B1 B2 ZN VDD VSS
MM6 net030 B2 VSS VPW N12LL W=860.00n L=60.00n
MM2 ZN net038 net030 VPW N12LL W=860.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=860.00n L=60.00n
MM1 net038 A1 net18 VPW N12LL W=350.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=350.00n L=60.00n
MM4 ZN B1 net063 VNW P12LL W=1.3u L=60.00n
MM5 ZN net038 VDD VNW P12LL W=1.3u L=60.00n
MM7 net063 B2 VDD VNW P12LL W=1.3u L=60.00n
MM0 net038 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net038 A1 VDD VNW P12LL W=520.00n L=60.00n
.ENDS IOA22HSV4
****Sub-Circuit for LAHHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHHSV1 D E Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c E VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 c pm VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c E VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=400.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHHSV1
****Sub-Circuit for LAHHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHHSV2 D E Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c E VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 c pm VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c E VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=570.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=570.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LAHHSV2
****Sub-Circuit for LAHHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHHSV4 D E Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c E VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 c pm VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c E VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=650.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LAHHSV4
****Sub-Circuit for LAHRNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRNHSV1 D E Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=340.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c E VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=340.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=340.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=600.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c E VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=560.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=560.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHRNHSV1
****Sub-Circuit for LAHRNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRNHSV2 D E Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=410.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=390.00n L=60.00n
MM27 c E VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=410.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c E VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=560.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=560.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHRNHSV2
****Sub-Circuit for LAHRNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRNHSV4 D E Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c E VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c E VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net117 cn pm VNW P12LL W=350.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=350.00n L=60.00n
MM10 pm c net128 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LAHRNHSV4
****Sub-Circuit for LAHRSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRSNHSV1 D E Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=330.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c E VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=330.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=330.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c E VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHRSNHSV1
****Sub-Circuit for LAHRSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHRSNHSV2 D E Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c E VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c E VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LAHRSNHSV2
****Sub-Circuit for LAHRSNHSV4, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT LAHRSNHSV4 D E Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM51 pm s VSS VPW N12LL W=240.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c E VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=360.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=650.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=640.00n L=60.00n
MM28 c E VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net0292 VNW P12LL W=640.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=510.00n L=60.00n
.ENDS LAHRSNHSV4
****Sub-Circuit for LAHSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHSNHSV1 D E Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=290.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c E VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 c net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 cn net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c E VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=430.00n L=60.00n
MM47 Q net0127 VDD VNW P12LL W=430.00n L=60.00n
MM14 net0285 cn net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 c net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=360.00n L=60.00n
.ENDS LAHSNHSV1
****Sub-Circuit for LAHSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHSNHSV2 D E Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=430.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c E VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 c net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 cn net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c E VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q net0127 VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 cn net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 c net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=440.00n L=60.00n
.ENDS LAHSNHSV2
****Sub-Circuit for LAHSNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LAHSNHSV4 D E Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=860.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=405.00n L=60.00n
MM27 c E VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 c net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 cn net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=320.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=650.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c E VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q net0127 VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 cn net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 c net0292 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=510.00n L=60.00n
.ENDS LAHSNHSV4
****Sub-Circuit for LALHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALHSV1 D EN Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c EN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c EN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=400.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALHSV1
****Sub-Circuit for LALHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALHSV2 D EN Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c EN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c EN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=570.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=570.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LALHSV2
****Sub-Circuit for LALHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALHSV4 D EN Q QN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c EN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c EN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net0285 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=650.00n L=60.00n
MM8 net0292 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LALHSV4
****Sub-Circuit for LALRNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRNHSV1 D EN Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=230.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c EN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=230.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=230.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=200.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c EN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS LALRNHSV1
****Sub-Circuit for LALRNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRNHSV2 D EN Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=310.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=390.00n L=60.00n
MM27 c EN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=310.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c EN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net117 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net128 VNW P12LL W=560.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=560.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALRNHSV2
****Sub-Circuit for LALRNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRNHSV4 D EN Q QN RDN VDD VSS
MM46 Q pm VSS VPW N12LL W=860.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=380.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c EN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=350.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=350.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c EN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q pm VDD VNW P12LL W=1.3u L=60.00n
MM14 net117 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net128 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=520.00n L=60.00n
.ENDS LALRNHSV4
****Sub-Circuit for LALRSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRSNHSV1 D EN Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=330.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c EN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=330.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=330.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c EN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALRSNHSV1
****Sub-Circuit for LALRSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALRSNHSV2 D EN Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=430.00n L=60.00n
MM51 pm s VSS VPW N12LL W=200.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=430.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c EN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 cn pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=380.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=550.00n L=60.00n
MM52 pm s net0252 VNW P12LL W=300.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=250.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c EN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS LALRSNHSV2
****Sub-Circuit for LALRSNHSV4, Mon May 30 19:34:53 CST 2011****
.SUBCKT LALRSNHSV4 D EN Q QN RDN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0145 VSS VPW N12LL W=860.00n L=60.00n
MM51 net0145 s VSS VPW N12LL W=200.00n L=60.00n
MM44 net_0104 D VSS VPW N12LL W=360.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c EN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 cn net0145 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 RDN net52 VPW N12LL W=200.00n L=60.00n
MM9 net0145 c net69 VPW N12LL W=420.00n L=60.00n
MM7 net69 RDN net_0104 VPW N12LL W=420.00n L=60.00n
MM0 net_0154 net0145 VSS VPW N12LL W=360.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM52 net0145 s net0252 VNW P12LL W=290.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net0252 RDN VDD VNW P12LL W=290.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=640.00n L=60.00n
MM28 c EN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q net0145 VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 c net0145 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0145 cn net0292 VNW P12LL W=605.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=550.00n L=60.00n
MM1 net_0154 net0145 VDD VNW P12LL W=510.00n L=60.00n
.ENDS LALRSNHSV4
****Sub-Circuit for LALSNHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALSNHSV1 D EN Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q pm VSS VPW N12LL W=290.00n L=60.00n
MM51 pm s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=260.00n L=60.00n
MM27 c EN VSS VPW N12LL W=200.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=290.00n L=60.00n
MM12 net_0119 cn pm VPW N12LL W=200.00n L=60.00n
MM9 pm c net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=290.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=240.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=440.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=390.00n L=60.00n
MM28 c EN VDD VNW P12LL W=300.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=440.00n L=60.00n
MM47 Q pm VDD VNW P12LL W=440.00n L=60.00n
MM14 net0285 c pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm cn net0292 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=360.00n L=60.00n
.ENDS LALSNHSV1
****Sub-Circuit for LALSNHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALSNHSV2 D EN Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=430.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=380.00n L=60.00n
MM27 c EN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=430.00n L=60.00n
MM12 net_0119 cn net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 c net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=290.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=600.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=570.00n L=60.00n
MM28 c EN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=650.00n L=60.00n
MM47 Q net0127 VDD VNW P12LL W=650.00n L=60.00n
MM14 net0285 c net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 cn net0292 VNW P12LL W=600.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=600.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=440.00n L=60.00n
.ENDS LALSNHSV2
****Sub-Circuit for LALSNHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT LALSNHSV4 D EN Q QN SDN VDD VSS
MM48 s SDN VSS VPW N12LL W=200.00n L=60.00n
MM46 Q net0127 VSS VPW N12LL W=860.00n L=60.00n
MM51 net0127 s VSS VPW N12LL W=250.00n L=60.00n
MM42 VSS net_0154 net_0119 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c EN VSS VPW N12LL W=290.00n L=60.00n
MM19 QN net_0154 VSS VPW N12LL W=860.00n L=60.00n
MM12 net_0119 cn net0127 VPW N12LL W=200.00n L=60.00n
MM9 net0127 c net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net0127 VSS VPW N12LL W=320.00n L=60.00n
MM50 net0292 s net128 VNW P12LL W=650.00n L=60.00n
MM49 s SDN VDD VNW P12LL W=300.00n L=60.00n
MM53 net117 s net0285 VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c EN VDD VNW P12LL W=440.00n L=60.00n
MM20 QN net_0154 VDD VNW P12LL W=1.3u L=60.00n
MM47 Q net0127 VDD VNW P12LL W=1.3u L=60.00n
MM14 net0285 c net0127 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net0127 cn net0292 VNW P12LL W=650.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=650.00n L=60.00n
MM1 net_0154 net0127 VDD VNW P12LL W=510.00n L=60.00n
.ENDS LALSNHSV4
****Sub-Circuit for MAJ23HSV0, Mon May 30 14:39:41 CST 2011****
.SUBCKT MAJ23HSV0 A1 A2 A3 Z VDD VSS
MM0 net100 A3 net_8 VNW P12LL W=180.00n L=60.00n
MM1 net_8 A2 VDD VNW P12LL W=260.00n L=60.00n
MM18 net_8 A1 VDD VNW P12LL W=260.00n L=60.00n
MM32 Z net100 VDD VNW P12LL W=250.00n L=60.00n
MM3 net_28 A2 VDD VNW P12LL W=180.00n L=60.00n
MM2 net100 A1 net_28 VNW P12LL W=180.00n L=60.00n
MM35 net_29 A1 VSS VPW N12LL W=220.00n L=60.00n
MM37 net_33 A2 VSS VPW N12LL W=180.00n L=60.00n
MM17 net100 A1 net_33 VPW N12LL W=180.00n L=60.00n
MM31 Z net100 VSS VPW N12LL W=200.00n L=60.00n
MM4 net_29 A2 VSS VPW N12LL W=220.00n L=60.00n
MM5 net100 A3 net_29 VPW N12LL W=180.00n L=60.00n
.ENDS MAJ23HSV0
****Sub-Circuit for MAJ23HSV1, Mon May 30 14:39:41 CST 2011****
.SUBCKT MAJ23HSV1 A1 A2 A3 Z VDD VSS
MM0 net100 A3 net_8 VNW P12LL W=200.00n L=60.00n
MM1 net_8 A2 VDD VNW P12LL W=290.00n L=60.00n
MM18 net_8 A1 VDD VNW P12LL W=290.00n L=60.00n
MM32 Z net100 VDD VNW P12LL W=440.00n L=60.00n
MM3 net_28 A2 VDD VNW P12LL W=200.00n L=60.00n
MM2 net100 A1 net_28 VNW P12LL W=200.00n L=60.00n
MM35 net_29 A1 VSS VPW N12LL W=250.00n L=60.00n
MM37 net_33 A2 VSS VPW N12LL W=180.00n L=60.00n
MM17 net100 A1 net_33 VPW N12LL W=180.00n L=60.00n
MM31 Z net100 VSS VPW N12LL W=350.00n L=60.00n
MM4 net_29 A2 VSS VPW N12LL W=250.00n L=60.00n
MM5 net100 A3 net_29 VPW N12LL W=180.00n L=60.00n
.ENDS MAJ23HSV1
****Sub-Circuit for MAJ23HSV2, Mon Jan 24 15:15:20 CST 2011****
.SUBCKT MAJ23HSV2 A1 A2 A3 Z VDD VSS
MM0 net100 A3 net_8 VNW P12LL W=220.00n L=60.00n
MM1 net_8 A2 VDD VNW P12LL W=350.00n L=60.00n
MM18 net_8 A1 VDD VNW P12LL W=350.00n L=60.00n
MM32 Z net100 VDD VNW P12LL W=540.00n L=60.00n
MM3 net_28 A2 VDD VNW P12LL W=220.00n L=60.00n
MM2 net100 A1 net_28 VNW P12LL W=220.00n L=60.00n
MM35 net_29 A1 VSS VPW N12LL W=320.00n L=60.00n
MM37 net_33 A2 VSS VPW N12LL W=180.00n L=60.00n
MM17 net100 A1 net_33 VPW N12LL W=180.00n L=60.00n
MM31 Z net100 VSS VPW N12LL W=430.00n L=60.00n
MM4 net_29 A2 VSS VPW N12LL W=320.00n L=60.00n
MM5 net100 A3 net_29 VPW N12LL W=180.00n L=60.00n
.ENDS MAJ23HSV2
****Sub-Circuit for MAJ23HSV4, Mon Jan 24 15:15:21 CST 2011****
.SUBCKT MAJ23HSV4 A1 A2 A3 Z VDD VSS
MM0 net100 A3 net_8 VNW P12LL W=440.00n L=60.00n
MM1 net_8 A2 VDD VNW P12LL W=650.00n L=60.00n
MM18 net_8 A1 VDD VNW P12LL W=650.00n L=60.00n
MM32 Z net100 VDD VNW P12LL W=1.08u L=60.00n
MM3 net_28 A2 VDD VNW P12LL W=440.00n L=60.00n
MM2 net100 A1 net_28 VNW P12LL W=440.00n L=60.00n
MM35 net_29 A1 VSS VPW N12LL W=430.00n L=60.00n
MM37 net_33 A2 VSS VPW N12LL W=350.00n L=60.00n
MM17 net100 A1 net_33 VPW N12LL W=350.00n L=60.00n
MM31 Z net100 VSS VPW N12LL W=860.00n L=60.00n
MM4 net_29 A2 VSS VPW N12LL W=430.00n L=60.00n
MM5 net100 A3 net_29 VPW N12LL W=350.00n L=60.00n
.ENDS MAJ23HSV4
****Sub-Circuit for MAOI222HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MAOI222HSV0 A B C ZN VDD VSS
MM6 ZN C net4 VPW N12LL W=200.00n L=60.00n
MM10 net4 B VSS VPW N12LL W=200.00n L=60.00n
MM9 net5 C VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN A net6 VPW N12LL W=200.00n L=60.00n
MM4 ZN A net5 VPW N12LL W=200.00n L=60.00n
MMN1 net6 B VSS VPW N12LL W=200.00n L=60.00n
MM8 net2 C net1 VNW P12LL W=300.0n L=60.00n
MM11 ZN B net2 VNW P12LL W=300.0n L=60.00n
MM7 net1 B VDD VNW P12LL W=300.0n L=60.00n
MM5 net1 C VDD VNW P12LL W=300.0n L=60.00n
MM0 net2 A net1 VNW P12LL W=300.0n L=60.00n
MMP1 ZN A net2 VNW P12LL W=300.0n L=60.00n
.ENDS MAOI222HSV0
****Sub-Circuit for MAOI222HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MAOI222HSV1 A B C ZN VDD VSS
MM6 ZN C net4 VPW N12LL W=290.00n L=60.00n
MM10 net4 B VSS VPW N12LL W=290.00n L=60.00n
MM9 net5 C VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN A net6 VPW N12LL W=290.00n L=60.00n
MM4 ZN A net5 VPW N12LL W=290.00n L=60.00n
MMN1 net6 B VSS VPW N12LL W=290.00n L=60.00n
MM8 net2 C net1 VNW P12LL W=440.0n L=60.00n
MM11 ZN B net2 VNW P12LL W=440.0n L=60.00n
MM7 net1 B VDD VNW P12LL W=440.0n L=60.00n
MM5 net1 C VDD VNW P12LL W=440.0n L=60.00n
MM0 net2 A net1 VNW P12LL W=440.0n L=60.00n
MMP1 ZN A net2 VNW P12LL W=440.0n L=60.00n
.ENDS MAOI222HSV1
****Sub-Circuit for MAOI222HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MAOI222HSV2 A B C ZN VDD VSS
MM6 ZN C net4 VPW N12LL W=430.00n L=60.00n
MM10 net4 B VSS VPW N12LL W=430.00n L=60.00n
MM9 net5 C VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN A net6 VPW N12LL W=430.00n L=60.00n
MM4 ZN A net5 VPW N12LL W=430.00n L=60.00n
MMN1 net6 B VSS VPW N12LL W=430.00n L=60.00n
MM8 net2 C net1 VNW P12LL W=650.0n L=60.00n
MM11 ZN B net2 VNW P12LL W=650.0n L=60.00n
MM7 net1 B VDD VNW P12LL W=650.0n L=60.00n
MM5 net1 C VDD VNW P12LL W=650.0n L=60.00n
MM0 net2 A net1 VNW P12LL W=650.0n L=60.00n
MMP1 ZN A net2 VNW P12LL W=650.0n L=60.00n
.ENDS MAOI222HSV2
****Sub-Circuit for MAOI222HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MAOI222HSV4 A B C ZN VDD VSS
MM6 ZN B net4 VPW N12LL W=860.00n L=60.00n
MM10 net4 C VSS VPW N12LL W=860.00n L=60.00n
MM9 net5 C VSS VPW N12LL W=860.00n L=60.00n
MM1 ZN A net6 VPW N12LL W=860.00n L=60.00n
MM4 ZN A net5 VPW N12LL W=860.00n L=60.00n
MMN1 net6 B VSS VPW N12LL W=860.00n L=60.00n
MM8 net2 C net1 VNW P12LL W=1.3u L=60.00n
MM11 ZN B net2 VNW P12LL W=1.3u L=60.00n
MM7 net1 B VDD VNW P12LL W=1.3u L=60.00n
MM5 net1 C VDD VNW P12LL W=1.3u L=60.00n
MM0 net2 A net1 VNW P12LL W=1.28u L=60.00n
MMP1 ZN A net2 VNW P12LL W=1.3u L=60.00n
.ENDS MAOI222HSV4
****Sub-Circuit for MAOI22HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MAOI22HSV0 A1 A2 B1 B2 ZN VDD VSS
MM3 net24 B2 VSS VPW N12LL W=200.00n L=60.00n
MM2 net24 B1 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN A1 net050 VPW N12LL W=200.00n L=60.00n
MM7 net050 A2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=200.00n L=60.00n
MM6 net061 A2 VDD VNW P12LL W=300.00n L=60.00n
MM4 net24 B2 net074 VNW P12LL W=300.00n L=60.00n
MM5 net074 B1 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net24 net061 VNW P12LL W=300.00n L=60.00n
MMP1 net061 A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS MAOI22HSV0
****Sub-Circuit for MAOI22HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MAOI22HSV1 A1 A2 B1 B2 ZN VDD VSS
MM3 net24 B2 VSS VPW N12LL W=200.00n L=60.00n
MM2 net24 B1 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN A1 net050 VPW N12LL W=290.00n L=60.00n
MM7 net050 A2 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=290.00n L=60.00n
MM6 net061 A2 VDD VNW P12LL W=440.00n L=60.00n
MM4 net24 B2 net074 VNW P12LL W=300.00n L=60.00n
MM5 net074 B1 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net24 net061 VNW P12LL W=440.00n L=60.00n
MMP1 net061 A1 VDD VNW P12LL W=440.00n L=60.00n
.ENDS MAOI22HSV1
****Sub-Circuit for MAOI22HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MAOI22HSV2 A1 A2 B1 B2 ZN VDD VSS
MM3 net24 B2 VSS VPW N12LL W=200.00n L=60.00n
MM2 net24 B1 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN A1 net050 VPW N12LL W=430.00n L=60.00n
MM7 net050 A2 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=430.00n L=60.00n
MM6 net061 A2 VDD VNW P12LL W=650.00n L=60.00n
MM4 net24 B2 net074 VNW P12LL W=300.00n L=60.00n
MM5 net074 B1 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN net24 net061 VNW P12LL W=650.00n L=60.00n
MMP1 net061 A1 VDD VNW P12LL W=650.00n L=60.00n
.ENDS MAOI22HSV2
****Sub-Circuit for MAOI22HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MAOI22HSV4 A1 A2 B1 B2 ZN VDD VSS
MM3 net24 B2 VSS VPW N12LL W=350.0n L=60.00n
MM2 net24 B1 VSS VPW N12LL W=350.0n L=60.00n
MM0 ZN A1 net050 VPW N12LL W=860.00n L=60.00n
MM7 net050 A2 VSS VPW N12LL W=860.00n L=60.00n
MMN1 ZN net24 VSS VPW N12LL W=860.00n L=60.00n
MM6 net061 A2 VDD VNW P12LL W=1.3u L=60.00n
MM4 net24 B2 net074 VNW P12LL W=520.0n L=60.00n
MM5 net074 B1 VDD VNW P12LL W=520.0n L=60.00n
MM1 ZN net24 net061 VNW P12LL W=1.3u L=60.00n
MMP1 net061 A1 VDD VNW P12LL W=1.3u L=60.00n
.ENDS MAOI22HSV4
****Sub-Circuit for MOAI22HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MOAI22HSV0 A1 A2 B1 B2 ZN VDD VSS
MM6 net030 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 ZN net038 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net038 B1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 B2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN A1 net063 VNW P12LL W=300.00n L=60.00n
MM5 ZN net038 VDD VNW P12LL W=300.00n L=60.00n
MM7 net063 A2 VDD VNW P12LL W=300.00n L=60.00n
MM0 net038 B2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net038 B1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS MOAI22HSV0
****Sub-Circuit for MOAI22HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MOAI22HSV1 A1 A2 B1 B2 ZN VDD VSS
MM6 net030 A2 VSS VPW N12LL W=290.00n L=60.00n
MM2 ZN net038 net030 VPW N12LL W=290.00n L=60.00n
MM3 net030 A1 VSS VPW N12LL W=290.00n L=60.00n
MM1 net038 B1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 B2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN A1 net063 VNW P12LL W=440.00n L=60.00n
MM5 ZN net038 VDD VNW P12LL W=440.00n L=60.00n
MM7 net063 A2 VDD VNW P12LL W=440.00n L=60.00n
MM0 net038 B2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net038 B1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS MOAI22HSV1
****Sub-Circuit for MOAI22HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MOAI22HSV2 A1 A2 B1 B2 ZN VDD VSS
MM6 net030 A2 VSS VPW N12LL W=430.00n L=60.00n
MM2 ZN net038 net030 VPW N12LL W=430.00n L=60.00n
MM3 net030 A1 VSS VPW N12LL W=430.00n L=60.00n
MM1 net038 B1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 B2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN A1 net063 VNW P12LL W=650.00n L=60.00n
MM5 ZN net038 VDD VNW P12LL W=650.00n L=60.00n
MM7 net063 A2 VDD VNW P12LL W=650.00n L=60.00n
MM0 net038 B2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net038 B1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS MOAI22HSV2
****Sub-Circuit for MOAI22HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MOAI22HSV4 A1 A2 B1 B2 ZN VDD VSS
MM6 net030 A2 VSS VPW N12LL W=860.00n L=60.00n
MM2 ZN net038 net030 VPW N12LL W=860.00n L=60.00n
MM3 net030 A1 VSS VPW N12LL W=860.00n L=60.00n
MM1 net038 B1 net18 VPW N12LL W=350.00n L=60.00n
MMN1 net18 B2 VSS VPW N12LL W=350.00n L=60.00n
MM4 ZN A1 net063 VNW P12LL W=1.3u L=60.00n
MM5 ZN net038 VDD VNW P12LL W=1.3u L=60.00n
MM7 net063 A2 VDD VNW P12LL W=1.3u L=60.00n
MM0 net038 B2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net038 B1 VDD VNW P12LL W=520.00n L=60.00n
.ENDS MOAI22HSV4
****Sub-Circuit for MUX2HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX2HSV0 I0 I1 S Z VDD VSS
MM47 net41 S net64 VPW N12LL W=200.00n L=60.00n
MM51 Z net64 VSS VPW N12LL W=200.00n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=200.00n L=60.00n
MM31 net41 I1 VSS VPW N12LL W=200.00n L=60.00n
MM53 net43 S VSS VPW N12LL W=200.00n L=60.00n
MM36 net39 net43 net64 VPW N12LL W=200.00n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=300.0n L=60.00n
MM52 Z net64 VDD VNW P12LL W=300.0n L=60.00n
MM48 net41 net43 net64 VNW P12LL W=300.00n L=60.00n
MM32 net41 I1 VDD VNW P12LL W=300.0n L=60.00n
MM54 net43 S VDD VNW P12LL W=300.00n L=60.00n
MM39 net39 S net64 VNW P12LL W=300.00n L=60.00n
.ENDS MUX2HSV0
****Sub-Circuit for MUX2HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX2HSV1 I0 I1 S Z VDD VSS
MM47 net41 S net64 VPW N12LL W=200.00n L=60.00n
MM51 Z net64 VSS VPW N12LL W=290.00n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=200.00n L=60.00n
MM31 net41 I1 VSS VPW N12LL W=200.00n L=60.00n
MM53 net43 S VSS VPW N12LL W=200.00n L=60.00n
MM36 net39 net43 net64 VPW N12LL W=200.00n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=300.0n L=60.00n
MM52 Z net64 VDD VNW P12LL W=440.0n L=60.00n
MM48 net41 net43 net64 VNW P12LL W=300.00n L=60.00n
MM32 net41 I1 VDD VNW P12LL W=300.0n L=60.00n
MM54 net43 S VDD VNW P12LL W=300.00n L=60.00n
MM39 net39 S net64 VNW P12LL W=300.00n L=60.00n
.ENDS MUX2HSV1
****Sub-Circuit for MUX2HSV2, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT MUX2HSV2 I0 I1 S Z VDD VSS
MM47 net41 S net64 VPW N12LL W=290.00n L=60.00n
MM51 Z net64 VSS VPW N12LL W=430.00n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=290.00n L=60.00n
MM31 net41 I1 VSS VPW N12LL W=290.00n L=60.00n
MM53 net43 S VSS VPW N12LL W=200.00n L=60.00n
MM36 net39 net43 net64 VPW N12LL W=290.00n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=410.00n L=60.00n
MM52 Z net64 VDD VNW P12LL W=650.0n L=60.00n
MM48 net41 net43 net64 VNW P12LL W=440.00n L=60.00n
MM32 net41 I1 VDD VNW P12LL W=440.00n L=60.00n
MM54 net43 S VDD VNW P12LL W=300.00n L=60.00n
MM39 net39 S net64 VNW P12LL W=440.00n L=60.00n
.ENDS MUX2HSV2
****Sub-Circuit for MUX2HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX2HSV4 I0 I1 S Z VDD VSS
MM47 net41 S net64 VPW N12LL W=600.00n L=60.00n
MM51 Z net64 VSS VPW N12LL W=860.00n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=570.00n L=60.00n
MM31 net41 I1 VSS VPW N12LL W=570.00n L=60.00n
MM53 net43 S VSS VPW N12LL W=430.00n L=60.00n
MM36 net39 net43 net64 VPW N12LL W=600.00n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=870.0n L=60.00n
MM52 Z net64 VDD VNW P12LL W=1.3u L=60.00n
MM48 net41 net43 net64 VNW P12LL W=870.0n L=60.00n
MM32 net41 I1 VDD VNW P12LL W=870.0n L=60.00n
MM54 net43 S VDD VNW P12LL W=650.000n L=60.00n
MM39 net39 S net64 VNW P12LL W=870.0n L=60.00n
.ENDS MUX2HSV4
****Sub-Circuit for MUX2NHSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX2NHSV0 I0 I1 S ZN VDD VSS
MM47 net41 S ZN VPW N12LL W=200.0n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=200.0n L=60.00n
MM31 net41 I1 VSS VPW N12LL W=200.0n L=60.00n
MM53 net43 S VSS VPW N12LL W=200.00n L=60.00n
MM36 net39 net43 ZN VPW N12LL W=200.0n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=300.00n L=60.00n
MM48 net41 net43 ZN VNW P12LL W=300.00n L=60.00n
MM32 net41 I1 VDD VNW P12LL W=300.00n L=60.00n
MM54 net43 S VDD VNW P12LL W=300.00n L=60.00n
MM39 net39 S ZN VNW P12LL W=300.00n L=60.00n
.ENDS MUX2NHSV0
****Sub-Circuit for MUX2NHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX2NHSV1 I0 I1 S ZN VDD VSS
MM47 net41 S ZN VPW N12LL W=290.0n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=290.0n L=60.00n
MM31 net41 I1 VSS VPW N12LL W=290.0n L=60.00n
MM53 net43 S VSS VPW N12LL W=200.00n L=60.00n
MM36 net39 net43 ZN VPW N12LL W=290.0n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=440.00n L=60.00n
MM48 net41 net43 ZN VNW P12LL W=440.00n L=60.00n
MM32 net41 I1 VDD VNW P12LL W=440.00n L=60.00n
MM54 net43 S VDD VNW P12LL W=300.00n L=60.00n
MM39 net39 S ZN VNW P12LL W=440.00n L=60.00n
.ENDS MUX2NHSV1
****Sub-Circuit for MUX2NHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX2NHSV2 I0 I1 S ZN VDD VSS
MM47 net41 S ZN VPW N12LL W=430.0n L=60.00n
MM49 net39 I0 VSS VPW N12LL W=430.0n L=60.00n
MM31 net41 I1 VSS VPW N12LL W=430.0n L=60.00n
MM53 net43 S VSS VPW N12LL W=290.00n L=60.00n
MM36 net39 net43 ZN VPW N12LL W=430.0n L=60.00n
MM50 net39 I0 VDD VNW P12LL W=650.00n L=60.00n
MM48 net41 net43 ZN VNW P12LL W=565.00n L=60.00n
MM32 net41 I1 VDD VNW P12LL W=650.00n L=60.00n
MM54 net43 S VDD VNW P12LL W=440.00n L=60.00n
MM39 net39 S ZN VNW P12LL W=640.00n L=60.00n
.ENDS MUX2NHSV2
****Sub-Circuit for MUX2NHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX2NHSV4 I0 I1 S ZN VDD VSS
MM2 net_045 I1 VSS VPW N12LL W=860.00n L=60.00n
MM47 net_045 S ZN VPW N12LL W=780.00n L=60.00n
MM0 net_041 I0 VSS VPW N12LL W=860.00n L=60.00n
MM53 net43 S VSS VPW N12LL W=430.00n L=60.00n
MM36 net_041 net43 ZN VPW N12LL W=780.00n L=60.00n
MM48 net_045 net43 ZN VNW P12LL W=970n L=60.00n
MM3 net_045 I1 VDD VNW P12LL W=1.1u L=60.00n
MM1 net_041 I0 VDD VNW P12LL W=1.1u L=60.00n
MM54 net43 S VDD VNW P12LL W=550n L=60.00n
MM39 net_041 S ZN VNW P12LL W=970n L=60.00n
.ENDS MUX2NHSV4
****Sub-Circuit for MUX3HSV0, Mon May 30 14:11:46 CST 2011****
.SUBCKT MUX3HSV0 I0 I1 I2 S0 S1 Z VDD VSS
MM2 S0N S0 VDD VNW P12LL W=250.00n L=60.00n
MM0 net67 I1 VDD VNW P12LL W=250.00n L=60.00n
MM39 net75 S0 net82 VNW P12LL W=250.00n L=60.00n
MM56 net75 I0 VDD VNW P12LL W=250.00n L=60.00n
MM48 net67 S0N net82 VNW P12LL W=250.00n L=60.00n
MM58 Z net54 VDD VNW P12LL W=250.00n L=60.00n
MM5 S1N S1 VDD VNW P12LL W=250.00n L=60.00n
MM7 net59 I2 VDD VNW P12LL W=250.00n L=60.00n
MM9 net59 S1N net54 VNW P12LL W=250.00n L=60.00n
MM13 net82 S1 net54 VNW P12LL W=250.00n L=60.00n
MM6 net59 I2 VSS VPW N12LL W=200.00n L=60.00n
MM3 S0N S0 VSS VPW N12LL W=200.00n L=60.00n
MM1 net67 I1 VSS VPW N12LL W=200.00n L=60.00n
MM36 net75 S0N net82 VPW N12LL W=200.00n L=60.00n
MM55 net75 I0 VSS VPW N12LL W=200.00n L=60.00n
MM47 net67 S0 net82 VPW N12LL W=200.00n L=60.00n
MM57 Z net54 VSS VPW N12LL W=200.00n L=60.00n
MM4 S1N S1 VSS VPW N12LL W=200.00n L=60.00n
MM8 net59 S1 net54 VPW N12LL W=200.00n L=60.00n
MM12 net82 S1N net54 VPW N12LL W=200.00n L=60.00n
.ENDS MUX3HSV0
****Sub-Circuit for MUX3HSV1, Mon May 30 14:11:46 CST 2011****
.SUBCKT MUX3HSV1 I0 I1 I2 S0 S1 Z VDD VSS
MM12 net26 S1N net14 VPW N12LL W=230.00n L=60.00n
MM8 net43 S1 net14 VPW N12LL W=230.00n L=60.00n
MM4 S1N S1 VSS VPW N12LL W=230.00n L=60.00n
MM57 Z net14 VSS VPW N12LL W=350.00n L=60.00n
MM47 net35 S0 net26 VPW N12LL W=230.00n L=60.00n
MM55 net27 I0 VSS VPW N12LL W=230.00n L=60.00n
MM36 net27 S0N net26 VPW N12LL W=230.00n L=60.00n
MM1 net35 I1 VSS VPW N12LL W=230.00n L=60.00n
MM3 S0N S0 VSS VPW N12LL W=230.00n L=60.00n
MM6 net43 I2 VSS VPW N12LL W=230.00n L=60.00n
MM13 net26 S1 net14 VNW P12LL W=290.00n L=60.00n
MM9 net43 S1N net14 VNW P12LL W=290.00n L=60.00n
MM7 net43 I2 VDD VNW P12LL W=290.00n L=60.00n
MM5 S1N S1 VDD VNW P12LL W=290.00n L=60.00n
MM58 Z net14 VDD VNW P12LL W=440.00n L=60.00n
MM48 net35 S0N net26 VNW P12LL W=290.00n L=60.00n
MM56 net27 I0 VDD VNW P12LL W=290.00n L=60.00n
MM39 net27 S0 net26 VNW P12LL W=290.00n L=60.00n
MM0 net35 I1 VDD VNW P12LL W=290.00n L=60.00n
MM2 S0N S0 VDD VNW P12LL W=290.00n L=60.00n
.ENDS MUX3HSV1
****Sub-Circuit for MUX3HSV2, Mon May 30 14:11:46 CST 2011****
.SUBCKT MUX3HSV2 I0 I1 I2 S0 S1 Z VDD VSS
MM12 net26 S1N net14 VPW N12LL W=290.00n L=60.00n
MM8 net43 S1 net14 VPW N12LL W=290.00n L=60.00n
MM4 S1N S1 VSS VPW N12LL W=290.00n L=60.00n
MM57 Z net14 VSS VPW N12LL W=430.00n L=60.00n
MM47 net35 S0 net26 VPW N12LL W=290.00n L=60.00n
MM55 net27 I0 VSS VPW N12LL W=290.00n L=60.00n
MM36 net27 S0N net26 VPW N12LL W=290.00n L=60.00n
MM1 net35 I1 VSS VPW N12LL W=290.00n L=60.00n
MM3 S0N S0 VSS VPW N12LL W=290.00n L=60.00n
MM6 net43 I2 VSS VPW N12LL W=290.00n L=60.00n
MM13 net26 S1 net14 VNW P12LL W=360.00n L=60.00n
MM9 net43 S1N net14 VNW P12LL W=360.00n L=60.00n
MM7 net43 I2 VDD VNW P12LL W=360.00n L=60.00n
MM5 S1N S1 VDD VNW P12LL W=360.00n L=60.00n
MM58 Z net14 VDD VNW P12LL W=540.00n L=60.00n
MM48 net35 S0N net26 VNW P12LL W=360.00n L=60.00n
MM56 net27 I0 VDD VNW P12LL W=360.00n L=60.00n
MM39 net27 S0 net26 VNW P12LL W=360.00n L=60.00n
MM0 net35 I1 VDD VNW P12LL W=360.00n L=60.00n
MM2 S0N S0 VDD VNW P12LL W=360.00n L=60.00n
.ENDS MUX3HSV2
****Sub-Circuit for MUX3HSV4, Mon May 30 14:26:44 CST 2011****
.SUBCKT MUX3HSV4 I0 I1 I2 S0 S1 Z VDD VSS
MM55 net99 S1 net73 VPW N12LL W=430.00n L=60.00n
MM58 net61 net111 net73 VPW N12LL W=570.00n L=60.00n
MM47 net97 S0 net61 VPW N12LL W=570.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=570.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=290.00n L=60.00n
MM67 net99 I2 VSS VPW N12LL W=430.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=570.00n L=60.00n
MM69 Z net73 VSS VPW N12LL W=860.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=430.00n L=60.00n
MM36 net95 net107 net61 VPW N12LL W=570.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=860.00n L=60.00n
MM60 net99 net111 net73 VNW P12LL W=640.00n L=60.00n
MM62 net61 S1 net73 VNW P12LL W=870.00n L=60.00n
MM48 net97 net107 net61 VNW P12LL W=860.00n L=60.00n
MM70 Z net73 VDD VNW P12LL W=1.3u L=60.00n
MM66 net111 S1 VDD VNW P12LL W=440.00n L=60.00n
MM68 net99 I2 VDD VNW P12LL W=650.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=860.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=605.00n L=60.00n
MM39 net95 S0 net61 VNW P12LL W=860.00n L=60.00n
.ENDS MUX3HSV4
****Sub-Circuit for MUX3NHSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX3NHSV0 I0 I1 I2 S0 S1 ZN VDD VSS
MM55 net105 S1 net73 VPW N12LL W=200.00n L=60.00n
MM56 net103 net61 VSS VPW N12LL W=200.00n L=60.00n
MM57 net105 net99 VSS VPW N12LL W=200.00n L=60.00n
MM58 net103 net111 net73 VPW N12LL W=200.00n L=60.00n
MM47 net97 S0 net61 VPW N12LL W=200.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=200.00n L=60.00n
MM63 ZN net73 VSS VPW N12LL W=200.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=200.00n L=60.00n
MM67 net99 I2 VSS VPW N12LL W=200.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=200.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=200.00n L=60.00n
MM36 net95 net107 net61 VPW N12LL W=200.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=300.00n L=60.00n
MM59 net103 net61 VDD VNW P12LL W=300.00n L=60.00n
MM60 net105 net111 net73 VNW P12LL W=300.00n L=60.00n
MM61 net105 net99 VDD VNW P12LL W=300.00n L=60.00n
MM62 net103 S1 net73 VNW P12LL W=300.00n L=60.00n
MM48 net97 net107 net61 VNW P12LL W=300.00n L=60.00n
MM64 ZN net73 VDD VNW P12LL W=300.00n L=60.00n
MM66 net111 S1 VDD VNW P12LL W=300.00n L=60.00n
MM68 net99 I2 VDD VNW P12LL W=300.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=300.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=300.00n L=60.00n
MM39 net95 S0 net61 VNW P12LL W=300.00n L=60.00n
.ENDS MUX3NHSV0
****Sub-Circuit for MUX3NHSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX3NHSV1 I0 I1 I2 S0 S1 ZN VDD VSS
MM55 net105 S1 net73 VPW N12LL W=290.00n L=60.00n
MM56 net103 net61 VSS VPW N12LL W=290.00n L=60.00n
MM57 net105 net99 VSS VPW N12LL W=290.00n L=60.00n
MM58 net103 net111 net73 VPW N12LL W=290.00n L=60.00n
MM47 net97 S0 net61 VPW N12LL W=290.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=290.00n L=60.00n
MM63 ZN net73 VSS VPW N12LL W=290.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=200.00n L=60.00n
MM67 net99 I2 VSS VPW N12LL W=200.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=290.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=200.00n L=60.00n
MM36 net95 net107 net61 VPW N12LL W=290.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=440.00n L=60.00n
MM59 net103 net61 VDD VNW P12LL W=440.00n L=60.00n
MM60 net105 net111 net73 VNW P12LL W=440.00n L=60.00n
MM61 net105 net99 VDD VNW P12LL W=440.00n L=60.00n
MM62 net103 S1 net73 VNW P12LL W=440.00n L=60.00n
MM48 net97 net107 net61 VNW P12LL W=440.00n L=60.00n
MM64 ZN net73 VDD VNW P12LL W=440.00n L=60.00n
MM66 net111 S1 VDD VNW P12LL W=300.00n L=60.00n
MM68 net99 I2 VDD VNW P12LL W=300.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=440.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=300.00n L=60.00n
MM39 net95 S0 net61 VNW P12LL W=440.00n L=60.00n
.ENDS MUX3NHSV1
****Sub-Circuit for MUX3NHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX3NHSV2 I0 I1 I2 S0 S1 ZN VDD VSS
MM55 net105 S1 net73 VPW N12LL W=290.00n L=60.00n
MM56 net103 net61 VSS VPW N12LL W=290.00n L=60.00n
MM57 net105 net99 VSS VPW N12LL W=290.00n L=60.00n
MM58 net103 net111 net73 VPW N12LL W=290.00n L=60.00n
MM47 net97 S0 net61 VPW N12LL W=290.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=290.00n L=60.00n
MM63 ZN net73 VSS VPW N12LL W=430.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=200.00n L=60.00n
MM67 net99 I2 VSS VPW N12LL W=200.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=290.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=290.00n L=60.00n
MM36 net95 net107 net61 VPW N12LL W=290.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=440.00n L=60.00n
MM59 net103 net61 VDD VNW P12LL W=440.00n L=60.00n
MM60 net105 net111 net73 VNW P12LL W=440.00n L=60.00n
MM61 net105 net99 VDD VNW P12LL W=440.00n L=60.00n
MM62 net103 S1 net73 VNW P12LL W=440.00n L=60.00n
MM48 net97 net107 net61 VNW P12LL W=440.00n L=60.00n
MM64 ZN net73 VDD VNW P12LL W=650.00n L=60.00n
MM66 net111 S1 VDD VNW P12LL W=300.00n L=60.00n
MM68 net99 I2 VDD VNW P12LL W=300.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=440.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=440.00n L=60.00n
MM39 net95 S0 net61 VNW P12LL W=440.00n L=60.00n
.ENDS MUX3NHSV2
****Sub-Circuit for MUX3NHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX3NHSV4 I0 I1 I2 S0 S1 ZN VDD VSS
MM55 net105 S1 net73 VPW N12LL W=570.00n L=60.00n
MM56 net103 net61 VSS VPW N12LL W=570.00n L=60.00n
MM57 net105 net99 VSS VPW N12LL W=570.00n L=60.00n
MM58 net103 net111 net73 VPW N12LL W=570.00n L=60.00n
MM47 net97 S0 net61 VPW N12LL W=430.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=430.00n L=60.00n
MM63 ZN net73 VSS VPW N12LL W=860.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=430.00n L=60.00n
MM67 net99 I2 VSS VPW N12LL W=380.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=430.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=430.00n L=60.00n
MM36 net95 net107 net61 VPW N12LL W=430.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=650.00n L=60.00n
MM59 net103 net61 VDD VNW P12LL W=870.00n L=60.00n
MM60 net105 net111 net73 VNW P12LL W=870.00n L=60.00n
MM61 net105 net99 VDD VNW P12LL W=870.00n L=60.00n
MM62 net103 S1 net73 VNW P12LL W=870.00n L=60.00n
MM48 net97 net107 net61 VNW P12LL W=650.00n L=60.00n
MM64 ZN net73 VDD VNW P12LL W=1.3u L=60.00n
MM66 net111 S1 VDD VNW P12LL W=650.00n L=60.00n
MM68 net99 I2 VDD VNW P12LL W=570.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=650.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=650.00n L=60.00n
MM39 net95 S0 net61 VNW P12LL W=650.00n L=60.00n
.ENDS MUX3NHSV4
****Sub-Circuit for MUX4HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX4HSV0 I0 I1 I2 I3 S0 S1 Z VDD VSS
MM58 net59 net111 net71 VPW N12LL W=200.00n L=60.00n
MM47 net97 S0 net59 VPW N12LL W=200.00n L=60.00n
MM69 net65 S1 net71 VPW N12LL W=200.00n L=60.00n
MM70 net101 S0 net65 VPW N12LL W=200.00n L=60.00n
MM72 net101 I3 VSS VPW N12LL W=200.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=200.00n L=60.00n
MM73 net99 net107 net65 VPW N12LL W=200.00n L=60.00n
MM63 Z net71 VSS VPW N12LL W=200.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=200.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=200.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=200.00n L=60.00n
MM71 net99 I2 VSS VPW N12LL W=200.00n L=60.00n
MM36 net95 net107 net59 VPW N12LL W=200.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=300.00n L=60.00n
MM62 net59 S1 net71 VNW P12LL W=300.00n L=60.00n
MM48 net97 net107 net59 VNW P12LL W=300.00n L=60.00n
MM74 net99 I2 VDD VNW P12LL W=300.00n L=60.00n
MM76 net65 net111 net71 VNW P12LL W=300.00n L=60.00n
MM77 net101 net107 net65 VNW P12LL W=300.00n L=60.00n
MM78 net101 I3 VDD VNW P12LL W=300.00n L=60.00n
MM79 net99 S0 net65 VNW P12LL W=300.00n L=60.00n
MM64 Z net71 VDD VNW P12LL W=300.00n L=60.00n
MM66 net111 S1 VDD VNW P12LL W=300.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=300.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=300.00n L=60.00n
MM39 net95 S0 net59 VNW P12LL W=300.00n L=60.00n
.ENDS MUX4HSV0
****Sub-Circuit for MUX4HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX4HSV1 I0 I1 I2 I3 S0 S1 Z VDD VSS
MM58 net59 net111 net71 VPW N12LL W=290.00n L=60.00n
MM47 net97 S0 net59 VPW N12LL W=290.00n L=60.00n
MM69 net65 S1 net71 VPW N12LL W=290.00n L=60.00n
MM70 net101 S0 net65 VPW N12LL W=290.00n L=60.00n
MM72 net101 I3 VSS VPW N12LL W=290.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=290.00n L=60.00n
MM73 net99 net107 net65 VPW N12LL W=290.00n L=60.00n
MM63 Z net71 VSS VPW N12LL W=290.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=290.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=290.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=430.00n L=60.00n
MM71 net99 I2 VSS VPW N12LL W=290.00n L=60.00n
MM36 net95 net107 net59 VPW N12LL W=290.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=440.00n L=60.00n
MM62 net59 S1 net71 VNW P12LL W=440.00n L=60.00n
MM48 net97 net107 net59 VNW P12LL W=440.00n L=60.00n
MM74 net99 I2 VDD VNW P12LL W=440.00n L=60.00n
MM76 net65 net111 net71 VNW P12LL W=440.00n L=60.00n
MM77 net101 net107 net65 VNW P12LL W=440.00n L=60.00n
MM78 net101 I3 VDD VNW P12LL W=440.00n L=60.00n
MM79 net99 S0 net65 VNW P12LL W=440.00n L=60.00n
MM64 Z net71 VDD VNW P12LL W=440.00n L=60.00n
MM66 net111 S1 VDD VNW P12LL W=440.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=440.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=650.00n L=60.00n
MM39 net95 S0 net59 VNW P12LL W=440.00n L=60.00n
.ENDS MUX4HSV1
****Sub-Circuit for MUX4HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX4HSV2 I0 I1 I2 I3 S0 S1 Z VDD VSS
MM58 net59 net111 net71 VPW N12LL W=290.00n L=60.00n
MM47 net97 S0 net59 VPW N12LL W=290.00n L=60.00n
MM69 net65 S1 net71 VPW N12LL W=290.00n L=60.00n
MM70 net101 S0 net65 VPW N12LL W=290.00n L=60.00n
MM72 net101 I3 VSS VPW N12LL W=290.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=290.00n L=60.00n
MM73 net99 net107 net65 VPW N12LL W=290.00n L=60.00n
MM63 Z net71 VSS VPW N12LL W=430.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=290.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=290.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=430.00n L=60.00n
MM71 net99 I2 VSS VPW N12LL W=290.00n L=60.00n
MM36 net95 net107 net59 VPW N12LL W=290.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=440.00n L=60.00n
MM62 net59 S1 net71 VNW P12LL W=440.00n L=60.00n
MM48 net97 net107 net59 VNW P12LL W=440.00n L=60.00n
MM74 net99 I2 VDD VNW P12LL W=440.00n L=60.00n
MM76 net65 net111 net71 VNW P12LL W=440.00n L=60.00n
MM77 net101 net107 net65 VNW P12LL W=440.00n L=60.00n
MM78 net101 I3 VDD VNW P12LL W=440.00n L=60.00n
MM79 net99 S0 net65 VNW P12LL W=440.00n L=60.00n
MM64 Z net71 VDD VNW P12LL W=650.00n L=60.00n
MM66 net111 S1 VDD VNW P12LL W=440.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=440.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=650.00n L=60.00n
MM39 net95 S0 net59 VNW P12LL W=440.00n L=60.00n
.ENDS MUX4HSV2
****Sub-Circuit for MUX4HSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX4HSV4 I0 I1 I2 I3 S0 S1 Z VDD VSS
MM58 net59 net111 net71 VPW N12LL W=430.00n L=60.00n
MM47 net97 S0 net59 VPW N12LL W=430.00n L=60.00n
MM69 net65 S1 net71 VPW N12LL W=430.00n L=60.00n
MM70 net101 S0 net65 VPW N12LL W=430.00n L=60.00n
MM72 net101 I3 VSS VPW N12LL W=430.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=430.00n L=60.00n
MM73 net99 net107 net65 VPW N12LL W=430.00n L=60.00n
MM63 Z net71 VSS VPW N12LL W=860.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=430.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=430.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=570.00n L=60.00n
MM71 net99 I2 VSS VPW N12LL W=430.00n L=60.00n
MM36 net95 net107 net59 VPW N12LL W=430.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=635.00n L=60.00n
MM62 net59 S1 net71 VNW P12LL W=640.00n L=60.00n
MM48 net97 net107 net59 VNW P12LL W=635.00n L=60.00n
MM74 net99 I2 VDD VNW P12LL W=640.00n L=60.00n
MM76 net65 net111 net71 VNW P12LL W=640.00n L=60.00n
MM77 net101 net107 net65 VNW P12LL W=640.00n L=60.00n
MM78 net101 I3 VDD VNW P12LL W=640.00n L=60.00n
MM79 net99 S0 net65 VNW P12LL W=640.00n L=60.00n
MM64 Z net71 VDD VNW P12LL W=1.3u L=60.00n
MM66 net111 S1 VDD VNW P12LL W=650.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=630.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=870.00n L=60.00n
MM39 net95 S0 net59 VNW P12LL W=635.00n L=60.00n
.ENDS MUX4HSV4
****Sub-Circuit for MUX4NHSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX4NHSV0 I0 I1 I2 I3 S0 S1 ZN VDD VSS
MM82 net105 net67 VSS VPW N12LL W=200.00n L=60.00n
MM75 net103 net61 VSS VPW N12LL W=200.00n L=60.00n
MM58 net103 net111 net73 VPW N12LL W=200.00n L=60.00n
MM47 net97 S0 net61 VPW N12LL W=200.00n L=60.00n
MM69 net105 S1 net73 VPW N12LL W=200.00n L=60.00n
MM70 net101 S0 net67 VPW N12LL W=200.00n L=60.00n
MM72 net101 I3 VSS VPW N12LL W=200.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=200.00n L=60.00n
MM73 net99 net107 net67 VPW N12LL W=200.00n L=60.00n
MM63 ZN net73 VSS VPW N12LL W=200.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=200.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=200.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=200.00n L=60.00n
MM71 net99 I2 VSS VPW N12LL W=200.00n L=60.00n
MM36 net95 net107 net61 VPW N12LL W=200.00n L=60.00n
MM81 net105 net67 VDD VNW P12LL W=300.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=300.00n L=60.00n
MM62 net103 S1 net73 VNW P12LL W=300.00n L=60.00n
MM48 net97 net107 net61 VNW P12LL W=300.00n L=60.00n
MM74 net99 I2 VDD VNW P12LL W=300.00n L=60.00n
MM76 net105 net111 net73 VNW P12LL W=300.00n L=60.00n
MM77 net101 net107 net67 VNW P12LL W=300.00n L=60.00n
MM78 net101 I3 VDD VNW P12LL W=300.00n L=60.00n
MM79 net99 S0 net67 VNW P12LL W=300.00n L=60.00n
MM64 ZN net73 VDD VNW P12LL W=300.00n L=60.00n
MM66 net111 S1 VDD VNW P12LL W=300.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=300.00n L=60.00n
MM80 net103 net61 VDD VNW P12LL W=300.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=300.00n L=60.00n
MM39 net95 S0 net61 VNW P12LL W=300.00n L=60.00n
.ENDS MUX4NHSV0
****Sub-Circuit for MUX4NHSV1, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT MUX4NHSV1 I0 I1 I2 I3 S0 S1 ZN VDD VSS
MM82 net105 net67 VSS VPW N12LL W=280.00n L=60.00n
MM75 net103 net61 VSS VPW N12LL W=290.00n L=60.00n
MM58 net103 net111 net73 VPW N12LL W=290.00n L=60.00n
MM47 net97 S0 net61 VPW N12LL W=200.00n L=60.00n
MM69 net105 S1 net73 VPW N12LL W=290.00n L=60.00n
MM70 net101 S0 net67 VPW N12LL W=200.00n L=60.00n
MM72 net101 I3 VSS VPW N12LL W=200.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=200.00n L=60.00n
MM73 net99 net107 net67 VPW N12LL W=200.00n L=60.00n
MM63 ZN net73 VSS VPW N12LL W=290.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=200.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=200.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=290.00n L=60.00n
MM71 net99 I2 VSS VPW N12LL W=200.00n L=60.00n
MM36 net95 net107 net61 VPW N12LL W=200.00n L=60.00n
MM81 net105 net67 VDD VNW P12LL W=420.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=300.00n L=60.00n
MM62 net103 S1 net73 VNW P12LL W=430.00n L=60.00n
MM48 net97 net107 net61 VNW P12LL W=300.00n L=60.00n
MM74 net99 I2 VDD VNW P12LL W=300.00n L=60.00n
MM76 net105 net111 net73 VNW P12LL W=410.00n L=60.00n
MM77 net101 net107 net67 VNW P12LL W=300.00n L=60.00n
MM78 net101 I3 VDD VNW P12LL W=300.00n L=60.00n
MM79 net99 S0 net67 VNW P12LL W=300.00n L=60.00n
MM64 ZN net73 VDD VNW P12LL W=440.00n L=60.00n
MM66 net111 S1 VDD VNW P12LL W=300.00n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=300.00n L=60.00n
MM80 net103 net61 VDD VNW P12LL W=430.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=440.00n L=60.00n
MM39 net95 S0 net61 VNW P12LL W=300.00n L=60.00n
.ENDS MUX4NHSV1
****Sub-Circuit for MUX4NHSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX4NHSV2 I0 I1 I2 I3 S0 S1 ZN VDD VSS
MM82 net105 net67 VSS VPW N12LL W=430.00n L=60.00n
MM75 net103 net61 VSS VPW N12LL W=430.00n L=60.00n
MM58 net103 net111 net73 VPW N12LL W=430.00n L=60.00n
MM47 net97 S0 net61 VPW N12LL W=290.00n L=60.00n
MM69 net105 S1 net73 VPW N12LL W=430.00n L=60.00n
MM70 net101 S0 net67 VPW N12LL W=290.00n L=60.00n
MM72 net101 I3 VSS VPW N12LL W=290.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=290.00n L=60.00n
MM73 net99 net107 net67 VPW N12LL W=290.00n L=60.00n
MM63 ZN net73 VSS VPW N12LL W=430.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=290.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=290.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=430.00n L=60.00n
MM71 net99 I2 VSS VPW N12LL W=290.00n L=60.00n
MM36 net95 net107 net61 VPW N12LL W=290.00n L=60.00n
MM81 net105 net67 VDD VNW P12LL W=640.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=440.00n L=60.00n
MM62 net103 S1 net73 VNW P12LL W=650.00n L=60.00n
MM48 net97 net107 net61 VNW P12LL W=440.00n L=60.00n
MM74 net99 I2 VDD VNW P12LL W=440.00n L=60.00n
MM76 net105 net111 net73 VNW P12LL W=650.00n L=60.00n
MM77 net101 net107 net67 VNW P12LL W=440.00n L=60.00n
MM78 net101 I3 VDD VNW P12LL W=440.00n L=60.00n
MM79 net99 S0 net67 VNW P12LL W=440.00n L=60.00n
MM64 ZN net73 VDD VNW P12LL W=650.00n L=60.00n
MM66 net111 S1 VDD VNW P12LL W=440.0n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=440.00n L=60.00n
MM80 net103 net61 VDD VNW P12LL W=650.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=650.00n L=60.00n
MM39 net95 S0 net61 VNW P12LL W=440.00n L=60.00n
.ENDS MUX4NHSV2
****Sub-Circuit for MUX4NHSV4, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT MUX4NHSV4 I0 I1 I2 I3 S0 S1 ZN VDD VSS
MM82 net105 net67 VSS VPW N12LL W=570.00n L=60.00n
MM75 net103 net61 VSS VPW N12LL W=570.00n L=60.00n
MM58 net103 net111 net73 VPW N12LL W=570.00n L=60.00n
MM47 net97 S0 net61 VPW N12LL W=430.00n L=60.00n
MM69 net105 S1 net73 VPW N12LL W=570.00n L=60.00n
MM70 net101 S0 net67 VPW N12LL W=430.00n L=60.00n
MM72 net101 I3 VSS VPW N12LL W=430.00n L=60.00n
MM49 net95 I0 VSS VPW N12LL W=430.00n L=60.00n
MM73 net99 net107 net67 VPW N12LL W=430.00n L=60.00n
MM63 ZN net73 VSS VPW N12LL W=860.00n L=60.00n
MM65 net111 S1 VSS VPW N12LL W=430.00n L=60.00n
MM31 net97 I1 VSS VPW N12LL W=430.00n L=60.00n
MM53 net107 S0 VSS VPW N12LL W=650.00n L=60.00n
MM71 net99 I2 VSS VPW N12LL W=430.00n L=60.00n
MM36 net95 net107 net61 VPW N12LL W=430.00n L=60.00n
MM81 net105 net67 VDD VNW P12LL W=960.00n L=60.00n
MM50 net95 I0 VDD VNW P12LL W=640.00n L=60.00n
MM62 net103 S1 net73 VNW P12LL W=870.00n L=60.00n
MM48 net97 net107 net61 VNW P12LL W=635.00n L=60.00n
MM74 net99 I2 VDD VNW P12LL W=640.00n L=60.00n
MM76 net105 net111 net73 VNW P12LL W=870.00n L=60.00n
MM77 net101 net107 net67 VNW P12LL W=635.00n L=60.00n
MM78 net101 I3 VDD VNW P12LL W=640.00n L=60.00n
MM79 net99 S0 net67 VNW P12LL W=635.00n L=60.00n
MM64 ZN net73 VDD VNW P12LL W=1.3u L=60.00n
MM66 net111 S1 VDD VNW P12LL W=650.0n L=60.00n
MM32 net97 I1 VDD VNW P12LL W=635.00n L=60.00n
MM80 net103 net61 VDD VNW P12LL W=870.00n L=60.00n
MM54 net107 S0 VDD VNW P12LL W=980.00n L=60.00n
MM39 net95 S0 net61 VNW P12LL W=640.00n L=60.00n
.ENDS MUX4NHSV4
****Sub-Circuit for NAND2HSV0, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT NAND2HSV0 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS NAND2HSV0
****Sub-Circuit for NAND2HSV0P5, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND2HSV0P5 A1 A2 ZN VDD VSS
MM1 net4 A2 VSS VPW N12LL W=350.00n L=60.00n
MM2 ZN A1 net4 VPW N12LL W=350.00n L=60.00n
MM3 ZN A2 VDD VNW P12LL W=310.00n L=60.00n
MM0 ZN A1 VDD VNW P12LL W=310.00n L=60.00n
.ENDS NAND2HSV0P5
****Sub-Circuit for NAND2HSV1, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT NAND2HSV1 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=290.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=290.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=440.00n L=60.00n
.ENDS NAND2HSV1
****Sub-Circuit for NAND2HSV12, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND2HSV12 A1 A2 ZN VDD VSS
MM1 net4 A2 VSS VPW N12LL W=3.24u L=60.00n
MM2 ZN A1 net4 VPW N12LL W=3.24u L=60.00n
MM3 ZN A2 VDD VNW P12LL W=2.88u L=60.00n
MM0 ZN A1 VDD VNW P12LL W=2.88u L=60.00n
.ENDS NAND2HSV12
****Sub-Circuit for NAND2HSV16, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND2HSV16 A1 A2 ZN VDD VSS
MM1 net4 A2 VSS VPW N12LL W=4.32u L=60.00n
MM2 ZN A1 net4 VPW N12LL W=4.32u L=60.00n
MM3 ZN A2 VDD VNW P12LL W=3.84u L=60.00n
MM0 ZN A1 VDD VNW P12LL W=3.84u L=60.00n
.ENDS NAND2HSV16
****Sub-Circuit for NAND2HSV2, Wed Dec  8 11:21:16 CST 2010****
.SUBCKT NAND2HSV2 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=430.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=430.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=650.00n L=60.00n
.ENDS NAND2HSV2
****Sub-Circuit for NAND2HSV24, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND2HSV24 A1 A2 ZN VDD VSS
MM1 net4 A2 VSS VPW N12LL W=6.48u L=60.00n
MM2 ZN A1 net4 VPW N12LL W=6.48u L=60.00n
MM3 ZN A2 VDD VNW P12LL W=5.76u L=60.00n
MM0 ZN A1 VDD VNW P12LL W=5.76u L=60.00n
.ENDS NAND2HSV24
****Sub-Circuit for NAND2HSV3, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND2HSV3 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=650.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=650.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=980.0n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=980.0n L=60.00n
.ENDS NAND2HSV3
****Sub-Circuit for NAND2HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND2HSV4 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=860.00n L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=860.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=1.30u L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=1.30u L=60.00n
.ENDS NAND2HSV4
****Sub-Circuit for NAND2HSV8, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND2HSV8 A1 A2 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=1.66u L=60.00n
MMN1 net18 A2 VSS VPW N12LL W=1.66u L=60.00n
MM0 ZN A2 VDD VNW P12LL W=2.54u L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=2.54u L=60.00n
.ENDS NAND2HSV8
****Sub-Circuit for NAND3HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND3HSV0 A1 A2 A3 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=200.00n L=60.00n
MM3 net022 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=200.00n L=60.00n
MM2 ZN A3 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS NAND3HSV0
****Sub-Circuit for NAND3HSV0P5, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND3HSV0P5 A1 A2 A3 ZN VDD VSS
MM3 ZN A2 VDD VNW P12LL W=240.00n L=60.00n
MM0 ZN A1 VDD VNW P12LL W=240.00n L=60.00n
MM4 ZN A3 VDD VNW P12LL W=240.00n L=60.00n
MM1 net17 A3 VSS VPW N12LL W=350.00n L=60.00n
MM2 net21 A2 net17 VPW N12LL W=350.00n L=60.00n
MM5 ZN A1 net21 VPW N12LL W=350.00n L=60.00n
.ENDS NAND3HSV0P5
****Sub-Circuit for NAND3HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND3HSV1 A1 A2 A3 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=290.00n L=60.00n
MM3 net022 A3 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=290.00n L=60.00n
MM2 ZN A3 VDD VNW P12LL W=440.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=440.00n L=60.00n
.ENDS NAND3HSV1
****Sub-Circuit for NAND3HSV12, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND3HSV12 A1 A2 A3 ZN VDD VSS
MM3 ZN A2 VDD VNW P12LL W=2.24u L=60.00n
MM0 ZN A1 VDD VNW P12LL W=2.24u L=60.00n
MM4 ZN A3 VDD VNW P12LL W=2.24u L=60.00n
MM1 net17 A3 VSS VPW N12LL W=3.24u L=60.00n
MM2 net21 A2 net17 VPW N12LL W=3.24u L=60.00n
MM5 ZN A1 net21 VPW N12LL W=3.24u L=60.00n
.ENDS NAND3HSV12
****Sub-Circuit for NAND3HSV16, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND3HSV16 A1 A2 A3 ZN VDD VSS
MM3 ZN A2 VDD VNW P12LL W=2.98u L=60.00n
MM0 ZN A1 VDD VNW P12LL W=2.98u L=60.00n
MM4 ZN A3 VDD VNW P12LL W=2.98u L=60.00n
MM1 net17 A3 VSS VPW N12LL W=4.32u L=60.00n
MM2 net21 A2 net17 VPW N12LL W=4.32u L=60.00n
MM5 ZN A1 net21 VPW N12LL W=4.32u L=60.00n
.ENDS NAND3HSV16
****Sub-Circuit for NAND3HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND3HSV2 A1 A2 A3 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=430.00n L=60.00n
MM3 net022 A3 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=430.00n L=60.00n
MM2 ZN A3 VDD VNW P12LL W=650.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=650.00n L=60.00n
.ENDS NAND3HSV2
****Sub-Circuit for NAND3HSV24, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND3HSV24 A1 A2 A3 ZN VDD VSS
MM3 ZN A2 VDD VNW P12LL W=4.47u L=60.00n
MM0 ZN A1 VDD VNW P12LL W=4.47u L=60.00n
MM4 ZN A3 VDD VNW P12LL W=4.47u L=60.00n
MM1 net17 A3 VSS VPW N12LL W=6.48u L=60.00n
MM2 net21 A2 net17 VPW N12LL W=6.48u L=60.00n
MM5 ZN A1 net21 VPW N12LL W=6.48u L=60.00n
.ENDS NAND3HSV24
****Sub-Circuit for NAND3HSV3, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND3HSV3 A1 A2 A3 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=650.00n L=60.00n
MM3 net022 A3 VSS VPW N12LL W=650.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=650.00n L=60.00n
MM2 ZN A3 VDD VNW P12LL W=980.0n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=980.0n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=980.0n L=60.00n
.ENDS NAND3HSV3
****Sub-Circuit for NAND3HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND3HSV4 A1 A2 A3 ZN VDD VSS
MM1 ZN A1 net18 VPW N12LL W=830.00n L=60.00n
MM3 net022 A3 VSS VPW N12LL W=830.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=830.00n L=60.00n
MM2 ZN A3 VDD VNW P12LL W=1.27u L=60.00n
MM0 ZN A2 VDD VNW P12LL W=1.27u L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=1.27u L=60.00n
.ENDS NAND3HSV4
****Sub-Circuit for NAND3HSV8, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND3HSV8 A1 A2 A3 ZN VDD VSS
MM6 ZN net029 VSS VPW N12LL W=1.72u L=60.00n
MM1 net053 A1 net18 VPW N12LL W=270.00n L=60.00n
MM4 net029 net053 VSS VPW N12LL W=680.00n L=60.00n
MM3 net022 A3 VSS VPW N12LL W=270.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=270.00n L=60.00n
MM5 net029 net053 VDD VNW P12LL W=1.0u L=60.00n
MM7 ZN net029 VDD VNW P12LL W=2.60u L=60.00n
MM2 net053 A3 VDD VNW P12LL W=400.00n L=60.00n
MM0 net053 A2 VDD VNW P12LL W=400.00n L=60.00n
MMP1 net053 A1 VDD VNW P12LL W=400.00n L=60.00n
.ENDS NAND3HSV8
****Sub-Circuit for NAND4HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND4HSV0 A1 A2 A3 A4 ZN VDD VSS
MM4 net026 A4 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 net18 VPW N12LL W=200.00n L=60.00n
MM3 net022 A3 net026 VPW N12LL W=200.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=200.00n L=60.00n
MM5 ZN A4 VDD VNW P12LL W=300.00n L=60.00n
MM2 ZN A3 VDD VNW P12LL W=300.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=300.00n L=60.00n
.ENDS NAND4HSV0
****Sub-Circuit for NAND4HSV0P5, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND4HSV0P5 A1 A2 A3 A4 ZN VDD VSS
MM3 ZN A3 VDD VNW P12LL W=190.00n L=60.00n
MM4 ZN A4 VDD VNW P12LL W=190.00n L=60.00n
MM7 ZN A1 VDD VNW P12LL W=190.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=190.00n L=60.00n
MM1 net22 A4 VSS VPW N12LL W=350.00n L=60.00n
MM2 net26 A3 net22 VPW N12LL W=350.00n L=60.00n
MM5 net30 A2 net26 VPW N12LL W=350.00n L=60.00n
MM6 ZN A1 net30 VPW N12LL W=350.00n L=60.00n
.ENDS NAND4HSV0P5
****Sub-Circuit for NAND4HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND4HSV1 A1 A2 A3 A4 ZN VDD VSS
MM4 net026 A4 VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 net18 VPW N12LL W=290.00n L=60.00n
MM3 net022 A3 net026 VPW N12LL W=290.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=290.00n L=60.00n
MM5 ZN A4 VDD VNW P12LL W=440.00n L=60.00n
MM2 ZN A3 VDD VNW P12LL W=440.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=440.00n L=60.00n
.ENDS NAND4HSV1
****Sub-Circuit for NAND4HSV12, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND4HSV12 A1 A2 A3 A4 ZN VDD VSS
MM3 ZN A3 VDD VNW P12LL W=1.75u L=60.00n
MM4 ZN A4 VDD VNW P12LL W=1.75u L=60.00n
MM7 ZN A1 VDD VNW P12LL W=1.75u L=60.00n
MM0 ZN A2 VDD VNW P12LL W=1.75u L=60.00n
MM1 net22 A4 VSS VPW N12LL W=3.24u L=60.00n
MM2 net26 A3 net22 VPW N12LL W=3.24u L=60.00n
MM5 net30 A2 net26 VPW N12LL W=3.24u L=60.00n
MM6 ZN A1 net30 VPW N12LL W=3.24u L=60.00n
.ENDS NAND4HSV12
****Sub-Circuit for NAND4HSV16, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND4HSV16 A1 A2 A3 A4 ZN VDD VSS
MM3 ZN A3 VDD VNW P12LL W=2.33u L=60.00n
MM4 ZN A4 VDD VNW P12LL W=2.33u L=60.00n
MM7 ZN A1 VDD VNW P12LL W=2.33u L=60.00n
MM0 ZN A2 VDD VNW P12LL W=2.33u L=60.00n
MM1 net22 A4 VSS VPW N12LL W=4.32u L=60.00n
MM2 net26 A3 net22 VPW N12LL W=4.32u L=60.00n
MM5 net30 A2 net26 VPW N12LL W=4.32u L=60.00n
MM6 ZN A1 net30 VPW N12LL W=4.32u L=60.00n
.ENDS NAND4HSV16
****Sub-Circuit for NAND4HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND4HSV2 A1 A2 A3 A4 ZN VDD VSS
MM4 net026 A4 VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 net18 VPW N12LL W=430.00n L=60.00n
MM3 net022 A3 net026 VPW N12LL W=430.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=430.00n L=60.00n
MM5 ZN A4 VDD VNW P12LL W=650.00n L=60.00n
MM2 ZN A3 VDD VNW P12LL W=650.00n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=650.00n L=60.00n
.ENDS NAND4HSV2
****Sub-Circuit for NAND4HSV24, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NAND4HSV24 A1 A2 A3 A4 ZN VDD VSS
MM3 ZN A3 VDD VNW P12LL W=3.5u L=60.00n
MM4 ZN A4 VDD VNW P12LL W=3.5u L=60.00n
MM7 ZN A1 VDD VNW P12LL W=3.5u L=60.00n
MM0 ZN A2 VDD VNW P12LL W=3.5u L=60.00n
MM1 net22 A4 VSS VPW N12LL W=6.48u L=60.00n
MM2 net26 A3 net22 VPW N12LL W=6.48u L=60.00n
MM5 net30 A2 net26 VPW N12LL W=6.48u L=60.00n
MM6 ZN A1 net30 VPW N12LL W=6.48u L=60.00n
.ENDS NAND4HSV24
****Sub-Circuit for NAND4HSV3, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND4HSV3 A1 A2 A3 A4 ZN VDD VSS
MM4 net026 A4 VSS VPW N12LL W=650.00n L=60.00n
MM1 ZN A1 net18 VPW N12LL W=650.00n L=60.00n
MM3 net022 A3 net026 VPW N12LL W=650.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=650.00n L=60.00n
MM5 ZN A4 VDD VNW P12LL W=980.0n L=60.00n
MM2 ZN A3 VDD VNW P12LL W=980.0n L=60.00n
MM0 ZN A2 VDD VNW P12LL W=980.0n L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=980.0n L=60.00n
.ENDS NAND4HSV3
****Sub-Circuit for NAND4HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND4HSV4 A1 A2 A3 A4 ZN VDD VSS
MM4 net026 A4 VSS VPW N12LL W=860.00n L=60.00n
MM1 ZN A1 net18 VPW N12LL W=860.00n L=60.00n
MM3 net022 A3 net026 VPW N12LL W=860.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=860.00n L=60.00n
MM5 ZN A4 VDD VNW P12LL W=1.29u L=60.00n
MM2 ZN A3 VDD VNW P12LL W=1.29u L=60.00n
MM0 ZN A2 VDD VNW P12LL W=1.29u L=60.00n
MMP1 ZN A1 VDD VNW P12LL W=1.29u L=60.00n
.ENDS NAND4HSV4
****Sub-Circuit for NAND4HSV8, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NAND4HSV8 A1 A2 A3 A4 ZN VDD VSS
MM6 net068 net096 VSS VPW N12LL W=680.00n L=60.00n
MM8 ZN net068 VSS VPW N12LL W=1.72u L=60.00n
MM4 net026 A4 VSS VPW N12LL W=270.00n L=60.00n
MM1 net096 A1 net18 VPW N12LL W=270.00n L=60.00n
MM3 net022 A3 net026 VPW N12LL W=270.00n L=60.00n
MMN1 net18 A2 net022 VPW N12LL W=270.00n L=60.00n
MM7 net068 net096 VDD VNW P12LL W=1.0u L=60.00n
MM9 ZN net068 VDD VNW P12LL W=2.60u L=60.00n
MM5 net096 A4 VDD VNW P12LL W=400n L=60.00n
MM2 net096 A3 VDD VNW P12LL W=400n L=60.00n
MM0 net096 A2 VDD VNW P12LL W=400n L=60.00n
MMP1 net096 A1 VDD VNW P12LL W=400n L=60.00n
.ENDS NAND4HSV8
****Sub-Circuit for NDHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDHSV1 CKN D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=290.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=290.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM43 QN s VDD VNW P12LL W=440.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDHSV1
****Sub-Circuit for NDHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDHSV2 CKN D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n
MM39 net43 c net_099 VPW N12LL W=230.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=230.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n
MM38 net43 cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=480.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDHSV2
****Sub-Circuit for NDHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDHSV4 CKN D Q QN VDD VSS
MM42 QN s VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 net43 c net_099 VPW N12LL W=400.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=400.00n L=60.00n
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM17 s net43 VSS VPW N12LL W=400.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 m pm VSS VPW N12LL W=200.00n L=60.00n
MM43 QN s VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 net43 cn net_0158 VNW P12LL W=450.00n L=60.00n m=2
MM41 net_0158 m VDD VNW P12LL W=450.00n L=60.00n m=2
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM18 s net43 VDD VNW P12LL W=600.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 m pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDHSV4
****Sub-Circuit for NDRNHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRNHSV1 CKN D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=200.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=200.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=440.00n L=60.00n
.ENDS NDRNHSV1
****Sub-Circuit for NDRNHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRNHSV2 CKN D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=200.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=300.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=200.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS NDRNHSV2
****Sub-Circuit for NDRNHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRNHSV4 CKN D Q QN RDN VDD VSS
MM45 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM3 net_0154 c net43 VPW N12LL W=360.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=200.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=190.00n L=60.00n
MM39 s net43 net_099 VPW N12LL W=280.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=280.00n L=60.00n m=2
MM30 cn c VSS VPW N12LL W=430.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=190.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=190.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D net_0104 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm VSS VPW N12LL W=260.00n L=60.00n
MM46 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM43 pm RDN VDD VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=560n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=650.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=650.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=530.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=300.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=610.00n L=60.00n
.ENDS NDRNHSV4
****Sub-Circuit for NDRSNHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRSNHSV1 CKN D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=200.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=200.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=380.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=440.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=350.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=440.00n L=60.00n
.ENDS NDRSNHSV1
****Sub-Circuit for NDRSNHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRSNHSV2 CKN D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=250.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=260.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=240.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=250.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=250.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=240.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=320.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=460.00n L=60.00n m=1
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=650.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=580.00n L=60.00n
.ENDS NDRSNHSV2
****Sub-Circuit for NDRSNHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDRSNHSV4 CKN D Q QN RDN SDN VDD VSS
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R net_0132 VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=260.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=240.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM40 net43 R net_0132 VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=420.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=430.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=240.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 s net43 VDD VNW P12LL W=470.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0243 R VDD VNW P12LL W=460n L=60.00n
MM29 cn c VDD VNW P12LL W=640.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=650.00n L=60.00n
MM26 net_0243 s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=430.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=400.00n L=60.00n
MM1 net_0154 pm net_0243 VNW P12LL W=620.00n L=60.00n
.ENDS NDRSNHSV4
****Sub-Circuit for NDSNHSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDSNHSV1 CKN D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=200.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=290.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=270.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=290.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=300.00n L=60.00n
.ENDS NDSNHSV1
****Sub-Circuit for NDSNHSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDSNHSV2 CKN D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=260.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=390.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM30 cn c VSS VPW N12LL W=200.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=390.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=300.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=395.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=395.00n L=60.00n
.ENDS NDSNHSV2
****Sub-Circuit for NDSNHSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NDSNHSV4 CKN D Q QN SDN VDD VSS
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=390.00n L=60.00n
MM30 cn c VSS VPW N12LL W=400.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=400.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 pm cn net69 VPW N12LL W=200.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=200.00n L=60.00n
MM0 net_0154 pm net_0132 VPW N12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM38 s net43 VDD VNW P12LL W=580.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=600.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=600.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 pm c net128 VNW P12LL W=440.00n L=60.00n
MM8 net128 D VDD VNW P12LL W=440.00n L=60.00n
MM1 net_0154 pm VDD VNW P12LL W=620.00n L=60.00n
.ENDS NDSNHSV4
****Sub-Circuit for NOR2HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR2HSV0 A1 A2 ZN VDD VSS
MM0 ZN A2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 net34 VNW P12LL W=300.00n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=300.00n L=60.00n
.ENDS NOR2HSV0
****Sub-Circuit for NOR2HSV0P5, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NOR2HSV0P5 A1 A2 ZN VDD VSS
MM3 net11 A2 VDD VNW P12LL W=320.00n L=60.00n
MM0 ZN A1 net11 VNW P12LL W=320.00n L=60.00n
MM1 ZN A1 VSS VPW N12LL W=240.00n L=60.00n
MM2 ZN A2 VSS VPW N12LL W=240.00n L=60.00n
.ENDS NOR2HSV0P5
****Sub-Circuit for NOR2HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR2HSV1 A1 A2 ZN VDD VSS
MM0 ZN A2 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 net34 VNW P12LL W=440.00n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=440.00n L=60.00n
.ENDS NOR2HSV1
****Sub-Circuit for NOR2HSV12, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NOR2HSV12 A1 A2 ZN VDD VSS
MM3 net11 A2 VDD VNW P12LL W=3.9u L=60.00n
MM0 ZN A1 net11 VNW P12LL W=3.9u L=60.00n
MM1 ZN A1 VSS VPW N12LL W=2.1u L=60.00n
MM2 ZN A2 VSS VPW N12LL W=2.1u L=60.00n
.ENDS NOR2HSV12
****Sub-Circuit for NOR2HSV16, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NOR2HSV16 A1 A2 ZN VDD VSS
MM3 net11 A2 VDD VNW P12LL W=5.2u L=60.00n
MM0 ZN A1 net11 VNW P12LL W=5.2u L=60.00n
MM1 ZN A1 VSS VPW N12LL W=2.8u L=60.00n
MM2 ZN A2 VSS VPW N12LL W=2.8u L=60.00n
.ENDS NOR2HSV16
****Sub-Circuit for NOR2HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR2HSV2 A1 A2 ZN VDD VSS
MM0 ZN A2 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 net34 VNW P12LL W=650.00n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=650.00n L=60.00n
.ENDS NOR2HSV2
****Sub-Circuit for NOR2HSV24, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NOR2HSV24 A1 A2 ZN VDD VSS
MM3 net11 A2 VDD VNW P12LL W=7.8u L=60.00n
MM0 ZN A1 net11 VNW P12LL W=7.8u L=60.00n
MM1 ZN A1 VSS VPW N12LL W=4.2u L=60.00n
MM2 ZN A2 VSS VPW N12LL W=4.2u L=60.00n
.ENDS NOR2HSV24
****Sub-Circuit for NOR2HSV3, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR2HSV3 A1 A2 ZN VDD VSS
MM0 ZN A2 VSS VPW N12LL W=650.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=650.00n L=60.00n
MM1 ZN A1 net34 VNW P12LL W=980.00n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=980.00n L=60.00n
.ENDS NOR2HSV3
****Sub-Circuit for NOR2HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR2HSV4 A1 A2 ZN VDD VSS
MM0 ZN A2 VSS VPW N12LL W=860.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=860.00n L=60.00n
MM1 ZN A1 net34 VNW P12LL W=1.3u L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=1.3u L=60.00n
.ENDS NOR2HSV4
****Sub-Circuit for NOR2HSV8, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR2HSV8 A1 A2 ZN VDD VSS
MM0 ZN A2 VSS VPW N12LL W=1.72u L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=1.72u L=60.00n
MM1 ZN A1 net34 VNW P12LL W=2.6u L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=2.6u L=60.00n
.ENDS NOR2HSV8
****Sub-Circuit for NOR3HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR3HSV0 A1 A2 A3 ZN VDD VSS
MM3 ZN A3 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=200.00n L=60.00n
MM2 net47 A3 VDD VNW P12LL W=300.00n L=60.00n
MM1 ZN A1 net43 VNW P12LL W=300.00n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=300.00n L=60.00n
.ENDS NOR3HSV0
****Sub-Circuit for NOR3HSV0P5, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NOR3HSV0P5 A1 A2 A3 ZN VDD VSS
MM4 ZN A3 VSS VPW N12LL W=190.00n L=60.00n
MM2 ZN A2 VSS VPW N12LL W=190.00n L=60.00n
MM1 ZN A1 VSS VPW N12LL W=190.00n L=60.00n
MM5 ZN A1 net20 VNW P12LL W=320.00n L=60.00n
MM0 net20 A2 net24 VNW P12LL W=320.00n L=60.00n
MM3 net24 A3 VDD VNW P12LL W=320.00n L=60.00n
.ENDS NOR3HSV0P5
****Sub-Circuit for NOR3HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR3HSV1 A1 A2 A3 ZN VDD VSS
MM3 ZN A3 VSS VPW N12LL W=290.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=290.00n L=60.00n
MM2 net47 A3 VDD VNW P12LL W=440.00n L=60.00n
MM1 ZN A1 net43 VNW P12LL W=440.00n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=440.00n L=60.00n
.ENDS NOR3HSV1
****Sub-Circuit for NOR3HSV12, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NOR3HSV12 A1 A2 A3 ZN VDD VSS
MM4 ZN A3 VSS VPW N12LL W=1.62u L=60.00n
MM2 ZN A2 VSS VPW N12LL W=1.62u L=60.00n
MM1 ZN A1 VSS VPW N12LL W=1.62u L=60.00n
MM5 ZN A1 net20 VNW P12LL W=3.9u L=60.00n
MM0 net20 A2 net24 VNW P12LL W=3.9u L=60.00n
MM3 net24 A3 VDD VNW P12LL W=3.9u L=60.00n
.ENDS NOR3HSV12
****Sub-Circuit for NOR3HSV16, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NOR3HSV16 A1 A2 A3 ZN VDD VSS
MM4 ZN A3 VSS VPW N12LL W=2.16u L=60.00n
MM2 ZN A2 VSS VPW N12LL W=2.16u L=60.00n
MM1 ZN A1 VSS VPW N12LL W=2.16u L=60.00n
MM5 ZN A1 net20 VNW P12LL W=5.2u L=60.00n
MM0 net20 A2 net24 VNW P12LL W=5.2u L=60.00n
MM3 net24 A3 VDD VNW P12LL W=5.2u L=60.00n
.ENDS NOR3HSV16
****Sub-Circuit for NOR3HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR3HSV2 A1 A2 A3 ZN VDD VSS
MM3 ZN A3 VSS VPW N12LL W=430.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=430.00n L=60.00n
MM2 net47 A3 VDD VNW P12LL W=650.00n L=60.00n
MM1 ZN A1 net43 VNW P12LL W=650.00n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=650.00n L=60.00n
.ENDS NOR3HSV2
****Sub-Circuit for NOR3HSV24, Wed Dec  8 16:10:28 CST 2010****
.SUBCKT NOR3HSV24 A1 A2 A3 ZN VDD VSS
MM4 ZN A3 VSS VPW N12LL W=3.24u L=60.00n
MM2 ZN A2 VSS VPW N12LL W=3.24u L=60.00n
MM1 ZN A1 VSS VPW N12LL W=3.24u L=60.00n
MM5 ZN A1 net20 VNW P12LL W=7.8u L=60.00n
MM0 net20 A2 net24 VNW P12LL W=7.8u L=60.00n
MM3 net24 A3 VDD VNW P12LL W=7.8u L=60.00n
.ENDS NOR3HSV24
****Sub-Circuit for NOR3HSV3, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR3HSV3 A1 A2 A3 ZN VDD VSS
MM3 ZN A3 VSS VPW N12LL W=650.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=650.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=650.00n L=60.00n
MM2 net47 A3 VDD VNW P12LL W=980.00n L=60.00n
MM1 ZN A1 net43 VNW P12LL W=980.00n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=980.00n L=60.00n
.ENDS NOR3HSV3
****Sub-Circuit for NOR3HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR3HSV4 A1 A2 A3 ZN VDD VSS
MM3 ZN A3 VSS VPW N12LL W=860.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=860.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=860.00n L=60.00n
MM2 net47 A3 VDD VNW P12LL W=1.3u L=60.00n
MM1 ZN A1 net43 VNW P12LL W=1.3u L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=1.3u L=60.00n
.ENDS NOR3HSV4
****Sub-Circuit for NOR3HSV8, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR3HSV8 A1 A2 A3 ZN VDD VSS
MM5 net027 net039 VSS VPW N12LL W=680.00n L=60.00n
MM3 net039 A3 VSS VPW N12LL W=270.0n L=60.00n
MM0 net039 A2 VSS VPW N12LL W=270.0n L=60.00n
MM6 ZN net027 VSS VPW N12LL W=1.72u L=60.00n
MMN1 net039 A1 VSS VPW N12LL W=270.0n L=60.00n
MM7 ZN net027 VDD VNW P12LL W=2.6u L=60.00n
MM4 net027 net039 VDD VNW P12LL W=1.02u L=60.00n
MM2 net47 A3 VDD VNW P12LL W=410.00n L=60.00n
MM1 net039 A1 net43 VNW P12LL W=410.00n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=410.00n L=60.00n
.ENDS NOR3HSV8
****Sub-Circuit for NOR4HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR4HSV0 A1 A2 A3 A4 ZN VDD VSS
MM4 ZN A4 VSS VPW N12LL W=200.00n L=60.00n
MM3 ZN A3 VSS VPW N12LL W=200.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=200.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=200.00n L=60.00n
MM5 net047 A4 VDD VNW P12LL W=300.0n L=60.00n
MM2 net47 A3 net047 VNW P12LL W=300.0n L=60.00n
MM1 ZN A1 net43 VNW P12LL W=300.0n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=300.0n L=60.00n
.ENDS NOR4HSV0
****Sub-Circuit for NOR4HSV0P5, Thu May 19 13:57:40 CST 2011****
.SUBCKT NOR4HSV0P5 A1 A2 A3 A4 ZN VDD VSS
MM3 net13 A3 net9 VNW P12LL W=320.00n L=60.00n
MM0 net17 A2 net13 VNW P12LL W=320.00n L=60.00n
MM5 ZN A1 net17 VNW P12LL W=320.00n L=60.00n
MM6 net9 A4 VDD VNW P12LL W=320.00n L=60.00n
MM1 ZN A1 VSS VPW N12LL W=180.00n L=60.00n
MM2 ZN A2 VSS VPW N12LL W=180.00n L=60.00n
MM4 ZN A3 VSS VPW N12LL W=180.00n L=60.00n
MM7 ZN A4 VSS VPW N12LL W=180.00n L=60.00n
.ENDS NOR4HSV0P5
****Sub-Circuit for NOR4HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR4HSV1 A1 A2 A3 A4 ZN VDD VSS
MM4 ZN A4 VSS VPW N12LL W=290.00n L=60.00n
MM3 ZN A3 VSS VPW N12LL W=290.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=290.00n L=60.00n
MM5 net047 A4 VDD VNW P12LL W=440.0n L=60.00n
MM2 net47 A3 net047 VNW P12LL W=440.0n L=60.00n
MM1 ZN A1 net43 VNW P12LL W=440.0n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=440.0n L=60.00n
.ENDS NOR4HSV1
****Sub-Circuit for NOR4HSV12, Wed Dec  8 16:10:29 CST 2010****
.SUBCKT NOR4HSV12 A1 A2 A3 A4 ZN VDD VSS
MM3 net13 A3 net9 VNW P12LL W=3.9u L=60.00n
MM0 net17 A2 net13 VNW P12LL W=3.9u L=60.00n
MM5 ZN A1 net17 VNW P12LL W=3.9u L=60.00n
MM6 net9 A4 VDD VNW P12LL W=3.9u L=60.00n
MM1 ZN A1 VSS VPW N12LL W=1.38u L=60.00n
MM2 ZN A2 VSS VPW N12LL W=1.38u L=60.00n
MM4 ZN A3 VSS VPW N12LL W=1.38u L=60.00n
MM7 ZN A4 VSS VPW N12LL W=1.38u L=60.00n
.ENDS NOR4HSV12
****Sub-Circuit for NOR4HSV16, Wed Dec  8 16:10:29 CST 2010****
.SUBCKT NOR4HSV16 A1 A2 A3 A4 ZN VDD VSS
MM3 net13 A3 net9 VNW P12LL W=5.2u L=60.00n
MM0 net17 A2 net13 VNW P12LL W=5.2u L=60.00n
MM5 ZN A1 net17 VNW P12LL W=5.2u L=60.00n
MM6 net9 A4 VDD VNW P12LL W=5.2u L=60.00n
MM1 ZN A1 VSS VPW N12LL W=1.84u L=60.00n
MM2 ZN A2 VSS VPW N12LL W=1.84u L=60.00n
MM4 ZN A3 VSS VPW N12LL W=1.84u L=60.00n
MM7 ZN A4 VSS VPW N12LL W=1.84u L=60.00n
.ENDS NOR4HSV16
****Sub-Circuit for NOR4HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR4HSV2 A1 A2 A3 A4 ZN VDD VSS
MM4 ZN A4 VSS VPW N12LL W=430.00n L=60.00n
MM3 ZN A3 VSS VPW N12LL W=430.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=430.00n L=60.00n
MM5 net047 A4 VDD VNW P12LL W=650.0n L=60.00n
MM2 net47 A3 net047 VNW P12LL W=650.0n L=60.00n
MM1 ZN A1 net43 VNW P12LL W=650.0n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=650.0n L=60.00n
.ENDS NOR4HSV2
****Sub-Circuit for NOR4HSV24, Wed Dec  8 16:10:29 CST 2010****
.SUBCKT NOR4HSV24 A1 A2 A3 A4 ZN VDD VSS
MM3 net13 A3 net9 VNW P12LL W=7.8u L=60.00n
MM0 net17 A2 net13 VNW P12LL W=7.8u L=60.00n
MM5 ZN A1 net17 VNW P12LL W=7.8u L=60.00n
MM6 net9 A4 VDD VNW P12LL W=7.8u L=60.00n
MM1 ZN A1 VSS VPW N12LL W=2.76u L=60.00n
MM2 ZN A2 VSS VPW N12LL W=2.76u L=60.00n
MM4 ZN A3 VSS VPW N12LL W=2.76u L=60.00n
MM7 ZN A4 VSS VPW N12LL W=2.76u L=60.00n
.ENDS NOR4HSV24
****Sub-Circuit for NOR4HSV3, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR4HSV3 A1 A2 A3 A4 ZN VDD VSS
MM4 ZN A4 VSS VPW N12LL W=650.00n L=60.00n
MM3 ZN A3 VSS VPW N12LL W=650.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=650.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=650.00n L=60.00n
MM5 net047 A4 VDD VNW P12LL W=980.0n L=60.00n
MM2 net47 A3 net047 VNW P12LL W=980.0n L=60.00n
MM1 ZN A1 net43 VNW P12LL W=980.0n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=980.0n L=60.00n
.ENDS NOR4HSV3
****Sub-Circuit for NOR4HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR4HSV4 A1 A2 A3 A4 ZN VDD VSS
MM4 ZN A4 VSS VPW N12LL W=860.00n L=60.00n
MM3 ZN A3 VSS VPW N12LL W=860.00n L=60.00n
MM0 ZN A2 VSS VPW N12LL W=860.00n L=60.00n
MMN1 ZN A1 VSS VPW N12LL W=860.00n L=60.00n
MM5 net047 A4 VDD VNW P12LL W=1.3u L=60.00n
MM2 net47 A3 net047 VNW P12LL W=1.3u L=60.00n
MM1 ZN A1 net43 VNW P12LL W=1.3u L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=1.3u L=60.00n
.ENDS NOR4HSV4
****Sub-Circuit for NOR4HSV8, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT NOR4HSV8 A1 A2 A3 A4 ZN VDD VSS
MM7 net033 net049 VSS VPW N12LL W=680.00n L=60.00n
MM8 ZN net033 VSS VPW N12LL W=1.72u L=60.00n
MM4 net049 A4 VSS VPW N12LL W=270.00n L=60.00n
MM3 net049 A3 VSS VPW N12LL W=270.00n L=60.00n
MM0 net049 A2 VSS VPW N12LL W=270.00n L=60.00n
MMN1 net049 A1 VSS VPW N12LL W=270.00n L=60.00n
MM6 net033 net049 VDD VNW P12LL W=1.02u L=60.00n
MM9 ZN net033 VDD VNW P12LL W=2.6u L=60.00n
MM5 net047 A4 VDD VNW P12LL W=410.00n L=60.00n
MM2 net47 A3 net047 VNW P12LL W=410.00n L=60.00n
MM1 net049 A1 net43 VNW P12LL W=410.00n L=60.00n
MMP1 net43 A2 net47 VNW P12LL W=410.00n L=60.00n
.ENDS NOR4HSV8
****Sub-Circuit for OA211HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA211HSV0 A1 A2 B C Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=200.00n L=60.00n
MM2 net18 B net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 C VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=300.00n L=60.00n
MM4 net064 B VDD VNW P12LL W=300.00n L=60.00n
MM5 net064 C VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA211HSV0
****Sub-Circuit for OA211HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA211HSV1 A1 A2 B C Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=290.00n L=60.00n
MM2 net18 B net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 C VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=440.00n L=60.00n
MM4 net064 B VDD VNW P12LL W=300.00n L=60.00n
MM5 net064 C VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA211HSV1
****Sub-Circuit for OA211HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA211HSV2 A1 A2 B C Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=430.00n L=60.00n
MM2 net18 B net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 C VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=440.00n L=60.00n
MM4 net064 B VDD VNW P12LL W=300.00n L=60.00n
MM5 net064 C VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA211HSV2
****Sub-Circuit for OA211HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA211HSV4 A1 A2 B C Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=860.00n L=60.00n
MM2 net18 B net030 VPW N12LL W=350.000n L=60.00n
MM3 net030 C VSS VPW N12LL W=350.000n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=350.000n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=350.000n L=60.00n
MM6 Z net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net064 B VDD VNW P12LL W=520.00n L=60.00n
MM5 net064 C VDD VNW P12LL W=520.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=520.00n L=60.00n
.ENDS OA211HSV4
****Sub-Circuit for OA21HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA21HSV0 A1 A2 B Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=200.00n L=60.00n
MM2 net064 B net029 VPW N12LL W=200.00n L=60.00n
MM1 net029 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net029 A2 VSS VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=300.00n L=60.00n
MM4 net064 B VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA21HSV0
****Sub-Circuit for OA21HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA21HSV1 A1 A2 B Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=290.00n L=60.00n
MM2 net064 B net029 VPW N12LL W=200.00n L=60.00n
MM1 net029 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net029 A2 VSS VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=440.00n L=60.00n
MM4 net064 B VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA21HSV1
****Sub-Circuit for OA21HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA21HSV2 A1 A2 B Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=430.00n L=60.00n
MM2 net064 B net029 VPW N12LL W=200.00n L=60.00n
MM1 net029 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net029 A2 VSS VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=650.00n L=60.00n
MM4 net064 B VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA21HSV2
****Sub-Circuit for OA21HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA21HSV4 A1 A2 B Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=860.00n L=60.00n
MM2 net064 B net029 VPW N12LL W=350.00n L=60.00n
MM1 net029 A1 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net029 A2 VSS VPW N12LL W=350.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net064 B VDD VNW P12LL W=520.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=520.00n L=60.00n
.ENDS OA21HSV4
****Sub-Circuit for OA221HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA221HSV0 A1 A2 B1 B2 C Z VDD VSS
MM9 net18 B2 net030 VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=200.00n L=60.00n
MM2 net18 B1 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 C VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=300.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM5 net064 C VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA221HSV0
****Sub-Circuit for OA221HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA221HSV1 A1 A2 B1 B2 C Z VDD VSS
MM9 net18 B2 net030 VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=290.00n L=60.00n
MM2 net18 B1 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 C VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=440.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM5 net064 C VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA221HSV1
****Sub-Circuit for OA221HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA221HSV2 A1 A2 B1 B2 C Z VDD VSS
MM9 net18 B2 net030 VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=430.00n L=60.00n
MM2 net18 B1 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 C VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=650.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM5 net064 C VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA221HSV2
****Sub-Circuit for OA221HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA221HSV4 A1 A2 B1 B2 C Z VDD VSS
MM9 net18 B2 net030 VPW N12LL W=350.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=860.00n L=60.00n
MM2 net18 B1 net030 VPW N12LL W=350.00n L=60.00n
MM3 net030 C VSS VPW N12LL W=350.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=350.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=350.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=520.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net064 B1 net071 VNW P12LL W=520.00n L=60.00n
MM5 net064 C VDD VNW P12LL W=520.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=520.00n L=60.00n
.ENDS OA221HSV4
****Sub-Circuit for OA222HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA222HSV0 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM12 net030 B2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net18 C2 net030 VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=200.00n L=60.00n
MM2 net18 C1 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM10 net073 C2 VDD VNW P12LL W=300.00n L=60.00n
MM11 net064 C1 net073 VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=300.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA222HSV0
****Sub-Circuit for OA222HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA222HSV1 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM12 net030 B2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net18 C2 net030 VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=290.00n L=60.00n
MM2 net18 C1 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM10 net073 C2 VDD VNW P12LL W=300.00n L=60.00n
MM11 net064 C1 net073 VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=440.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA222HSV1
****Sub-Circuit for OA222HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA222HSV2 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM12 net030 B2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net18 C2 net030 VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=430.00n L=60.00n
MM2 net18 C1 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM10 net073 C2 VDD VNW P12LL W=300.00n L=60.00n
MM11 net064 C1 net073 VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=650.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA222HSV2
****Sub-Circuit for OA222HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA222HSV4 A1 A2 B1 B2 C1 C2 Z VDD VSS
MM12 net030 B2 VSS VPW N12LL W=350.00n L=60.00n
MM9 net18 C2 net030 VPW N12LL W=350.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=860.00n L=60.00n
MM2 net18 C1 net030 VPW N12LL W=350.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=350.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=350.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=350.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=520.00n L=60.00n
MM10 net073 C2 VDD VNW P12LL W=520.00n L=60.00n
MM11 net064 C1 net073 VNW P12LL W=520.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net064 B1 net071 VNW P12LL W=520.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=520.00n L=60.00n
.ENDS OA222HSV4
****Sub-Circuit for OA22HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA22HSV0 A1 A2 B1 B2 Z VDD VSS
MM9 net18 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=200.00n L=60.00n
MM2 net18 B1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=300.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA22HSV0
****Sub-Circuit for OA22HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA22HSV1 A1 A2 B1 B2 Z VDD VSS
MM9 net18 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=290.00n L=60.00n
MM2 net18 B1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=440.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA22HSV1
****Sub-Circuit for OA22HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA22HSV2 A1 A2 B1 B2 Z VDD VSS
MM9 net18 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=430.00n L=60.00n
MM2 net18 B1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=650.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA22HSV2
****Sub-Circuit for OA22HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA22HSV4 A1 A2 B1 B2 Z VDD VSS
MM9 net18 B2 VSS VPW N12LL W=350.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=860.00n L=60.00n
MM2 net18 B1 VSS VPW N12LL W=350.00n L=60.00n
MM1 net064 A1 net18 VPW N12LL W=350.00n L=60.00n
MMN1 net064 A2 net18 VPW N12LL W=350.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=520.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net064 B1 net071 VNW P12LL W=520.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=520.00n L=60.00n
.ENDS OA22HSV4
****Sub-Circuit for OA31HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA31HSV0 A1 A2 A3 B Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=200.00n L=60.00n
MM2 net041 B VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=300.00n L=60.00n
MM4 net064 B VDD VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA31HSV0
****Sub-Circuit for OA31HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA31HSV1 A1 A2 A3 B Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=290.0n L=60.00n
MM2 net041 B VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=440.00n L=60.00n
MM4 net064 B VDD VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA31HSV1
****Sub-Circuit for OA31HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA31HSV2 A1 A2 A3 B Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=430.0n L=60.00n
MM2 net041 B VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=650.00n L=60.00n
MM4 net064 B VDD VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA31HSV2
****Sub-Circuit for OA31HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA31HSV4 A1 A2 A3 B Z VDD VSS
MM7 Z net064 VSS VPW N12LL W=860.00n L=60.00n
MM2 net041 B VSS VPW N12LL W=350.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=350.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=350.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=350.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net064 B VDD VNW P12LL W=520.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=520.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=520.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=520.00n L=60.00n
.ENDS OA31HSV4
****Sub-Circuit for OA32HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA32HSV0 A1 A2 A3 B1 B2 Z VDD VSS
MM11 net041 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=200.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=300.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA32HSV0
****Sub-Circuit for OA32HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA32HSV1 A1 A2 A3 B1 B2 Z VDD VSS
MM11 net041 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=290.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=440.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA32HSV1
****Sub-Circuit for OA32HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA32HSV2 A1 A2 A3 B1 B2 Z VDD VSS
MM11 net041 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=430.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=200.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=650.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA32HSV2
****Sub-Circuit for OA32HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA32HSV4 A1 A2 A3 B1 B2 Z VDD VSS
MM11 net041 B2 VSS VPW N12LL W=350.0n L=60.00n
MM7 Z net064 VSS VPW N12LL W=860.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=350.0n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=350.0n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=350.0n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=350.0n L=60.00n
MM6 Z net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net064 B1 net071 VNW P12LL W=520.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=520.00n L=60.00n
MM10 net071 B2 VDD VNW P12LL W=520.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=520.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=520.00n L=60.00n
.ENDS OA32HSV4
****Sub-Circuit for OA33HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA33HSV0 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM11 net041 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=200.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=200.00n L=60.00n
MM13 net041 B3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=200.00n L=60.00n
MM12 net076 B3 VDD VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=300.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net071 B2 net076 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA33HSV0
****Sub-Circuit for OA33HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA33HSV1 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM11 net041 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=290.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=200.00n L=60.00n
MM13 net041 B3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=200.00n L=60.00n
MM12 net076 B3 VDD VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=440.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net071 B2 net076 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA33HSV1
****Sub-Circuit for OA33HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA33HSV2 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM11 net041 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=430.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=200.00n L=60.00n
MM13 net041 B3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=200.00n L=60.00n
MM12 net076 B3 VDD VNW P12LL W=300.00n L=60.00n
MM6 Z net064 VDD VNW P12LL W=650.00n L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net071 B2 net076 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OA33HSV2
****Sub-Circuit for OA33HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OA33HSV4 A1 A2 A3 B1 B2 B3 Z VDD VSS
MM11 net041 B2 VSS VPW N12LL W=350.00n L=60.00n
MM7 Z net064 VSS VPW N12LL W=860.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=350.00n L=60.00n
MM9 net064 A3 net041 VPW N12LL W=350.00n L=60.00n
MM1 net064 A1 net041 VPW N12LL W=350.00n L=60.00n
MM13 net041 B3 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net064 A2 net041 VPW N12LL W=350.00n L=60.00n
MM12 net076 B3 VDD VNW P12LL W=520.0n L=60.00n
MM6 Z net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net064 B1 net071 VNW P12LL W=520.0n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=520.0n L=60.00n
MM10 net071 B2 net076 VNW P12LL W=520.0n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=520.0n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=520.0n L=60.00n
.ENDS OA33HSV4
****Sub-Circuit for OAI211HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI211HSV0 A1 A2 B C ZN VDD VSS
MM2 ZN B net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 C net027 VPW N12LL W=200.00n L=60.00n
MM1 net027 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net027 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=300.00n L=60.00n
MM5 ZN C VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI211HSV0
****Sub-Circuit for OAI211HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI211HSV1 A1 A2 B C ZN VDD VSS
MM2 ZN B net030 VPW N12LL W=290.00n L=60.00n
MM3 net030 C net027 VPW N12LL W=290.00n L=60.00n
MM1 net027 A1 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net027 A2 VSS VPW N12LL W=290.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=440.00n L=60.00n
MM5 ZN C VDD VNW P12LL W=440.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=440.00n L=60.00n
.ENDS OAI211HSV1
****Sub-Circuit for OAI211HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI211HSV2 A1 A2 B C ZN VDD VSS
MM2 ZN B net030 VPW N12LL W=430.00n L=60.00n
MM3 net030 C net027 VPW N12LL W=430.00n L=60.00n
MM1 net027 A1 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net027 A2 VSS VPW N12LL W=430.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=650.00n L=60.00n
MM5 ZN C VDD VNW P12LL W=650.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=650.00n L=60.00n
.ENDS OAI211HSV2
****Sub-Circuit for OAI211HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI211HSV4 A1 A2 B C ZN VDD VSS
MM7 ZN net064 VSS VPW N12LL W=860.00n L=60.00n
MM8 net064 net079 VSS VPW N12LL W=350.00n L=60.00n
MM2 net079 B net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 C net044 VPW N12LL W=200.00n L=60.00n
MM1 net044 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net044 A2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net064 net079 VDD VNW P12LL W=530.00n L=60.00n
MM6 ZN net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net079 B VDD VNW P12LL W=300.00n L=60.00n
MM5 net079 C VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net079 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI211HSV4
****Sub-Circuit for OAI21HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI21HSV0 A1 A2 B ZN VDD VSS
MM2 ZN B net029 VPW N12LL W=200.00n L=60.00n
MM1 net029 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net029 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI21HSV0
****Sub-Circuit for OAI21HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI21HSV1 A1 A2 B ZN VDD VSS
MM2 ZN B net029 VPW N12LL W=290.00n L=60.00n
MM1 net029 A1 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net029 A2 VSS VPW N12LL W=290.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=440.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=440.00n L=60.00n
.ENDS OAI21HSV1
****Sub-Circuit for OAI21HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI21HSV2 A1 A2 B ZN VDD VSS
MM2 ZN B net029 VPW N12LL W=430.00n L=60.00n
MM1 net029 A1 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net029 A2 VSS VPW N12LL W=430.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=650.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=650.00n L=60.00n
.ENDS OAI21HSV2
****Sub-Circuit for OAI21HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI21HSV4 A1 A2 B ZN VDD VSS
MM2 ZN B net029 VPW N12LL W=860.00n L=60.00n
MM1 net029 A1 VSS VPW N12LL W=860.00n L=60.00n
MMN1 net029 A2 VSS VPW N12LL W=860.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=1.3u L=60.00n
MM0 net067 A2 VDD VNW P12LL W=1.3u L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=1.3u L=60.00n
.ENDS OAI21HSV4
****Sub-Circuit for OAI221HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI221HSV0 A1 A2 B1 B2 C ZN VDD VSS
MM9 net18 B2 VSS VPW N12LL W=200.00n L=60.00n
MM2 net18 B1 VSS VPW N12LL W=200.00n L=60.00n
MM3 ZN C net045 VPW N12LL W=200.00n L=60.00n
MM1 net045 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net045 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.000n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=300.000n L=60.00n
MM5 ZN C VDD VNW P12LL W=300.000n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.000n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=300.000n L=60.00n
.ENDS OAI221HSV0
****Sub-Circuit for OAI221HSV1, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT OAI221HSV1 A1 A2 B1 B2 C ZN VDD VSS
MM9 net18 B2 VSS VPW N12LL W=275.00n L=60.00n
MM2 net18 B1 VSS VPW N12LL W=290.00n L=60.00n
MM3 ZN C net045 VPW N12LL W=290.00n L=60.00n
MM1 net045 A1 net18 VPW N12LL W=290.00n L=60.00n
MMN1 net045 A2 net18 VPW N12LL W=290.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=425.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=440.00n L=60.00n
MM5 ZN C VDD VNW P12LL W=440.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=440.00n L=60.00n
.ENDS OAI221HSV1
****Sub-Circuit for OAI221HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI221HSV2 A1 A2 B1 B2 C ZN VDD VSS
MM9 net18 B2 VSS VPW N12LL W=430.00n L=60.00n
MM2 net18 B1 VSS VPW N12LL W=430.00n L=60.00n
MM3 ZN C net045 VPW N12LL W=430.00n L=60.00n
MM1 net045 A1 net18 VPW N12LL W=430.00n L=60.00n
MMN1 net045 A2 net18 VPW N12LL W=430.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=640.0n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=640.0n L=60.00n
MM5 ZN C VDD VNW P12LL W=640.0n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=640.0n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=640.0n L=60.00n
.ENDS OAI221HSV2
****Sub-Circuit for OAI221HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI221HSV4 A1 A2 B1 B2 C ZN VDD VSS
MM9 net18 B2 VSS VPW N12LL W=200.00n L=60.00n
MM7 ZN net064 VSS VPW N12LL W=860.00n L=60.00n
MM10 net064 net093 VSS VPW N12LL W=350.00n L=60.00n
MM2 net18 B1 VSS VPW N12LL W=200.00n L=60.00n
MM3 net093 C net062 VPW N12LL W=200.00n L=60.00n
MM1 net062 A1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net062 A2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM6 ZN net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net093 B1 net071 VNW P12LL W=300.00n L=60.00n
MM5 net093 C VDD VNW P12LL W=300.00n L=60.00n
MM11 net064 net093 VDD VNW P12LL W=530.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net093 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI221HSV4
****Sub-Circuit for OAI222HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI222HSV0 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM12 net030 B2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net18 A2 net030 VPW N12LL W=200.00n L=60.00n
MM2 net18 A1 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=200.00n L=60.00n
MM1 ZN C1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 ZN C2 net18 VPW N12LL W=200.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM10 net073 C2 VDD VNW P12LL W=300.00n L=60.00n
MM11 ZN C1 net073 VNW P12LL W=300.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI222HSV0
****Sub-Circuit for OAI222HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI222HSV1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM12 net030 B2 VSS VPW N12LL W=290.00n L=60.00n
MM9 net18 A2 net030 VPW N12LL W=290.00n L=60.00n
MM2 net18 A1 net030 VPW N12LL W=290.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=290.00n L=60.00n
MM1 ZN C1 net18 VPW N12LL W=290.00n L=60.00n
MMN1 ZN C2 net18 VPW N12LL W=290.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=440.00n L=60.00n
MM10 net073 C2 VDD VNW P12LL W=440.00n L=60.00n
MM11 ZN C1 net073 VNW P12LL W=440.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=440.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=440.00n L=60.00n
.ENDS OAI222HSV1
****Sub-Circuit for OAI222HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI222HSV2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM12 net030 B2 VSS VPW N12LL W=430.00n L=60.00n
MM9 net18 A2 net030 VPW N12LL W=430.00n L=60.00n
MM2 net18 A1 net030 VPW N12LL W=430.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=430.00n L=60.00n
MM1 ZN C1 net18 VPW N12LL W=430.00n L=60.00n
MMN1 ZN C2 net18 VPW N12LL W=430.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=650.00n L=60.00n
MM10 net073 C2 VDD VNW P12LL W=650.00n L=60.00n
MM11 ZN C1 net073 VNW P12LL W=650.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=650.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=650.00n L=60.00n
.ENDS OAI222HSV2
****Sub-Circuit for OAI222HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI222HSV4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
MM12 net030 B2 VSS VPW N12LL W=200.00n L=60.00n
MM9 net18 A2 net030 VPW N12LL W=200.00n L=60.00n
MM7 ZN net051 VSS VPW N12LL W=860.00n L=60.00n
MM2 net18 A1 net030 VPW N12LL W=200.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=200.00n L=60.00n
MM13 net051 net064 VSS VPW N12LL W=350.00n L=60.00n
MM1 net064 C1 net18 VPW N12LL W=200.00n L=60.00n
MMN1 net064 C2 net18 VPW N12LL W=200.00n L=60.00n
MM14 net051 net064 VDD VNW P12LL W=530.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM10 net073 C2 VDD VNW P12LL W=300.00n L=60.00n
MM11 net064 C1 net073 VNW P12LL W=300.00n L=60.00n
MM6 ZN net051 VDD VNW P12LL W=1.3u L=60.00n
MM4 net064 B1 net071 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net064 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI222HSV4
****Sub-Circuit for OAI22HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI22HSV0 A1 A2 B1 B2 ZN VDD VSS
MM12 net030 B2 VSS VPW N12LL W=200.0n L=60.00n
MM9 ZN A2 net030 VPW N12LL W=200.0n L=60.00n
MM2 ZN A1 net030 VPW N12LL W=200.0n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=200.0n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=300.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI22HSV0
****Sub-Circuit for OAI22HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI22HSV1 A1 A2 B1 B2 ZN VDD VSS
MM12 net030 B2 VSS VPW N12LL W=290.00n L=60.00n
MM9 ZN A2 net030 VPW N12LL W=290.00n L=60.00n
MM2 ZN A1 net030 VPW N12LL W=290.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=255.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=440.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=405.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=440.00n L=60.00n
.ENDS OAI22HSV1
****Sub-Circuit for OAI22HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI22HSV2 A1 A2 B1 B2 ZN VDD VSS
MM12 net030 B2 VSS VPW N12LL W=430.00n L=60.00n
MM9 ZN A2 net030 VPW N12LL W=430.00n L=60.00n
MM2 ZN A1 net030 VPW N12LL W=430.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=430.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=650.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=650.00n L=60.00n
MM0 net067 A2 VDD VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=650.00n L=60.00n
.ENDS OAI22HSV2
****Sub-Circuit for OAI22HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI22HSV4 A1 A2 B1 B2 ZN VDD VSS
MM12 net030 B2 VSS VPW N12LL W=860.00n L=60.00n
MM9 ZN A2 net030 VPW N12LL W=860.00n L=60.00n
MM2 ZN A1 net030 VPW N12LL W=860.00n L=60.00n
MM3 net030 B1 VSS VPW N12LL W=860.00n L=60.00n
MM8 net071 B2 VDD VNW P12LL W=1.3u L=60.00n
MM4 ZN B1 net071 VNW P12LL W=1.3u L=60.00n
MM0 net067 A2 VDD VNW P12LL W=1.3u L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=1.3u L=60.00n
.ENDS OAI22HSV4
****Sub-Circuit for OAI31HSV0, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI31HSV0 A1 A2 A3 B ZN VDD VSS
MM2 ZN B net064 VPW N12LL W=200.00n L=60.00n
MM9 net064 A3 VSS VPW N12LL W=200.00n L=60.00n
MM1 net064 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net064 A2 VSS VPW N12LL W=200.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI31HSV0
****Sub-Circuit for OAI31HSV1, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI31HSV1 A1 A2 A3 B ZN VDD VSS
MM2 ZN B net064 VPW N12LL W=290.00n L=60.00n
MM9 net064 A3 VSS VPW N12LL W=290.00n L=60.00n
MM1 net064 A1 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net064 A2 VSS VPW N12LL W=290.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=440.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=440.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=440.00n L=60.00n
.ENDS OAI31HSV1
****Sub-Circuit for OAI31HSV2, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI31HSV2 A1 A2 A3 B ZN VDD VSS
MM2 ZN B net064 VPW N12LL W=430.00n L=60.00n
MM9 net064 A3 VSS VPW N12LL W=430.00n L=60.00n
MM1 net064 A1 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net064 A2 VSS VPW N12LL W=430.00n L=60.00n
MM4 ZN B VDD VNW P12LL W=650.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=650.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=650.00n L=60.00n
.ENDS OAI31HSV2
****Sub-Circuit for OAI31HSV4, Wed Dec  8 11:21:17 CST 2010****
.SUBCKT OAI31HSV4 A1 A2 A3 B ZN VDD VSS
MM7 ZN net064 VSS VPW N12LL W=860.00n L=60.00n
MM10 net064 net055 VSS VPW N12LL W=350.00n L=60.00n
MM2 net055 B net058 VPW N12LL W=200.00n L=60.00n
MM9 net058 A3 VSS VPW N12LL W=200.00n L=60.00n
MM1 net058 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net058 A2 VSS VPW N12LL W=200.00n L=60.00n
MM11 net064 net055 VDD VNW P12LL W=530.00n L=60.00n
MM6 ZN net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net055 B VDD VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net055 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI31HSV4
****Sub-Circuit for OAI32HSV0, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OAI32HSV0 A1 A2 A3 B1 B2 ZN VDD VSS
MM11 net041 B2 VSS VPW N12LL W=200.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=200.00n L=60.00n
MM9 ZN A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 ZN A1 net041 VPW N12LL W=200.00n L=60.00n
MMN1 ZN A2 net041 VPW N12LL W=200.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=300.0n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.0n L=60.00n
MM10 net071 B2 VDD VNW P12LL W=300.0n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.0n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=300.0n L=60.00n
.ENDS OAI32HSV0
****Sub-Circuit for OAI32HSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OAI32HSV1 A1 A2 A3 B1 B2 ZN VDD VSS
MM11 net041 B2 VSS VPW N12LL W=290.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=290.00n L=60.00n
MM9 ZN A3 net041 VPW N12LL W=290.00n L=60.00n
MM1 ZN A1 net041 VPW N12LL W=290.00n L=60.00n
MMN1 ZN A2 net041 VPW N12LL W=290.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=440.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=440.00n L=60.00n
MM10 net071 B2 VDD VNW P12LL W=440.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=440.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=440.00n L=60.00n
.ENDS OAI32HSV1
****Sub-Circuit for OAI32HSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OAI32HSV2 A1 A2 A3 B1 B2 ZN VDD VSS
MM11 net041 B2 VSS VPW N12LL W=430.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=430.00n L=60.00n
MM9 ZN A3 net041 VPW N12LL W=430.00n L=60.00n
MM1 ZN A1 net041 VPW N12LL W=430.00n L=60.00n
MMN1 ZN A2 net041 VPW N12LL W=430.00n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=650.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=650.00n L=60.00n
MM10 net071 B2 VDD VNW P12LL W=650.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=650.00n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=650.00n L=60.00n
.ENDS OAI32HSV2
****Sub-Circuit for OAI32HSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OAI32HSV4 A1 A2 A3 B1 B2 ZN VDD VSS
MM11 net041 B2 VSS VPW N12LL W=200.00n L=60.00n
MM12 net064 net0104 VSS VPW N12LL W=350.00n L=60.00n
MM7 ZN net064 VSS VPW N12LL W=860.00n L=60.00n
MM2 net041 B1 VSS VPW N12LL W=200.00n L=60.00n
MM9 net0104 A3 net041 VPW N12LL W=200.00n L=60.00n
MM1 net0104 A1 net041 VPW N12LL W=200.00n L=60.00n
MMN1 net0104 A2 net041 VPW N12LL W=200.00n L=60.00n
MM13 net064 net0104 VDD VNW P12LL W=530.00n L=60.00n
MM6 ZN net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net0104 B1 net071 VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net071 B2 VDD VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net0104 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI32HSV4
****Sub-Circuit for OAI33HSV0, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OAI33HSV0 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM11 net041 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 net041 A1 VSS VPW N12LL W=200.00n L=60.00n
MM9 ZN B3 net041 VPW N12LL W=200.00n L=60.00n
MM1 ZN B1 net041 VPW N12LL W=200.00n L=60.00n
MM13 net041 A3 VSS VPW N12LL W=200.00n L=60.00n
MMN1 ZN B2 net041 VPW N12LL W=200.00n L=60.00n
MM12 net076 B3 VDD VNW P12LL W=300.0n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=300.0n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.0n L=60.00n
MM10 net071 B2 net076 VNW P12LL W=300.0n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.0n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=300.0n L=60.00n
.ENDS OAI33HSV0
****Sub-Circuit for OAI33HSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OAI33HSV1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM11 net041 A2 VSS VPW N12LL W=290.00n L=60.00n
MM2 net041 A1 VSS VPW N12LL W=290.00n L=60.00n
MM9 ZN B3 net041 VPW N12LL W=290.00n L=60.00n
MM1 ZN B1 net041 VPW N12LL W=290.00n L=60.00n
MM13 net041 A3 VSS VPW N12LL W=290.00n L=60.00n
MMN1 ZN B2 net041 VPW N12LL W=290.00n L=60.00n
MM12 net076 B3 VDD VNW P12LL W=440.0n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=440.0n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=440.0n L=60.00n
MM10 net071 B2 net076 VNW P12LL W=440.0n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=440.0n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=440.0n L=60.00n
.ENDS OAI33HSV1
****Sub-Circuit for OAI33HSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OAI33HSV2 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM11 net041 A2 VSS VPW N12LL W=430.00n L=60.00n
MM2 net041 A1 VSS VPW N12LL W=430.00n L=60.00n
MM9 ZN B3 net041 VPW N12LL W=430.00n L=60.00n
MM1 ZN B1 net041 VPW N12LL W=430.00n L=60.00n
MM13 net041 A3 VSS VPW N12LL W=430.00n L=60.00n
MMN1 ZN B2 net041 VPW N12LL W=430.00n L=60.00n
MM12 net076 B3 VDD VNW P12LL W=650.0n L=60.00n
MM4 ZN B1 net071 VNW P12LL W=650.0n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=650.0n L=60.00n
MM10 net071 B2 net076 VNW P12LL W=650.0n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=650.0n L=60.00n
MMP1 ZN A1 net067 VNW P12LL W=650.0n L=60.00n
.ENDS OAI33HSV2
****Sub-Circuit for OAI33HSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OAI33HSV4 A1 A2 A3 B1 B2 B3 ZN VDD VSS
MM11 net041 B2 net077 VPW N12LL W=200.0n L=60.00n
MM7 ZN net064 VSS VPW N12LL W=860.00n L=60.00n
MM14 net064 net041 VSS VPW N12LL W=350.00n L=60.00n
MM2 net041 B1 net077 VPW N12LL W=200.0n L=60.00n
MM9 net077 A3 VSS VPW N12LL W=200.0n L=60.00n
MM1 net077 A1 VSS VPW N12LL W=200.0n L=60.00n
MM13 net041 B3 net077 VPW N12LL W=200.0n L=60.00n
MMN1 net077 A2 VSS VPW N12LL W=200.0n L=60.00n
MM12 net076 B3 VDD VNW P12LL W=300.00n L=60.00n
MM15 net064 net041 VDD VNW P12LL W=530.00n L=60.00n
MM6 ZN net064 VDD VNW P12LL W=1.3u L=60.00n
MM4 net041 B1 net071 VNW P12LL W=300.00n L=60.00n
MM8 net065 A3 VDD VNW P12LL W=300.00n L=60.00n
MM10 net071 B2 net076 VNW P12LL W=300.00n L=60.00n
MM0 net067 A2 net065 VNW P12LL W=300.00n L=60.00n
MMP1 net041 A1 net067 VNW P12LL W=300.00n L=60.00n
.ENDS OAI33HSV4
****Sub-Circuit for OAO211HSV0, Thu May 19 13:57:40 CST 2011****
.SUBCKT OAO211HSV0 A1 A2 B C Z VDD VSS
MM7 Z net18 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net14 A2 VSS VPW N12LL W=180.00n L=60.00n
MM1 net14 A1 VSS VPW N12LL W=180.00n L=60.00n
MM2 net18 B net14 VPW N12LL W=180.00n L=60.00n
MM5 net18 C VSS VPW N12LL W=180.00n L=60.00n
MM6 Z net18 VDD VNW P12LL W=250.00n L=60.00n
MMP1 net30 A1 net33 VNW P12LL W=200.00n L=60.00n
MM0 net33 A2 VDD VNW P12LL W=200.00n L=60.00n
MM4 net30 B VDD VNW P12LL W=200.00n L=60.00n
MM3 net18 C net30 VNW P12LL W=200.00n L=60.00n
.ENDS OAO211HSV0
****Sub-Circuit for OAO211HSV1, Thu May 19 13:57:40 CST 2011****
.SUBCKT OAO211HSV1 A1 A2 B C Z VDD VSS
MM6 Z net30 VDD VNW P12LL W=440.00n L=60.00n
MMP1 net18 A1 net21 VNW P12LL W=200.00n L=60.00n
MM0 net21 A2 VDD VNW P12LL W=200.00n L=60.00n
MM4 net18 B VDD VNW P12LL W=200.00n L=60.00n
MM3 net30 C net18 VNW P12LL W=200.00n L=60.00n
MM7 Z net30 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net34 A2 VSS VPW N12LL W=180.00n L=60.00n
MM1 net34 A1 VSS VPW N12LL W=180.00n L=60.00n
MM2 net30 B net34 VPW N12LL W=180.00n L=60.00n
MM5 net30 C VSS VPW N12LL W=180.00n L=60.00n
.ENDS OAO211HSV1
****Sub-Circuit for OAO211HSV2, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAO211HSV2 A1 A2 B C Z VDD VSS
MM3 net30 C net18 VNW P12LL W=220.00n L=60.00n
MM4 net18 B VDD VNW P12LL W=220.00n L=60.00n
MM0 net21 A2 VDD VNW P12LL W=220.00n L=60.00n
MMP1 net18 A1 net21 VNW P12LL W=220.00n L=60.00n
MM6 Z net30 VDD VNW P12LL W=540.00n L=60.00n
MM5 net30 C VSS VPW N12LL W=180.00n L=60.00n
MM2 net30 B net34 VPW N12LL W=180.00n L=60.00n
MM1 net34 A1 VSS VPW N12LL W=180.00n L=60.00n
MMN1 net34 A2 VSS VPW N12LL W=180.00n L=60.00n
MM7 Z net30 VSS VPW N12LL W=430.00n L=60.00n
.ENDS OAO211HSV2
****Sub-Circuit for OAO211HSV4, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAO211HSV4 A1 A2 B C Z VDD VSS
MM3 net30 C net18 VNW P12LL W=440.00n L=60.00n
MM4 net18 B VDD VNW P12LL W=440.00n L=60.00n
MM0 net21 A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 net18 A1 net21 VNW P12LL W=440.00n L=60.00n
MM6 Z net30 VDD VNW P12LL W=1.08u L=60.00n
MM5 net30 C VSS VPW N12LL W=350.00n L=60.00n
MM2 net30 B net34 VPW N12LL W=350.00n L=60.00n
MM1 net34 A1 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net34 A2 VSS VPW N12LL W=350.00n L=60.00n
MM7 Z net30 VSS VPW N12LL W=860.00n L=60.00n
.ENDS OAO211HSV4
****Sub-Circuit for OAOAI2111HSV0, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOAI2111HSV0 A1 A2 B C D ZN VDD VSS
MM7 ZN D net19 VPW N12LL W=200.00n L=60.00n
MMN1 net15 A2 VSS VPW N12LL W=200.00n L=60.00n
MM1 net15 A1 VSS VPW N12LL W=200.00n L=60.00n
MM2 net19 B net15 VPW N12LL W=200.00n L=60.00n
MM5 net19 C VSS VPW N12LL W=200.00n L=60.00n
MM6 ZN D VDD VNW P12LL W=250.00n L=60.00n
MMP1 net31 A1 net34 VNW P12LL W=250.00n L=60.00n
MM0 net34 A2 VDD VNW P12LL W=250.00n L=60.00n
MM4 net31 B VDD VNW P12LL W=250.00n L=60.00n
MM3 ZN C net31 VNW P12LL W=250.00n L=60.00n
.ENDS OAOAI2111HSV0
****Sub-Circuit for OAOAI2111HSV1, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOAI2111HSV1 A1 A2 B C D ZN VDD VSS
MM3 ZN C net19 VNW P12LL W=440.00n L=60.00n
MM4 net19 B VDD VNW P12LL W=440.00n L=60.00n
MM0 net22 A2 VDD VNW P12LL W=440.00n L=60.00n
MMP1 net19 A1 net22 VNW P12LL W=440.00n L=60.00n
MM6 ZN D VDD VNW P12LL W=440.00n L=60.00n
MM5 net31 C VSS VPW N12LL W=350.00n L=60.00n
MM2 net31 B net35 VPW N12LL W=350.00n L=60.00n
MM1 net35 A1 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net35 A2 VSS VPW N12LL W=350.00n L=60.00n
MM7 ZN D net31 VPW N12LL W=350.00n L=60.00n
.ENDS OAOAI2111HSV1
****Sub-Circuit for OAOAI2111HSV2, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOAI2111HSV2 A1 A2 B C D ZN VDD VSS
MM3 ZN C net19 VNW P12LL W=540.00n L=60.00n
MM4 net19 B VDD VNW P12LL W=540.00n L=60.00n
MM0 net22 A2 VDD VNW P12LL W=540.00n L=60.00n
MMP1 net19 A1 net22 VNW P12LL W=540.00n L=60.00n
MM6 ZN D VDD VNW P12LL W=540.00n L=60.00n
MM5 net31 C VSS VPW N12LL W=430.00n L=60.00n
MM2 net31 B net35 VPW N12LL W=430.00n L=60.00n
MM1 net35 A1 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net35 A2 VSS VPW N12LL W=430.00n L=60.00n
MM7 ZN D net31 VPW N12LL W=430.00n L=60.00n
.ENDS OAOAI2111HSV2
****Sub-Circuit for OAOAI2111HSV4, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOAI2111HSV4 A1 A2 B C D ZN VDD VSS
MM3 ZN C net19 VNW P12LL W=1.08u L=60.00n
MM4 net19 B VDD VNW P12LL W=1.08u L=60.00n
MM0 net22 A2 VDD VNW P12LL W=1.08u L=60.00n
MMP1 net19 A1 net22 VNW P12LL W=1.08u L=60.00n
MM6 ZN D VDD VNW P12LL W=1.08u L=60.00n
MM5 net31 C VSS VPW N12LL W=860.00n L=60.00n
MM2 net31 B net35 VPW N12LL W=860.00n L=60.00n
MM1 net35 A1 VSS VPW N12LL W=860.00n L=60.00n
MMN1 net35 A2 VSS VPW N12LL W=860.00n L=60.00n
MM7 ZN D net31 VPW N12LL W=860.00n L=60.00n
.ENDS OAOAI2111HSV4
****Sub-Circuit for OAOAOAI211111HSV0, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOAOAI211111HSV0 A1 A2 B C D E F ZN VDD VSS
MM9 ZN F VDD VNW P12LL W=250.00n L=60.00n
MM8 ZN E net14 VNW P12LL W=250.00n L=60.00n
MM3 net14 C net27 VNW P12LL W=250.00n L=60.00n
MM4 net27 B VDD VNW P12LL W=250.00n L=60.00n
MM0 net30 A2 VDD VNW P12LL W=250.00n L=60.00n
MMP1 net27 A1 net30 VNW P12LL W=250.00n L=60.00n
MM6 net14 D VDD VNW P12LL W=250.00n L=60.00n
MM11 ZN F net59 VPW N12LL W=200.00n L=60.00n
MM10 net59 E VSS VPW N12LL W=200.00n L=60.00n
MM5 net47 C VSS VPW N12LL W=200.00n L=60.00n
MM2 net47 B net51 VPW N12LL W=200.00n L=60.00n
MM1 net51 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net51 A2 VSS VPW N12LL W=200.00n L=60.00n
MM7 net59 D net47 VPW N12LL W=200.00n L=60.00n
.ENDS OAOAOAI211111HSV0
****Sub-Circuit for OAOAOAI211111HSV1, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOAOAI211111HSV1 A1 A2 B C D E F ZN VDD VSS
MM7 net9 D net21 VPW N12LL W=350.00n L=60.00n
MMN1 net17 A2 VSS VPW N12LL W=350.00n L=60.00n
MM1 net17 A1 VSS VPW N12LL W=350.00n L=60.00n
MM2 net21 B net17 VPW N12LL W=350.00n L=60.00n
MM5 net21 C VSS VPW N12LL W=350.00n L=60.00n
MM10 net9 E VSS VPW N12LL W=350.00n L=60.00n
MM11 ZN F net9 VPW N12LL W=350.00n L=60.00n
MM6 net60 D VDD VNW P12LL W=440.00n L=60.00n
MMP1 net41 A1 net44 VNW P12LL W=440.00n L=60.00n
MM0 net44 A2 VDD VNW P12LL W=440.00n L=60.00n
MM4 net41 B VDD VNW P12LL W=440.00n L=60.00n
MM3 net60 C net41 VNW P12LL W=440.00n L=60.00n
MM8 ZN E net60 VNW P12LL W=440.00n L=60.00n
MM9 ZN F VDD VNW P12LL W=440.00n L=60.00n
.ENDS OAOAOAI211111HSV1
****Sub-Circuit for OAOAOAI211111HSV2, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOAOAI211111HSV2 A1 A2 B C D E F ZN VDD VSS
MM7 net9 D net21 VPW N12LL W=430.00n L=60.00n
MMN1 net17 A2 VSS VPW N12LL W=430.00n L=60.00n
MM1 net17 A1 VSS VPW N12LL W=430.00n L=60.00n
MM2 net21 B net17 VPW N12LL W=430.00n L=60.00n
MM5 net21 C VSS VPW N12LL W=430.00n L=60.00n
MM10 net9 E VSS VPW N12LL W=430.00n L=60.00n
MM11 ZN F net9 VPW N12LL W=430.00n L=60.00n
MM6 net60 D VDD VNW P12LL W=540.00n L=60.00n
MMP1 net41 A1 net44 VNW P12LL W=540.00n L=60.00n
MM0 net44 A2 VDD VNW P12LL W=540.00n L=60.00n
MM4 net41 B VDD VNW P12LL W=540.00n L=60.00n
MM3 net60 C net41 VNW P12LL W=540.00n L=60.00n
MM8 ZN E net60 VNW P12LL W=540.00n L=60.00n
MM9 ZN F VDD VNW P12LL W=540.00n L=60.00n
.ENDS OAOAOAI211111HSV2
****Sub-Circuit for OAOAOAI211111HSV4, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOAOAI211111HSV4 A1 A2 B C D E F ZN VDD VSS
MM7 net9 D net21 VPW N12LL W=860.00n L=60.00n
MMN1 net17 A2 VSS VPW N12LL W=860.00n L=60.00n
MM1 net17 A1 VSS VPW N12LL W=860.00n L=60.00n
MM2 net21 B net17 VPW N12LL W=860.00n L=60.00n
MM5 net21 C VSS VPW N12LL W=860.00n L=60.00n
MM10 net9 E VSS VPW N12LL W=860.00n L=60.00n
MM11 ZN F net9 VPW N12LL W=860.00n L=60.00n
MM6 net60 D VDD VNW P12LL W=1.08u L=60.00n
MMP1 net41 A1 net44 VNW P12LL W=1.08u L=60.00n
MM0 net44 A2 VDD VNW P12LL W=1.08u L=60.00n
MM4 net41 B VDD VNW P12LL W=1.08u L=60.00n
MM3 net60 C net41 VNW P12LL W=1.08u L=60.00n
MM8 ZN E net60 VNW P12LL W=1.08u L=60.00n
MM9 ZN F VDD VNW P12LL W=1.08u L=60.00n
.ENDS OAOAOAI211111HSV4
****Sub-Circuit for OAOI211HSV0, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOI211HSV0 A1 A2 B C ZN VDD VSS
MM3 ZN C net18 VNW P12LL W=250.00n L=60.00n
MM4 net18 B VDD VNW P12LL W=250.00n L=60.00n
MM0 net21 A2 VDD VNW P12LL W=250.00n L=60.00n
MMP1 net18 A1 net21 VNW P12LL W=250.00n L=60.00n
MM5 ZN C VSS VPW N12LL W=200.00n L=60.00n
MM2 ZN B net30 VPW N12LL W=200.00n L=60.00n
MM1 net30 A1 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net30 A2 VSS VPW N12LL W=200.00n L=60.00n
.ENDS OAOI211HSV0
****Sub-Circuit for OAOI211HSV1, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOI211HSV1 A1 A2 B C ZN VDD VSS
MMN1 net10 A2 VSS VPW N12LL W=350.00n L=60.00n
MM1 net10 A1 VSS VPW N12LL W=350.00n L=60.00n
MM2 ZN B net10 VPW N12LL W=350.00n L=60.00n
MM5 ZN C VSS VPW N12LL W=350.00n L=60.00n
MMP1 net22 A1 net25 VNW P12LL W=440.00n L=60.00n
MM0 net25 A2 VDD VNW P12LL W=440.00n L=60.00n
MM4 net22 B VDD VNW P12LL W=440.00n L=60.00n
MM3 ZN C net22 VNW P12LL W=440.00n L=60.00n
.ENDS OAOI211HSV1
****Sub-Circuit for OAOI211HSV2, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOI211HSV2 A1 A2 B C ZN VDD VSS
MMN1 net10 A2 VSS VPW N12LL W=430.00n L=60.00n
MM1 net10 A1 VSS VPW N12LL W=430.00n L=60.00n
MM2 ZN B net10 VPW N12LL W=430.00n L=60.00n
MM5 ZN C VSS VPW N12LL W=430.00n L=60.00n
MMP1 net22 A1 net25 VNW P12LL W=540.00n L=60.00n
MM0 net25 A2 VDD VNW P12LL W=540.00n L=60.00n
MM4 net22 B VDD VNW P12LL W=540.00n L=60.00n
MM3 ZN C net22 VNW P12LL W=540.00n L=60.00n
.ENDS OAOI211HSV2
****Sub-Circuit for OAOI211HSV4, Fri Dec 24 10:49:43 CST 2010****
.SUBCKT OAOI211HSV4 A1 A2 B C ZN VDD VSS
MMN1 net10 A2 VSS VPW N12LL W=860.00n L=60.00n
MM1 net10 A1 VSS VPW N12LL W=860.00n L=60.00n
MM2 ZN B net10 VPW N12LL W=860.00n L=60.00n
MM5 ZN C VSS VPW N12LL W=860.00n L=60.00n
MMP1 net22 A1 net25 VNW P12LL W=1.08u L=60.00n
MM0 net25 A2 VDD VNW P12LL W=1.08u L=60.00n
MM4 net22 B VDD VNW P12LL W=1.08u L=60.00n
MM3 ZN C net22 VNW P12LL W=1.08u L=60.00n
.ENDS OAOI211HSV4
****Sub-Circuit for OR2HSV0, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR2HSV0 A1 A2 Z VDD VSS
MM0 net31 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=300.0n L=60.00n
MM4 Z net31 VDD VNW P12LL W=300.0n L=60.00n
MMP1 net42 A2 VDD VNW P12LL W=300.0n L=60.00n
.ENDS OR2HSV0
****Sub-Circuit for OR2HSV0RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR2HSV0RD A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=200.00n L=60.00n
MM0 net16 A2 VSS VPW N12LL W=180.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=270.0n L=60.00n
MM4 Z net16 VDD VNW P12LL W=250.0n L=60.00n
MM1 net16 A1 net15 VNW P12LL W=270.0n L=60.00n
.ENDS OR2HSV0RD
****Sub-Circuit for OR2HSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR2HSV1 A1 A2 Z VDD VSS
MM0 net31 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=300.0n L=60.00n
MM4 Z net31 VDD VNW P12LL W=440.0n L=60.00n
MMP1 net42 A2 VDD VNW P12LL W=300.0n L=60.00n
.ENDS OR2HSV1
****Sub-Circuit for OR2HSV12, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV12 A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=710.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=2.58u L=60.00n
MM0 net16 A2 VSS VPW N12LL W=710.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=1.30u L=60.00n
MM4 Z net16 VDD VNW P12LL W=3.24u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=1.30u L=60.00n
.ENDS OR2HSV12
****Sub-Circuit for OR2HSV12RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV12RD A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=1.13u L=60.00n
MM2 Z net16 VSS VPW N12LL W=2.58u L=60.00n
MM0 net16 A2 VSS VPW N12LL W=1.13u L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=2.06u L=60.00n
MM4 Z net16 VDD VNW P12LL W=3.24u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=2.05u L=60.00n
.ENDS OR2HSV12RD
****Sub-Circuit for OR2HSV12RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV12RQ A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=440.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=2.58u L=60.00n
MM0 net16 A2 VSS VPW N12LL W=440.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=810n L=60.00n
MM4 Z net16 VDD VNW P12LL W=3.24u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=810n L=60.00n
.ENDS OR2HSV12RQ
****Sub-Circuit for OR2HSV16, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV16 A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=950.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=3.44u L=60.00n
MM0 net16 A2 VSS VPW N12LL W=950.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=1.76u L=60.00n
MM4 Z net16 VDD VNW P12LL W=4.32u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=1.76u L=60.00n
.ENDS OR2HSV16
****Sub-Circuit for OR2HSV16RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV16RD A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=1.51u L=60.00n
MM2 Z net16 VSS VPW N12LL W=3.44u L=60.00n
MM0 net16 A2 VSS VPW N12LL W=1.51u L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=2.8u L=60.00n
MM4 Z net16 VDD VNW P12LL W=4.32u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=2.8u L=60.00n
.ENDS OR2HSV16RD
****Sub-Circuit for OR2HSV16RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV16RQ A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=580.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=3.44u L=60.00n
MM0 net16 A2 VSS VPW N12LL W=580.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=1.08u L=60.00n
MM4 Z net16 VDD VNW P12LL W=4.32u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=1.08u L=60.00n
.ENDS OR2HSV16RQ
****Sub-Circuit for OR2HSV1RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR2HSV1RD A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=350.00n L=60.00n
MM0 net16 A2 VSS VPW N12LL W=180.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=280.0n L=60.00n
MM4 Z net16 VDD VNW P12LL W=440.0n L=60.00n
MM1 net16 A1 net15 VNW P12LL W=280.0n L=60.00n
.ENDS OR2HSV1RD
****Sub-Circuit for OR2HSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR2HSV2 A1 A2 Z VDD VSS
MM0 net31 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=300.0n L=60.00n
MM4 Z net31 VDD VNW P12LL W=650.0n L=60.00n
MMP1 net42 A2 VDD VNW P12LL W=300.0n L=60.00n
.ENDS OR2HSV2
****Sub-Circuit for OR2HSV2RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV2RD A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=190.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=430.00n L=60.00n
MM0 net16 A2 VSS VPW N12LL W=190.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=350.0n L=60.00n
MM4 Z net16 VDD VNW P12LL W=540.0n L=60.00n
MM1 net16 A1 net15 VNW P12LL W=350.0n L=60.00n
.ENDS OR2HSV2RD
****Sub-Circuit for OR2HSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR2HSV4 A1 A2 Z VDD VSS
MM0 net31 A2 VSS VPW N12LL W=350.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=860.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=350.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=520.0n L=60.00n
MM4 Z net31 VDD VNW P12LL W=1.3u L=60.00n
MMP1 net42 A2 VDD VNW P12LL W=520.0n L=60.00n
.ENDS OR2HSV4
****Sub-Circuit for OR2HSV4RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV4RD A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=380.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=860.00n L=60.00n
MM0 net16 A2 VSS VPW N12LL W=380.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=650.0n L=60.00n
MM4 Z net16 VDD VNW P12LL W=1.08u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=650.0n L=60.00n
.ENDS OR2HSV4RD
****Sub-Circuit for OR2HSV4RQ, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR2HSV4RQ A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=860.00n L=60.00n
MM0 net16 A2 VSS VPW N12LL W=180.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=270.0n L=60.00n
MM4 Z net16 VDD VNW P12LL W=1.08u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=270.0n L=60.00n
.ENDS OR2HSV4RQ
****Sub-Circuit for OR2HSV8, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR2HSV8 A1 A2 Z VDD VSS
MM0 net31 A2 VSS VPW N12LL W=690.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=1.72u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=690.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=1.04u L=60.00n
MM4 Z net31 VDD VNW P12LL W=2.6u L=60.00n
MMP1 net42 A2 VDD VNW P12LL W=1.04u L=60.00n
.ENDS OR2HSV8
****Sub-Circuit for OR2HSV8RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV8RD A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=750.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=1.72u L=60.00n
MM0 net16 A2 VSS VPW N12LL W=750.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=1.3u L=60.00n
MM4 Z net16 VDD VNW P12LL W=2.16u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=1.3u L=60.00n
.ENDS OR2HSV8RD
****Sub-Circuit for OR2HSV8RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR2HSV8RQ A1 A2 Z VDD VSS
MMN1 net16 A1 VSS VPW N12LL W=290.00n L=60.00n
MM2 Z net16 VSS VPW N12LL W=1.72u L=60.00n
MM0 net16 A2 VSS VPW N12LL W=290.00n L=60.00n
MMP1 net15 A2 VDD VNW P12LL W=540.0n L=60.00n
MM4 Z net16 VDD VNW P12LL W=2.16u L=60.00n
MM1 net16 A1 net15 VNW P12LL W=540.0n L=60.00n
.ENDS OR2HSV8RQ
****Sub-Circuit for OR3HSV0, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR3HSV0 A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=200.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=300.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=300.00n L=60.00n
MM5 net054 A3 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=300.00n L=60.00n
.ENDS OR3HSV0
****Sub-Circuit for OR3HSV0RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR3HSV0RD A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=180.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=180.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=275.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=250.00n L=60.00n
MM5 net054 A3 VDD VNW P12LL W=275.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=275.00n L=60.00n
.ENDS OR3HSV0RD
****Sub-Circuit for OR3HSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR3HSV1 A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=200.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=300.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=440.00n L=60.00n
MM5 net054 A3 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=300.00n L=60.00n
.ENDS OR3HSV1
****Sub-Circuit for OR3HSV12, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR3HSV12 A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=550.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=550.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=2.58u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=550.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=1.3u L=60.00n
MM4 Z net31 VDD VNW P12LL W=3.24u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=1.3u L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=1.3u L=60.00n
.ENDS OR3HSV12
****Sub-Circuit for OR3HSV12RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR3HSV12RD A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=880.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=880.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=2.58u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=880.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=2.1u L=60.00n
MM4 Z net31 VDD VNW P12LL W=3.24u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=2.1u L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=2.1u L=60.00n
.ENDS OR3HSV12RD
****Sub-Circuit for OR3HSV12RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR3HSV12RQ A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=360.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=360.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=2.58u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=360.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=810n L=60.00n
MM4 Z net31 VDD VNW P12LL W=3.24u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=810n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=810n L=60.00n
.ENDS OR3HSV12RQ
****Sub-Circuit for OR3HSV16, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR3HSV16 A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=740.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=740.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=3.44u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=740.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=1.76u L=60.00n
MM4 Z net31 VDD VNW P12LL W=4.32u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=1.76u L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=1.76u L=60.00n
.ENDS OR3HSV16
****Sub-Circuit for OR3HSV16RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR3HSV16RD A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=1.175u L=60.00n
MM0 net31 A2 VSS VPW N12LL W=1.175u L=60.00n
MM2 Z net31 VSS VPW N12LL W=3.44u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=1.175u L=60.00n
MM1 net31 A1 net42 VNW P12LL W=2.8u L=60.00n
MM4 Z net31 VDD VNW P12LL W=4.32u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=2.8u L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=2.8u L=60.00n
.ENDS OR3HSV16RD
****Sub-Circuit for OR3HSV16RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR3HSV16RQ A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=450.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=450.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=3.44u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=450.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=1.08u L=60.00n
MM4 Z net31 VDD VNW P12LL W=4.32u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=1.08u L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=1.08u L=60.00n
.ENDS OR3HSV16RQ
****Sub-Circuit for OR3HSV1RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR3HSV1RD A1 A2 A3 Z VDD VSS
MM3 net050 A3 VSS VPW N12LL W=180.00n L=60.00n
MM0 net050 A2 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net050 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net050 A1 VSS VPW N12LL W=180.00n L=60.00n
MM1 net050 A1 net42 VNW P12LL W=355.00n L=60.00n
MM4 Z net050 VDD VNW P12LL W=440.00n L=60.00n
MM5 net054 A3 VDD VNW P12LL W=355.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=355.00n L=60.00n
.ENDS OR3HSV1RD
****Sub-Circuit for OR3HSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR3HSV2 A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=200.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=200.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=300.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=650.00n L=60.00n
MM5 net054 A3 VDD VNW P12LL W=300.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=300.00n L=60.00n
.ENDS OR3HSV2
****Sub-Circuit for OR3HSV2RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR3HSV2RD A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=180.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=180.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=360.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=540.00n L=60.00n
MM5 net054 A3 VDD VNW P12LL W=360.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=360.00n L=60.00n
.ENDS OR3HSV2RD
****Sub-Circuit for OR3HSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR3HSV4 A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=350.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=350.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=860.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=350.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=520.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=1.3u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=520.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=520.00n L=60.00n
.ENDS OR3HSV4
****Sub-Circuit for OR3HSV4RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR3HSV4RD A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=290.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=290.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=860.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=290.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=650.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=1.08u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=650.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=650.00n L=60.00n
.ENDS OR3HSV4RD
****Sub-Circuit for OR3HSV4RQ, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR3HSV4RQ A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=180.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=860.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=180.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=270.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=1.08u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=270.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=270.00n L=60.00n
.ENDS OR3HSV4RQ
****Sub-Circuit for OR3HSV8, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR3HSV8 A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=690.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=690.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=1.72u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=690.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=1.04u L=60.00n
MM4 Z net31 VDD VNW P12LL W=2.6u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=1.04u L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=1.04u L=60.00n
.ENDS OR3HSV8
****Sub-Circuit for OR3HSV8RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR3HSV8RD A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=590.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=590.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=1.72u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=590.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=1.3u L=60.00n
MM4 Z net31 VDD VNW P12LL W=2.16u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=1.3u L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=1.3u L=60.00n
.ENDS OR3HSV8RD
****Sub-Circuit for OR3HSV8RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR3HSV8RQ A1 A2 A3 Z VDD VSS
MM3 net31 A3 VSS VPW N12LL W=230.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=230.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=1.72u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=230.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=540.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=2.16u L=60.00n
MM5 net054 A3 VDD VNW P12LL W=540.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=540.00n L=60.00n
.ENDS OR3HSV8RQ
****Sub-Circuit for OR4HSV0, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR4HSV0 A1 A2 A3 A4 Z VDD VSS
MM6 net31 A4 VSS VPW N12LL W=200.00n L=60.00n
MM3 net31 A3 VSS VPW N12LL W=200.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=200.00n L=60.00n
MM7 net067 A4 VDD VNW P12LL W=300.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=300.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=300.00n L=60.00n
MM5 net054 A3 net067 VNW P12LL W=300.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=300.00n L=60.00n
.ENDS OR4HSV0
****Sub-Circuit for OR4HSV0RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR4HSV0RD A1 A2 A3 A4 Z VDD VSS
MM6 net31 A4 VSS VPW N12LL W=180.00n L=60.00n
MM3 net31 A3 VSS VPW N12LL W=180.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=200.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=180.00n L=60.00n
MM7 net067 A4 VDD VNW P12LL W=350.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=350.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=250.00n L=60.00n
MM5 net054 A3 net067 VNW P12LL W=350.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=350.00n L=60.00n
.ENDS OR4HSV0RD
****Sub-Circuit for OR4HSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR4HSV1 A1 A2 A3 A4 Z VDD VSS
MM6 net31 A4 VSS VPW N12LL W=200.00n L=60.00n
MM3 net31 A3 VSS VPW N12LL W=200.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=200.00n L=60.00n
MM7 net067 A4 VDD VNW P12LL W=300.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=300.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=440.00n L=60.00n
MM5 net054 A3 net067 VNW P12LL W=300.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=300.00n L=60.00n
.ENDS OR4HSV1
****Sub-Circuit for OR4HSV12RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR4HSV12RQ A1 A2 A3 A4 Z VDD VSS
MM7 net37 net49 VSS VPW N12LL W=3.77u L=60.00n
MM1 net53 A1 VSS VPW N12LL W=280.00n L=60.00n
MM8 net49 A4 VSS VPW N12LL W=280.00n L=60.00n
MM9 net49 A3 VSS VPW N12LL W=280.00n L=60.00n
MM2 net53 A2 VSS VPW N12LL W=280.00n L=60.00n
MM6 Z net53 net37 VPW N12LL W=3.77u L=60.00n
MM3 net80 A2 VDD VNW P12LL W=810n L=60.00n
MM11 net76 A4 VDD VNW P12LL W=810n L=60.00n
MM10 net49 A3 net76 VNW P12LL W=810n L=60.00n
MM5 Z net49 VDD VNW P12LL W=3.24u L=60.00n
MM4 Z net53 VDD VNW P12LL W=3.24u L=60.00n
MM0 net53 A1 net80 VNW P12LL W=810n L=60.00n
.ENDS OR4HSV12RQ
****Sub-Circuit for OR4HSV16RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR4HSV16RQ A1 A2 A3 A4 Z VDD VSS
MM11 net48 A4 VDD VNW P12LL W=1.08u L=60.00n
MM10 net69 A3 net48 VNW P12LL W=1.08u L=60.00n
MM0 net65 A1 net44 VNW P12LL W=1.08u L=60.00n
MM3 net44 A2 VDD VNW P12LL W=1.08u L=60.00n
MM5 Z net69 VDD VNW P12LL W=4.32u L=60.00n
MM4 Z net65 VDD VNW P12LL W=4.32u L=60.00n
MM8 net69 A4 VSS VPW N12LL W=375.00n L=60.00n
MM7 net81 net69 VSS VPW N12LL W=5.02u L=60.00n
MM1 net65 A1 VSS VPW N12LL W=375.00n L=60.00n
MM9 net69 A3 VSS VPW N12LL W=375.00n L=60.00n
MM2 net65 A2 VSS VPW N12LL W=375.00n L=60.00n
MM6 Z net65 net81 VPW N12LL W=5.02u L=60.00n
.ENDS OR4HSV16RQ
****Sub-Circuit for OR4HSV1RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR4HSV1RD A1 A2 A3 A4 Z VDD VSS
MM6 net31 A4 VSS VPW N12LL W=180.00n L=60.00n
MM3 net31 A3 VSS VPW N12LL W=180.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=350.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=180.00n L=60.00n
MM7 net067 A4 VDD VNW P12LL W=350.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=350.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=440.00n L=60.00n
MM5 net054 A3 net067 VNW P12LL W=350.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=350.00n L=60.00n
.ENDS OR4HSV1RD
****Sub-Circuit for OR4HSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR4HSV2 A1 A2 A3 A4 Z VDD VSS
MM6 net31 A4 VSS VPW N12LL W=200.00n L=60.00n
MM3 net31 A3 VSS VPW N12LL W=200.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=200.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=200.00n L=60.00n
MM7 net067 A4 VDD VNW P12LL W=300.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=300.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=650.00n L=60.00n
MM5 net054 A3 net067 VNW P12LL W=300.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=300.00n L=60.00n
.ENDS OR4HSV2
****Sub-Circuit for OR4HSV2RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR4HSV2RD A1 A2 A3 A4 Z VDD VSS
MM6 net31 A4 VSS VPW N12LL W=180.00n L=60.00n
MM3 net31 A3 VSS VPW N12LL W=180.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=430.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=180.00n L=60.00n
MM7 net067 A4 VDD VNW P12LL W=350.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=350.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=540.00n L=60.00n
MM5 net054 A3 net067 VNW P12LL W=350.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=350.00n L=60.00n
.ENDS OR4HSV2RD
****Sub-Circuit for OR4HSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR4HSV4 A1 A2 A3 A4 Z VDD VSS
MM6 net31 A4 VSS VPW N12LL W=350.00n L=60.00n
MM3 net31 A3 VSS VPW N12LL W=350.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=350.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=860.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=350.00n L=60.00n
MM7 net067 A4 VDD VNW P12LL W=520.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=520.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=1.3u L=60.00n
MM5 net054 A3 net067 VNW P12LL W=520.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=520.00n L=60.00n
.ENDS OR4HSV4
****Sub-Circuit for OR4HSV4RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR4HSV4RD A1 A2 A3 A4 Z VDD VSS
MM11 net48 A4 VDD VNW P12LL W=700n L=60.00n
MM10 net69 A3 net48 VNW P12LL W=700n L=60.00n
MM0 net65 A1 net44 VNW P12LL W=700n L=60.00n
MM3 net44 A2 VDD VNW P12LL W=700n L=60.00n
MM5 Z net69 VDD VNW P12LL W=1.08u L=60.00n
MM4 Z net65 VDD VNW P12LL W=1.08u L=60.00n
MM8 net69 A4 VSS VPW N12LL W=245.00n L=60.00n
MM7 net81 net69 VSS VPW N12LL W=1.26u L=60.00n
MM1 net65 A1 VSS VPW N12LL W=245.00n L=60.00n
MM9 net69 A3 VSS VPW N12LL W=245.00n L=60.00n
MM2 net65 A2 VSS VPW N12LL W=245.00n L=60.00n
MM6 Z net65 net81 VPW N12LL W=1.26u L=60.00n
.ENDS OR4HSV4RD
****Sub-Circuit for OR4HSV4RQ, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR4HSV4RQ A1 A2 A3 A4 Z VDD VSS
MM6 net31 A4 VSS VPW N12LL W=180.00n L=60.00n
MM3 net31 A3 VSS VPW N12LL W=180.00n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=180.00n L=60.00n
MM2 Z net31 VSS VPW N12LL W=860.00n L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=180.00n L=60.00n
MM7 net067 A4 VDD VNW P12LL W=270.00n L=60.00n
MM1 net31 A1 net42 VNW P12LL W=270.00n L=60.00n
MM4 Z net31 VDD VNW P12LL W=1.08u L=60.00n
MM5 net054 A3 net067 VNW P12LL W=270.00n L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=270.00n L=60.00n
.ENDS OR4HSV4RQ
****Sub-Circuit for OR4HSV8, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT OR4HSV8 A1 A2 A3 A4 Z VDD VSS
MM6 net31 A4 VSS VPW N12LL W=690.0n L=60.00n
MM3 net31 A3 VSS VPW N12LL W=690.0n L=60.00n
MM0 net31 A2 VSS VPW N12LL W=690.0n L=60.00n
MM2 Z net31 VSS VPW N12LL W=1.72u L=60.00n
MMN1 net31 A1 VSS VPW N12LL W=690.0n L=60.00n
MM7 net067 A4 VDD VNW P12LL W=1.04u L=60.00n
MM1 net31 A1 net42 VNW P12LL W=1.04u L=60.00n
MM4 Z net31 VDD VNW P12LL W=2.6u L=60.00n
MM5 net054 A3 net067 VNW P12LL W=1.04u L=60.00n
MMP1 net42 A2 net054 VNW P12LL W=1.04u L=60.00n
.ENDS OR4HSV8
****Sub-Circuit for OR4HSV8RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR4HSV8RD A1 A2 A3 A4 Z VDD VSS
MM8 net49 A4 VSS VPW N12LL W=490.00n L=60.00n
MM9 net49 A3 VSS VPW N12LL W=490.00n L=60.00n
MM6 Z net53 net37 VPW N12LL W=2.51u L=60.00n
MM1 net53 A1 VSS VPW N12LL W=490.00n L=60.00n
MM7 net37 net49 VSS VPW N12LL W=2.51u L=60.00n
MM2 net53 A2 VSS VPW N12LL W=490.00n L=60.00n
MM0 net53 A1 net80 VNW P12LL W=1.4u L=60.00n
MM11 net76 A4 VDD VNW P12LL W=1.4u L=60.00n
MM10 net49 A3 net76 VNW P12LL W=1.4u L=60.00n
MM4 Z net53 VDD VNW P12LL W=2.16u L=60.00n
MM5 Z net49 VDD VNW P12LL W=2.16u L=60.00n
MM3 net80 A2 VDD VNW P12LL W=1.4u L=60.00n
.ENDS OR4HSV8RD
****Sub-Circuit for OR4HSV8RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR4HSV8RQ A1 A2 A3 A4 Z VDD VSS
MM11 net48 A4 VDD VNW P12LL W=540n L=60.00n
MM10 net69 A3 net48 VNW P12LL W=540n L=60.00n
MM0 net65 A1 net44 VNW P12LL W=540n L=60.00n
MM3 net44 A2 VDD VNW P12LL W=540n L=60.00n
MM5 Z net69 VDD VNW P12LL W=2.16u L=60.00n
MM4 Z net65 VDD VNW P12LL W=2.16u L=60.00n
MM8 net69 A4 VSS VPW N12LL W=190.00n L=60.00n
MM7 net81 net69 VSS VPW N12LL W=2.51u L=60.00n
MM1 net65 A1 VSS VPW N12LL W=190.00n L=60.00n
MM9 net69 A3 VSS VPW N12LL W=190.00n L=60.00n
MM2 net65 A2 VSS VPW N12LL W=190.00n L=60.00n
MM6 Z net65 net81 VPW N12LL W=2.51u L=60.00n
.ENDS OR4HSV8RQ
****Sub-Circuit for OR5HSV0RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR5HSV0RD A1 A2 A3 A4 A5 Z VDD VSS
MM13 Z net43 VDD VNW P12LL W=250.00n L=60.00n
MM12 Z net55 VDD VNW P12LL W=250.00n L=60.00n
MM11 net26 A4 net18 VNW P12LL W=350.0n L=60.00n
MM10 net18 A5 VDD VNW P12LL W=350.0n L=60.00n
MM7 net43 A3 net26 VNW P12LL W=350.0n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=200.0n L=60.00n
MM1 net55 A1 net34 VNW P12LL W=200.0n L=60.00n
MM15 net35 net43 VSS VPW N12LL W=290.00n L=60.00n
MM14 Z net55 net35 VPW N12LL W=290.00n L=60.00n
MM6 net43 A3 VSS VPW N12LL W=180.00n L=60.00n
MM5 net43 A4 VSS VPW N12LL W=180.00n L=60.00n
MM3 net43 A5 VSS VPW N12LL W=180.00n L=60.00n
MMN1 net55 A1 VSS VPW N12LL W=180.00n L=60.00n
MM0 net55 A2 VSS VPW N12LL W=180.00n L=60.00n
.ENDS OR5HSV0RD
****Sub-Circuit for OR5HSV12RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR5HSV12RQ A1 A2 A3 A4 A5 Z VDD VSS
MM13 Z net43 VDD VNW P12LL W=3.24u L=60.00n
MM12 Z net55 VDD VNW P12LL W=3.24u L=60.00n
MM11 net26 A4 net18 VNW P12LL W=810.0n L=60.00n
MM10 net18 A5 VDD VNW P12LL W=810.0n L=60.00n
MM7 net43 A3 net26 VNW P12LL W=810.0n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=810.0n L=60.00n
MM1 net55 A1 net34 VNW P12LL W=810.0n L=60.00n
MM15 net35 net43 VSS VPW N12LL W=3.77u L=60.00n
MM14 Z net55 net35 VPW N12LL W=3.77u L=60.00n
MM6 net43 A3 VSS VPW N12LL W=340.00n L=60.00n
MM5 net43 A4 VSS VPW N12LL W=340.00n L=60.00n
MM3 net43 A5 VSS VPW N12LL W=340.00n L=60.00n
MMN1 net55 A1 VSS VPW N12LL W=440.00n L=60.00n
MM0 net55 A2 VSS VPW N12LL W=440.00n L=60.00n
.ENDS OR5HSV12RQ
****Sub-Circuit for OR5HSV16RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR5HSV16RQ A1 A2 A3 A4 A5 Z VDD VSS
MM13 Z net43 VDD VNW P12LL W=4.16u L=60.00n
MM12 Z net55 VDD VNW P12LL W=4.16u L=60.00n
MM11 net26 A4 net18 VNW P12LL W=1.08u L=60.00n
MM10 net18 A5 VDD VNW P12LL W=1.08u L=60.00n
MM7 net43 A3 net26 VNW P12LL W=1.08u L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=1.08u L=60.00n
MM1 net55 A1 net34 VNW P12LL W=1.08u L=60.00n
MM15 net35 net43 VSS VPW N12LL W=5.02u L=60.00n
MM14 Z net55 net35 VPW N12LL W=5.02u L=60.00n
MM6 net43 A3 VSS VPW N12LL W=450.00n L=60.00n
MM5 net43 A4 VSS VPW N12LL W=450.00n L=60.00n
MM3 net43 A5 VSS VPW N12LL W=450.00n L=60.00n
MMN1 net55 A1 VSS VPW N12LL W=580.00n L=60.00n
MM0 net55 A2 VSS VPW N12LL W=580.00n L=60.00n
.ENDS OR5HSV16RQ
****Sub-Circuit for OR5HSV1RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR5HSV1RD A1 A2 A3 A4 A5 Z VDD VSS
MM13 Z net43 VDD VNW P12LL W=440.00n L=60.00n
MM12 Z net55 VDD VNW P12LL W=440.00n L=60.00n
MM11 net26 A4 net18 VNW P12LL W=350.0n L=60.00n
MM10 net18 A5 VDD VNW P12LL W=350.0n L=60.00n
MM7 net43 A3 net26 VNW P12LL W=350.0n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=280.0n L=60.00n
MM1 net55 A1 net34 VNW P12LL W=280.0n L=60.00n
MM15 net35 net43 VSS VPW N12LL W=510.00n L=60.00n
MM14 Z net55 net35 VPW N12LL W=510.00n L=60.00n
MM6 net43 A3 VSS VPW N12LL W=180.00n L=60.00n
MM5 net43 A4 VSS VPW N12LL W=180.00n L=60.00n
MM3 net43 A5 VSS VPW N12LL W=180.00n L=60.00n
MMN1 net55 A1 VSS VPW N12LL W=180.00n L=60.00n
MM0 net55 A2 VSS VPW N12LL W=180.00n L=60.00n
.ENDS OR5HSV1RD
****Sub-Circuit for OR5HSV2RD, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR5HSV2RD A1 A2 A3 A4 A5 Z VDD VSS
MM13 Z net43 VDD VNW P12LL W=540.00n L=60.00n
MM12 Z net55 VDD VNW P12LL W=540.00n L=60.00n
MM11 net26 A4 net18 VNW P12LL W=350.0n L=60.00n
MM10 net18 A5 VDD VNW P12LL W=350.0n L=60.00n
MM7 net43 A3 net26 VNW P12LL W=350.0n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=350.0n L=60.00n
MM1 net55 A1 net34 VNW P12LL W=350.0n L=60.00n
MM15 net35 net43 VSS VPW N12LL W=630.00n L=60.00n
MM14 Z net55 net35 VPW N12LL W=630.00n L=60.00n
MM6 net43 A3 VSS VPW N12LL W=180.00n L=60.00n
MM5 net43 A4 VSS VPW N12LL W=180.00n L=60.00n
MM3 net43 A5 VSS VPW N12LL W=180.00n L=60.00n
MMN1 net55 A1 VSS VPW N12LL W=190.00n L=60.00n
MM0 net55 A2 VSS VPW N12LL W=190.00n L=60.00n
.ENDS OR5HSV2RD
****Sub-Circuit for OR5HSV4RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR5HSV4RD A1 A2 A3 A4 A5 Z VDD VSS
MM13 Z net43 VDD VNW P12LL W=1.08u L=60.00n
MM12 Z net55 VDD VNW P12LL W=1.08u L=60.00n
MM11 net26 A4 net18 VNW P12LL W=650.0n L=60.00n
MM10 net18 A5 VDD VNW P12LL W=650.0n L=60.00n
MM7 net43 A3 net26 VNW P12LL W=650.0n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=650.0n L=60.00n
MM1 net55 A1 net34 VNW P12LL W=650.0n L=60.00n
MM15 net35 net43 VSS VPW N12LL W=1.25u L=60.00n
MM14 Z net55 net35 VPW N12LL W=1.25u L=60.00n
MM6 net43 A3 VSS VPW N12LL W=290.00n L=60.00n
MM5 net43 A4 VSS VPW N12LL W=290.00n L=60.00n
MM3 net43 A5 VSS VPW N12LL W=290.00n L=60.00n
MMN1 net55 A1 VSS VPW N12LL W=380.00n L=60.00n
MM0 net55 A2 VSS VPW N12LL W=380.00n L=60.00n
.ENDS OR5HSV4RD
****Sub-Circuit for OR5HSV4RQ, Thu May 19 13:57:40 CST 2011****
.SUBCKT OR5HSV4RQ A1 A2 A3 A4 A5 Z VDD VSS
MM13 Z net43 VDD VNW P12LL W=1.08u L=60.00n
MM12 Z net55 VDD VNW P12LL W=1.08u L=60.00n
MM11 net26 A4 net18 VNW P12LL W=270.0n L=60.00n
MM10 net18 A5 VDD VNW P12LL W=270.0n L=60.00n
MM7 net43 A3 net26 VNW P12LL W=270.0n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=270.0n L=60.00n
MM1 net55 A1 net34 VNW P12LL W=270.0n L=60.00n
MM15 net35 net43 VSS VPW N12LL W=1.25u L=60.00n
MM14 Z net55 net35 VPW N12LL W=1.25u L=60.00n
MM6 net43 A3 VSS VPW N12LL W=180.00n L=60.00n
MM5 net43 A4 VSS VPW N12LL W=180.00n L=60.00n
MM3 net43 A5 VSS VPW N12LL W=180.00n L=60.00n
MMN1 net55 A1 VSS VPW N12LL W=180.00n L=60.00n
MM0 net55 A2 VSS VPW N12LL W=180.00n L=60.00n
.ENDS OR5HSV4RQ
****Sub-Circuit for OR5HSV8RD, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR5HSV8RD A1 A2 A3 A4 A5 Z VDD VSS
MM13 Z net43 VDD VNW P12LL W=2.16u L=60.00n
MM12 Z net55 VDD VNW P12LL W=2.16u L=60.00n
MM11 net26 A4 net18 VNW P12LL W=1.3u L=60.00n
MM10 net18 A5 VDD VNW P12LL W=1.3u L=60.00n
MM7 net43 A3 net26 VNW P12LL W=1.3u L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=1.3u L=60.00n
MM1 net55 A1 net34 VNW P12LL W=1.3u L=60.00n
MM15 net35 net43 VSS VPW N12LL W=2.51u L=60.00n
MM14 Z net55 net35 VPW N12LL W=2.51u L=60.00n
MM6 net43 A3 VSS VPW N12LL W=590.00n L=60.00n
MM5 net43 A4 VSS VPW N12LL W=590.00n L=60.00n
MM3 net43 A5 VSS VPW N12LL W=590.00n L=60.00n
MMN1 net55 A1 VSS VPW N12LL W=750.00n L=60.00n
MM0 net55 A2 VSS VPW N12LL W=750.00n L=60.00n
.ENDS OR5HSV8RD
****Sub-Circuit for OR5HSV8RQ, Thu Dec 23 11:14:06 CST 2010****
.SUBCKT OR5HSV8RQ A1 A2 A3 A4 A5 Z VDD VSS
MM13 Z net43 VDD VNW P12LL W=2.16u L=60.00n
MM12 Z net55 VDD VNW P12LL W=2.16u L=60.00n
MM11 net26 A4 net18 VNW P12LL W=540.0n L=60.00n
MM10 net18 A5 VDD VNW P12LL W=540.0n L=60.00n
MM7 net43 A3 net26 VNW P12LL W=540.0n L=60.00n
MMP1 net34 A2 VDD VNW P12LL W=540.0n L=60.00n
MM1 net55 A1 net34 VNW P12LL W=540.0n L=60.00n
MM15 net35 net43 VSS VPW N12LL W=2.51u L=60.00n
MM14 Z net55 net35 VPW N12LL W=2.51u L=60.00n
MM6 net43 A3 VSS VPW N12LL W=230.00n L=60.00n
MM5 net43 A4 VSS VPW N12LL W=230.00n L=60.00n
MM3 net43 A5 VSS VPW N12LL W=230.00n L=60.00n
MMN1 net55 A1 VSS VPW N12LL W=290.00n L=60.00n
MM0 net55 A2 VSS VPW N12LL W=290.00n L=60.00n
.ENDS OR5HSV8RQ
****Sub-Circuit for PULLHS0, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT PULLHS0 Z VDD VSS
MMN1 Z net18 VSS VPW N12LL W=300.00n L=60.00n
MMP1 net18 net18 VDD VNW P12LL W=300.00n L=60.00n
.ENDS PULLHS0
****Sub-Circuit for PULLHS1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT PULLHS1 Z VDD VSS
MMN1 net14 net14 VSS VPW N12LL W=200.00n L=60.00n
MMP1 Z net14 VDD VNW P12LL W=450.00n L=60.00n
.ENDS PULLHS1
****Sub-Circuit for SDGRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNHSV1 CK D Q QN RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM52 QN ps VSS VPW N12LL W=290.00n L=60.00n
MM3 m c ps VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=410.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=270.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=410.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM53 QN ps VDD VNW P12LL W=440.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=530.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=410.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=530.00n L=60.00n
MM1 m pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS SDGRNHSV1
****Sub-Circuit for SDGRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNHSV2 CK D Q QN RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM52 QN ps VSS VPW N12LL W=430.00n L=60.00n
MM3 m c ps VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=340.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=340.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=410.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=340.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=270.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=410.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM53 QN ps VDD VNW P12LL W=650.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=530.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=410.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=530.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRNHSV2
****Sub-Circuit for SDGRNHSV4, Fri Dec 10 10:21:28 CST 2010****
.SUBCKT SDGRNHSV4 CK D Q QN RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM52 QN ps VSS VPW N12LL W=860.00n L=60.00n
MM3 m c ps VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=360.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=410.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=270.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=410.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=410.00n L=60.00n
MM0 m pm VSS VPW N12LL W=390.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM53 QN ps VDD VNW P12LL W=1.3u L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=540.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=530.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=410.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=530.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRNHSV4
****Sub-Circuit for SDGRNQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNQHSV1 CK D Q RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM3 m c ps VPW N12LL W=350.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=380.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=260.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=250.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=380.00n L=60.00n
MM0 m pm VSS VPW N12LL W=350.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=530.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=500.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=390.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=380.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=530.00n L=60.00n
.ENDS SDGRNQHSV1
****Sub-Circuit for SDGRNQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRNQHSV2 CK D Q RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM3 m c ps VPW N12LL W=360.00n L=60.00n
MM30 c cn VSS VPW N12LL W=330.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=330.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=380.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=340.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=250.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=380.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=500.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=500.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=500.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=380.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRNQHSV2
****Sub-Circuit for SDGRNQHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SDGRNQHSV4 CK D Q RN SE SI VDD VSS
MM41 net_0127 SE net_0123 VPW N12LL W=300.00n L=60.00n
MM43 net_0123 SI VSS VPW N12LL W=300.00n L=60.00n
MM46 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM3 m c ps VPW N12LL W=370.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=360.00n L=60.00n
MM38 net_0162 RN VSS VPW N12LL W=380.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=300.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=300.00n L=60.00n
MM48 net_0127 cn pm VPW N12LL W=250.00n L=60.00n
MM40 net_0127 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D net_0162 VPW N12LL W=380.00n L=60.00n
MM0 m pm VSS VPW N12LL W=390.00n L=60.00n
MM44 net_0202 SI VDD VNW P12LL W=450.00n L=60.00n
MM45 net_0127 SEN net_0202 VNW P12LL W=450.00n L=60.00n
MM47 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM50 net_0178 SE VDD VNW P12LL W=300.0n L=60.00n
MM51 net_0127 RN net_0178 VNW P12LL W=300.0n L=60.00n
MM4 m cn ps VNW P12LL W=540.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=540.00n L=60.00n
MM37 net128 D VDD VNW P12LL W=500.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=450.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=450.00n L=60.00n
MM49 net_0127 c pm VNW P12LL W=360.00n L=60.00n
MM39 net_0127 SE net128 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=580.00n L=60.00n
.ENDS SDGRNQHSV4
****Sub-Circuit for SDGRSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRSNHSV1 CK D Q QN RN SE SI SN VDD VSS
MM45 net0370 SE net201 VPW N12LL W=300.00n L=60.00n
MM46 net201 SI VSS VPW N12LL W=300.00n L=60.00n
MM47 net0172 RN VSS VPW N12LL W=390.00n L=60.00n
MM48 net0370 SEN net213 VPW N12LL W=340.00n L=60.00n
MM49 net213 D net205 VPW N12LL W=390.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=300.00n L=60.00n
MM39 QN OS VSS VPW N12LL W=290.00n L=60.00n
MM62 OS c net181 VPW N12LL W=260.00n L=60.00n
MM63 net181 S VSS VPW N12LL W=260.00n L=60.00n
MM61 M cn net193 VPW N12LL W=300.00n L=60.00n
MM58 SEN SE VSS VPW N12LL W=300.00n L=60.00n
MM70 net205 SN net0172 VPW N12LL W=390.00n L=60.00n
MM60 net193 net0370 VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=230.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=230.00n L=60.00n
MM24 net172 cn OS VPW N12LL W=200.00n L=60.00n
MM23 VSS NET64 net172 VPW N12LL W=200.00n L=60.00n
MM69 net213 SNN net0172 VPW N12LL W=300.00n L=60.00n
MM19 Q NET64 VSS VPW N12LL W=290.00n L=60.00n
MM17 NET64 OS VSS VPW N12LL W=260.00n L=60.00n
MM12 net240 c M VPW N12LL W=200.00n L=60.00n
MM11 VSS S net240 VPW N12LL W=200.00n L=60.00n
MM0 S M VSS VPW N12LL W=300.00n L=60.00n
MM66 net0418 SNN net296 VNW P12LL W=590.00n L=60.00n
MM50 net288 SI VDD VNW P12LL W=420.00n L=60.00n
MM51 net0370 SEN net288 VNW P12LL W=420.00n L=60.00n
MM52 net296 D VDD VNW P12LL W=590.00n L=60.00n
MM53 net0370 SE net0418 VNW P12LL W=590.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=450.00n L=60.00n
MM40 QN OS VDD VNW P12LL W=440.00n L=60.00n
MM64 net268 S VDD VNW P12LL W=390.00n L=60.00n
MM65 OS cn net268 VNW P12LL W=390.00n L=60.00n
MM67 net0418 RN VDD VNW P12LL W=450.00n L=60.00n
MM59 SEN SE VDD VNW P12LL W=450.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=360.00n L=60.00n
MM26 VDD NET64 net253 VNW P12LL W=300.00n L=60.00n
MM25 net253 c OS VNW P12LL W=300.00n L=60.00n
MM20 Q NET64 VDD VNW P12LL W=440.00n L=60.00n
MM18 NET64 OS VDD VNW P12LL W=390.00n L=60.00n
MM14 net313 cn M VNW P12LL W=300.00n L=60.00n
MM13 VDD S net313 VNW P12LL W=300.00n L=60.00n
MM55 net280 net0370 VDD VNW P12LL W=450.00n L=60.00n
MM56 M c net280 VNW P12LL W=450.00n L=60.00n
MM1 S M VDD VNW P12LL W=450.00n L=60.00n
.ENDS SDGRSNHSV1
****Sub-Circuit for SDGRSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRSNHSV2 CK D Q QN RN SE SI SN VDD VSS
MM45 net0370 SE net201 VPW N12LL W=270.00n L=60.00n
MM46 net201 SI VSS VPW N12LL W=270.00n L=60.00n
MM47 net0172 RN VSS VPW N12LL W=350.00n L=60.00n
MM48 net0370 SEN net213 VPW N12LL W=350.00n L=60.00n
MM49 net213 D net205 VPW N12LL W=350.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=290.00n L=60.00n
MM39 QN OS VSS VPW N12LL W=430.00n L=60.00n
MM62 OS c net181 VPW N12LL W=400.00n L=60.00n
MM63 net181 S VSS VPW N12LL W=400.00n L=60.00n
MM61 M cn net193 VPW N12LL W=260.00n L=60.00n
MM58 SEN SE VSS VPW N12LL W=290.00n L=60.00n
MM70 net205 SN net0172 VPW N12LL W=350.00n L=60.00n
MM60 net193 net0370 VSS VPW N12LL W=260.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net172 cn OS VPW N12LL W=200.00n L=60.00n
MM23 VSS NET64 net172 VPW N12LL W=200.00n L=60.00n
MM69 net213 SNN net0172 VPW N12LL W=300.00n L=60.00n
MM19 Q NET64 VSS VPW N12LL W=430.00n L=60.00n
MM17 NET64 OS VSS VPW N12LL W=300.00n L=60.00n
MM12 net240 c M VPW N12LL W=200.00n L=60.00n
MM11 VSS S net240 VPW N12LL W=200.00n L=60.00n
MM0 S M VSS VPW N12LL W=360.00n L=60.00n
MM66 net0418 SNN net296 VNW P12LL W=590.00n L=60.00n
MM50 net288 SI VDD VNW P12LL W=410.00n L=60.00n
MM51 net0370 SEN net288 VNW P12LL W=410.00n L=60.00n
MM52 net296 D VDD VNW P12LL W=590.00n L=60.00n
MM53 net0370 SE net0418 VNW P12LL W=590.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=440.00n L=60.00n
MM40 QN OS VDD VNW P12LL W=650.00n L=60.00n
MM64 net268 S VDD VNW P12LL W=480.00n L=60.00n
MM65 OS cn net268 VNW P12LL W=480.00n L=60.00n
MM67 net0418 RN VDD VNW P12LL W=400.00n L=60.00n
MM59 SEN SE VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD NET64 net253 VNW P12LL W=300.00n L=60.00n
MM25 net253 c OS VNW P12LL W=300.00n L=60.00n
MM20 Q NET64 VDD VNW P12LL W=650.00n L=60.00n
MM18 NET64 OS VDD VNW P12LL W=450.00n L=60.00n
MM14 net313 cn M VNW P12LL W=300.00n L=60.00n
MM13 VDD S net313 VNW P12LL W=300.00n L=60.00n
MM55 net280 net0370 VDD VNW P12LL W=390.00n L=60.00n
MM56 M c net280 VNW P12LL W=390.00n L=60.00n
MM1 S M VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRSNHSV2
****Sub-Circuit for SDGRSNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGRSNHSV4 CK D Q QN RN SE SI SN VDD VSS
MM45 net0370 SE net201 VPW N12LL W=300.00n L=60.00n
MM46 net201 SI VSS VPW N12LL W=300.00n L=60.00n
MM47 net0172 RN VSS VPW N12LL W=350.00n L=60.00n
MM48 net0370 SEN net213 VPW N12LL W=350.00n L=60.00n
MM49 net213 D net205 VPW N12LL W=350.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=290.00n L=60.00n
MM39 QN OS VSS VPW N12LL W=860.00n L=60.00n
MM62 OS c net181 VPW N12LL W=450.00n L=60.00n
MM63 net181 S VSS VPW N12LL W=450.00n L=60.00n
MM61 M cn net193 VPW N12LL W=260.00n L=60.00n
MM58 SEN SE VSS VPW N12LL W=290.00n L=60.00n
MM70 net205 SN net0172 VPW N12LL W=350.00n L=60.00n
MM60 net193 net0370 VSS VPW N12LL W=260.00n L=60.00n
MM30 c cn VSS VPW N12LL W=260.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net172 cn OS VPW N12LL W=200.00n L=60.00n
MM23 VSS NET64 net172 VPW N12LL W=200.00n L=60.00n
MM69 net213 SNN net0172 VPW N12LL W=300.00n L=60.00n
MM19 Q NET64 VSS VPW N12LL W=860.00n L=60.00n
MM17 NET64 OS VSS VPW N12LL W=360.00n L=60.00n
MM12 net240 c M VPW N12LL W=200.00n L=60.00n
MM11 VSS S net240 VPW N12LL W=200.00n L=60.00n
MM0 S M VSS VPW N12LL W=360.00n L=60.00n
MM66 net0418 SNN net296 VNW P12LL W=590.00n L=60.00n
MM50 net288 SI VDD VNW P12LL W=450.00n L=60.00n
MM51 net0370 SEN net288 VNW P12LL W=450.00n L=60.00n
MM52 net296 D VDD VNW P12LL W=590.00n L=60.00n
MM53 net0370 SE net0418 VNW P12LL W=590.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=440.00n L=60.00n
MM40 QN OS VDD VNW P12LL W=1.3u L=60.00n
MM64 net268 S VDD VNW P12LL W=570.00n L=60.00n
MM65 OS cn net268 VNW P12LL W=570.00n L=60.00n
MM67 net0418 RN VDD VNW P12LL W=400.00n L=60.00n
MM59 SEN SE VDD VNW P12LL W=440.00n L=60.00n
MM29 c cn VDD VNW P12LL W=390.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD NET64 net253 VNW P12LL W=300.00n L=60.00n
MM25 net253 c OS VNW P12LL W=300.00n L=60.00n
MM20 Q NET64 VDD VNW P12LL W=1.3u L=60.00n
MM18 NET64 OS VDD VNW P12LL W=540.00n L=60.00n
MM14 net313 cn M VNW P12LL W=300.00n L=60.00n
MM13 VDD S net313 VNW P12LL W=300.00n L=60.00n
MM55 net280 net0370 VDD VNW P12LL W=390.00n L=60.00n
MM56 M c net280 VNW P12LL W=390.00n L=60.00n
MM1 S M VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDGRSNHSV4
****Sub-Circuit for SDGSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGSNHSV1 CK D Q QN SE SI SN VDD VSS
MM39 QN PS VSS VPW N12LL W=290.00n L=60.00n
MM45 N74 SE net0128 VPW N12LL W=200.00n L=60.00n
MM46 net0128 SI VSS VPW N12LL W=200.00n L=60.00n
MM48 N74 cn PM VPW N12LL W=270.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=200.00n L=60.00n
MM52 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM3 M c PS VPW N12LL W=270.00n L=60.00n
MM42 net69 SNN VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=250.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn PS VPW N12LL W=200.00n L=60.00n
MM23 VSS S net48 VPW N12LL W=200.00n L=60.00n
MM19 Q S VSS VPW N12LL W=290.00n L=60.00n
MM17 S PS VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c PM VPW N12LL W=200.00n L=60.00n
MM11 VSS M net52 VPW N12LL W=200.00n L=60.00n
MM9 N74 SEN net69 VPW N12LL W=250.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=250.00n L=60.00n
MM0 M PM VSS VPW N12LL W=270.00n L=60.00n
MM41 net_0231 SNN VDD VNW P12LL W=400.00n L=60.00n
MM40 QN PS VDD VNW P12LL W=440.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=300.00n L=60.00n
MM50 net0207 SI VDD VNW P12LL W=300.00n L=60.00n
MM51 N74 SEN net0207 VNW P12LL W=300.00n L=60.00n
MM54 N74 c PM VNW P12LL W=400.00n L=60.00n
MM4 M cn PS VNW P12LL W=400.00n L=60.00n
MM29 c cn VDD VNW P12LL W=380.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD S net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c PS VNW P12LL W=300.00n L=60.00n
MM20 Q S VDD VNW P12LL W=440.00n L=60.00n
MM18 S PS VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn PM VNW P12LL W=300.00n L=60.00n
MM13 VDD M net117 VNW P12LL W=300.00n L=60.00n
MM10 N74 SE net128 VNW P12LL W=400.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=400.00n L=60.00n
MM56 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM1 M PM VDD VNW P12LL W=400.00n L=60.00n
.ENDS SDGSNHSV1
****Sub-Circuit for SDGSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGSNHSV2 CK D Q QN SE SI SN VDD VSS
MM39 QN PS VSS VPW N12LL W=430.00n L=60.00n
MM45 N74 SE net0128 VPW N12LL W=200.00n L=60.00n
MM46 net0128 SI VSS VPW N12LL W=200.00n L=60.00n
MM48 N74 cn PM VPW N12LL W=360.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=200.00n L=60.00n
MM52 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM3 M c PS VPW N12LL W=390.00n L=60.00n
MM42 net69 SNN VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=380.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn PS VPW N12LL W=200.00n L=60.00n
MM23 VSS S net48 VPW N12LL W=200.00n L=60.00n
MM19 Q S VSS VPW N12LL W=430.00n L=60.00n
MM17 S PS VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c PM VPW N12LL W=200.00n L=60.00n
MM11 VSS M net52 VPW N12LL W=200.00n L=60.00n
MM9 N74 SEN net69 VPW N12LL W=380.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=380.00n L=60.00n
MM0 M PM VSS VPW N12LL W=390.00n L=60.00n
MM41 net_0231 SNN VDD VNW P12LL W=600.0n L=60.00n
MM40 QN PS VDD VNW P12LL W=650.00n L=60.00n
MM44 SNN SN VDD VNW P12LL W=300.00n L=60.00n
MM50 net0207 SI VDD VNW P12LL W=300.00n L=60.00n
MM51 N74 SEN net0207 VNW P12LL W=300.00n L=60.00n
MM54 N74 c PM VNW P12LL W=540.00n L=60.00n
MM4 M cn PS VNW P12LL W=580.00n L=60.00n
MM29 c cn VDD VNW P12LL W=570.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD S net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c PS VNW P12LL W=300.00n L=60.00n
MM20 Q S VDD VNW P12LL W=650.00n L=60.00n
MM18 S PS VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn PM VNW P12LL W=300.00n L=60.00n
MM13 VDD M net117 VNW P12LL W=300.00n L=60.00n
MM10 N74 SE net128 VNW P12LL W=600.0n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=600.0n L=60.00n
MM56 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM1 M PM VDD VNW P12LL W=580.00n L=60.00n
.ENDS SDGSNHSV2
****Sub-Circuit for SDGSNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDGSNHSV4 CK D Q QN SE SI SN VDD VSS
MM39 QN PS VSS VPW N12LL W=860.00n L=60.00n
MM45 N74 SE net0128 VPW N12LL W=200.00n L=60.00n
MM46 net0128 SI VSS VPW N12LL W=200.00n L=60.00n
MM48 N74 cn PM VPW N12LL W=400.00n L=60.00n
MM43 SNN SN VSS VPW N12LL W=200.00n L=60.00n
MM52 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM3 M c PS VPW N12LL W=430.00n L=60.00n
MM42 net69 SNN VSS VPW N12LL W=250.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn PS VPW N12LL W=200.00n L=60.00n
MM23 VSS S net48 VPW N12LL W=200.00n L=60.00n
MM19 Q S VSS VPW N12LL W=860.00n L=60.00n
MM17 S PS VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c PM VPW N12LL W=200.00n L=60.00n
MM11 VSS M net52 VPW N12LL W=200.00n L=60.00n
MM9 N74 SEN net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D VSS VPW N12LL W=430.00n L=60.00n
MM0 M PM VSS VPW N12LL W=430.00n L=60.00n
MM41 net_0231 SNN VDD VNW P12LL W=650.00n L=60.00n
MM40 QN PS VDD VNW P12LL W=1.3u L=60.00n
MM44 SNN SN VDD VNW P12LL W=300.00n L=60.00n
MM50 net0207 SI VDD VNW P12LL W=300.00n L=60.00n
MM51 N74 SEN net0207 VNW P12LL W=300.00n L=60.00n
MM54 N74 c PM VNW P12LL W=600.0n L=60.00n
MM4 M cn PS VNW P12LL W=650.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD S net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c PS VNW P12LL W=300.00n L=60.00n
MM20 Q S VDD VNW P12LL W=1.3u L=60.00n
MM18 S PS VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn PM VNW P12LL W=300.00n L=60.00n
MM13 VDD M net117 VNW P12LL W=300.00n L=60.00n
MM10 N74 SE net128 VNW P12LL W=650.00n L=60.00n
MM8 net128 D net_0231 VNW P12LL W=650.00n L=60.00n
MM56 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM1 M PM VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDGSNHSV4
****Sub-Circuit for SDHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDHSV1 CK D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=290.00n L=60.00n
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=280.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=280.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=290.00n L=60.00n
MM53 QN s VDD VNW P12LL W=440.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=300.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=300.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDHSV1
****Sub-Circuit for SDHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDHSV2 CK D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=430.00n L=60.00n
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=400.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=400.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM53 QN s VDD VNW P12LL W=650.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDHSV2
****Sub-Circuit for SDHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDHSV4 CK D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=860.00n L=60.00n
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=420.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=300.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=300.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM53 QN s VDD VNW P12LL W=1.3u L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=520.0n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=520.0n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.0n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDHSV4
****Sub-Circuit for SDQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDQHSV1 CK D Q SE SI VDD VSS
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=280.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=280.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=290.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=300.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=300.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDQHSV1
****Sub-Circuit for SDQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDQHSV2 CK D Q SE SI VDD VSS
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=400.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=400.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=440.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=440.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDQHSV2
****Sub-Circuit for SDQHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SDQHSV4 CK D Q SE SI VDD VSS
MM46 net_0107 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0163 SE net_0107 VPW N12LL W=200.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=430.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=430.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=300.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=300.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=300.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=300.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=300.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM51 net128 SEN net_0174 VNW P12LL W=300.00n L=60.00n
MM50 net_0174 SI VDD VNW P12LL W=300.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=490.0n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=490.0n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.0n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=450.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=450.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=450.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SDQHSV4
****Sub-Circuit for SDRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNHSV1 CK D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=290.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=290.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=290.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=290.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=440.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=330.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=330.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=330.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDRNHSV1
****Sub-Circuit for SDRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNHSV2 CK D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=430.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=320.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=320.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=650.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=350.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=350.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=350.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNHSV2
****Sub-Circuit for SDRNHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SDRNHSV4 CK D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=430.00n L=60.00n m=2
MM45 net_0137 sen net_0133 VPW N12LL W=430.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=400.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=300.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=300.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=650.00n L=60.00n m=2
MM47 net_0137 SE net_0212 VNW P12LL W=500n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=450.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=500n L=60.00n
MM8 net128 SI VDD VNW P12LL W=500n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNHSV4
****Sub-Circuit for SDRNQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNQHSV1 CK D Q RDN SE SI VDD VSS
MM45 net_0137 sen net_0133 VPW N12LL W=290.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=290.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=290.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=290.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=290.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=290.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=290.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=290.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=290.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=330.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=330.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=300.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=330.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=330.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDRNQHSV1
****Sub-Circuit for SDRNQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNQHSV2 CK D Q RDN SE SI VDD VSS
MM45 net_0137 sen net_0133 VPW N12LL W=320.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=320.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=200.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=320.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=390.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=390.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200n L=60.00n
MM27 cn CK VSS VPW N12LL W=200n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=320.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=320.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=350.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=350.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=400.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=350.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=350.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNQHSV2
****Sub-Circuit for SDRNQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRNQHSV4 CK D Q RDN SE SI VDD VSS
MM45 net_0137 sen net_0133 VPW N12LL W=430.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=430.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=360.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=340.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=400.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=200n L=60.00n
MM39 s ps net_099 VPW N12LL W=300.00n L=60.00n m=2
MM40 net_099 RDN VSS VPW N12LL W=300.00n L=60.00n m=2
MM30 c cn VSS VPW N12LL W=430n L=60.00n
MM27 cn CK VSS VPW N12LL W=300n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=430.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=350.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=500n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM38 s ps VDD VNW P12LL W=450.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=530.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn ps VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=500n L=60.00n
MM8 net128 SI VDD VNW P12LL W=500n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=540.00n L=60.00n
.ENDS SDRNQHSV4
****Sub-Circuit for SDRSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRSNHSV1 CK D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=250.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=290.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=200.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=260.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=260.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=260.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=260.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=280.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=330.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=420.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=380.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=330.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=330.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=330.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=440.00n L=60.00n
.ENDS SDRSNHSV1
****Sub-Circuit for SDRSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDRSNHSV2 CK D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=280.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=250.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=360.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=390.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=200.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=220.00n L=60.00n
MM40 net43 R L VPW N12LL W=280.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=220.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=220.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=220.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=300.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=510.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=380.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=300.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=300.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=300.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=600.00n L=60.00n
.ENDS SDRSNHSV2
****Sub-Circuit for SDRSNHSV4, Mon May 30 16:10:14 CST 2011****
.SUBCKT SDRSNHSV4 CK D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=200.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=280.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=250.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=320.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n m=2
MM39 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=430.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=400.00n L=60.00n
MM40 net43 R L VPW N12LL W=280.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=400.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=400.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=400.00n L=60.00n
MM30 c cn VSS VPW N12LL W=430.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n m=2
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=500.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n m=2
MM57 net_0140 c net_0139 VNW P12LL W=580.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=600.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=520.00n L=60.00n
MM29 c cn VDD VNW P12LL W=620.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=450.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n m=2
MM4 net_0154 cn net43 VNW P12LL W=380.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=500.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=500.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=500.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=650.00n L=60.00n
.ENDS SDRSNHSV4
****Sub-Circuit for SDSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDSNHSV1 CK D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=300.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=300.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=200.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=290.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=400.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=200.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=400.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=300.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=450.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=450.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=400.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=400.00n L=60.00n
.ENDS SDSNHSV1
****Sub-Circuit for SDSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDSNHSV2 CK D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=300.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=300.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=200.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=420.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=420.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=300.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=450.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=450.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=500.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=650.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=390.00n L=60.00n
.ENDS SDSNHSV2
****Sub-Circuit for SDSNHSV4, Mon May 30 17:13:17 CST 2011****
.SUBCKT SDSNHSV4 CK D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=300.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=300.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=200.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=200.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=360.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=300.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=450.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=450.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=300.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM38 s net43 VDD VNW P12LL W=650.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=300.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=625.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=480.00n L=60.00n
.ENDS SDSNHSV4
****Sub-Circuit for SDXHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDXHSV1 CK DA DB Q QN SA SE SI VDD VSS
MM5 net41 SB net_0171 VPW N12LL W=240.00n L=60.00n
MM49 net39 DA VSS VPW N12LL W=350.00n L=60.00n
MM48 net39 SA net_0171 VPW N12LL W=240.00n L=60.00n
MM37 SEN SE VSS VPW N12LL W=240.00n L=60.00n
MM41 net41 DB VSS VPW N12LL W=350.00n L=60.00n
MM31 SB SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=350.00n L=60.00n
MM19 QN s VSS VPW N12LL W=350.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM7 m c net43 VPW N12LL W=350.00n L=60.00n
MM12 net52 c net_0157 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM46 net_0169 SE VSS VPW N12LL W=240.00n L=60.00n
MM45 net_0153 sin net_0169 VPW N12LL W=240.00n L=60.00n
MM43 net_0161 SEN VSS VPW N12LL W=300.00n L=60.00n
MM9 net_0157 cn net_0153 VPW N12LL W=300.00n L=60.00n
MM42 net_0153 net_0171 net_0161 VPW N12LL W=300.00n L=60.00n
MM6 sin SI VSS VPW N12LL W=350.00n L=60.00n
MM0 m net_0157 VSS VPW N12LL W=350.00n L=60.00n
MM52 net39 DA VDD VNW P12LL W=440.0n L=60.00n
MM53 sin SI VDD VNW P12LL W=440.0n L=60.00n
MM54 net41 SA net_0171 VNW P12LL W=300.0n L=60.00n
MM55 net41 DB VDD VNW P12LL W=440.0n L=60.00n
MM56 net39 SB net_0171 VNW P12LL W=300.0n L=60.00n
MM38 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM4 m cn net43 VNW P12LL W=440.0n L=60.00n
MM44 net_0236 SE VDD VNW P12LL W=450.00n L=60.00n
MM32 SB SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=440.00n L=60.00n
MM20 QN s VDD VNW P12LL W=440.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=300.00n L=60.00n
MM47 net_0233 net_0171 net_0236 VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0157 VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM51 net_0233 sin net_0252 VNW P12LL W=300.00n L=60.00n
MM50 net_0252 SEN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0157 c net_0233 VNW P12LL W=450.00n L=60.00n
MM1 m net_0157 VDD VNW P12LL W=440.00n L=60.00n
.ENDS SDXHSV1
****Sub-Circuit for SDXHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDXHSV2 CK DA DB Q QN SA SE SI VDD VSS
MM8 sin SI VSS VPW N12LL W=350.00n L=60.00n
MM41 net41 DB VSS VPW N12LL W=430.00n L=60.00n
MM37 SEN SE VSS VPW N12LL W=240.00n L=60.00n
MM31 SB SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=430.00n L=60.00n
MM19 QN s VSS VPW N12LL W=430.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=350.00n L=60.00n
MM2 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0157 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM46 net_0169 SE VSS VPW N12LL W=240.00n L=60.00n
MM45 net_0153 sin net_0169 VPW N12LL W=240.00n L=60.00n
MM43 net_0161 SEN VSS VPW N12LL W=350.00n L=60.00n
MM9 net_0157 cn net_0153 VPW N12LL W=350.00n L=60.00n
MM42 net_0153 net_0152 net_0161 VPW N12LL W=350.00n L=60.00n
MM48 net39 SA net_0152 VPW N12LL W=240.00n L=60.00n
MM5 net41 SB net_0152 VPW N12LL W=240.00n L=60.00n
MM49 net39 DA VSS VPW N12LL W=430.00n L=60.00n
MM0 m net_0157 VSS VPW N12LL W=430.00n L=60.00n
MM38 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM53 sin SI VDD VNW P12LL W=440.0n L=60.00n
MM44 net_0236 SE VDD VNW P12LL W=440.00n L=60.00n
MM32 SB SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=550.00n L=60.00n
MM20 QN s VDD VNW P12LL W=550.00n L=60.00n
MM18 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM7 m cn net43 VNW P12LL W=540.00n L=60.00n
MM47 net_0233 net_0152 net_0236 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0157 VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM51 net_0233 sin net_0252 VNW P12LL W=300.00n L=60.00n
MM50 net_0252 SEN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0157 c net_0233 VNW P12LL W=440.00n L=60.00n
MM56 net39 SB net_0152 VNW P12LL W=300.0n L=60.00n
MM54 net41 SA net_0152 VNW P12LL W=300.0n L=60.00n
MM55 net41 DB VDD VNW P12LL W=550.0n L=60.00n
MM52 net39 DA VDD VNW P12LL W=550.0n L=60.00n
MM1 m net_0157 VDD VNW P12LL W=550.00n L=60.00n
.ENDS SDXHSV2
****Sub-Circuit for SDXHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SDXHSV4 CK DA DB Q QN SA SE SI VDD VSS
MM8 sin SI VSS VPW N12LL W=350.00n L=60.00n
MM41 net41 DB VSS VPW N12LL W=430.00n L=60.00n
MM37 SEN SE VSS VPW N12LL W=240.00n L=60.00n
MM31 SB SA VSS VPW N12LL W=240.00n L=60.00n
MM30 c cn VSS VPW N12LL W=350.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=240.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q net43 VSS VPW N12LL W=860.00n L=60.00n
MM19 QN s VSS VPW N12LL W=860.00n L=60.00n
MM17 s net43 VSS VPW N12LL W=430.00n L=60.00n
MM2 m c net43 VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0157 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM46 net_0169 SE VSS VPW N12LL W=240.00n L=60.00n
MM45 net_0153 sin net_0169 VPW N12LL W=240.00n L=60.00n
MM43 net_0161 SEN VSS VPW N12LL W=350.00n L=60.00n
MM9 net_0157 cn net_0153 VPW N12LL W=350.00n L=60.00n
MM42 net_0153 net_0152 net_0161 VPW N12LL W=350.00n L=60.00n
MM49 net39 DA VSS VPW N12LL W=430.00n L=60.00n
MM5 net41 SB net_0152 VPW N12LL W=240.00n L=60.00n
MM48 net39 SA net_0152 VPW N12LL W=240.00n L=60.00n
MM0 m net_0157 VSS VPW N12LL W=430.00n L=60.00n
MM38 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM44 net_0236 SE VDD VNW P12LL W=440.00n L=60.00n
MM56 net39 SB net_0152 VNW P12LL W=300.0n L=60.00n
MM54 net41 SA net_0152 VNW P12LL W=300.0n L=60.00n
MM52 net39 DA VDD VNW P12LL W=550.0n L=60.00n
MM55 net41 DB VDD VNW P12LL W=550.0n L=60.00n
MM32 SB SA VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=200.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=200.00n L=60.00n
MM21 Q net43 VDD VNW P12LL W=1.1u L=60.00n
MM20 QN s VDD VNW P12LL W=1.1u L=60.00n
MM18 s net43 VDD VNW P12LL W=550.00n L=60.00n
MM53 sin SI VDD VNW P12LL W=440.0n L=60.00n
MM7 m cn net43 VNW P12LL W=540.00n L=60.00n
MM47 net_0233 net_0152 net_0236 VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0157 VNW P12LL W=200.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=200.00n L=60.00n
MM51 net_0233 sin net_0252 VNW P12LL W=300.00n L=60.00n
MM50 net_0252 SEN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0157 c net_0233 VNW P12LL W=440.00n L=60.00n
MM1 m net_0157 VDD VNW P12LL W=550.00n L=60.00n
.ENDS SDXHSV4
****Sub-Circuit for SEDGRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNHSV1 CK D E Q QN RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM64 QN s VSS VPW N12LL W=290.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=290.00n L=60.00n
MM17 sp s VSS VPW N12LL W=280.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM65 QN s VDD VNW P12LL W=440.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=440.00n L=60.00n
MM18 sp s VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNHSV1
****Sub-Circuit for SEDGRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNHSV2 CK D E Q QN RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM64 QN s VSS VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=430.00n L=60.00n
MM17 sp s VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM65 QN s VDD VNW P12LL W=650.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=650.00n L=60.00n
MM18 sp s VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNHSV2
****Sub-Circuit for SEDGRNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNHSV4 CK D E Q QN RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM64 QN s VSS VPW N12LL W=860.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=860.00n L=60.00n
MM17 sp s VSS VPW N12LL W=400.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM65 QN s VDD VNW P12LL W=1.3u L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=1.3u L=60.00n
MM18 sp s VDD VNW P12LL W=480.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNHSV4
****Sub-Circuit for SEDGRNQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNQHSV1 CK D E Q RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=290.00n L=60.00n
MM17 sp s VSS VPW N12LL W=220.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=440.00n L=60.00n
MM18 sp s VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNQHSV1
****Sub-Circuit for SEDGRNQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNQHSV2 CK D E Q RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=240.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=430.00n L=60.00n
MM17 sp s VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=360.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=650.00n L=60.00n
MM18 sp s VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNQHSV2
****Sub-Circuit for SEDGRNQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDGRNQHSV4 CK D E Q RN SE SI VDD VSS
MM55 m c s VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net_0157 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM62 net_0157 cn pm VPW N12LL W=400.00n L=60.00n
MM40 net_0157 sen net_0149 VPW N12LL W=430.00n L=60.00n
MM41 net_0149 s net_0164 VPW N12LL W=430.00n L=60.00n
MM59 net0172 E net0175 VPW N12LL W=430.00n L=60.00n
MM42 net0175 RN VSS VPW N12LL W=430.00n L=60.00n
MM58 net_0164 en net0175 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn s VPW N12LL W=200.00n L=60.00n
MM23 VSS sp net48 VPW N12LL W=200.00n L=60.00n
MM22 Q sp VSS VPW N12LL W=860.00n L=60.00n
MM17 sp s VSS VPW N12LL W=310.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0157 sen net69 VPW N12LL W=430.00n L=60.00n
MM7 net69 D net0172 VPW N12LL W=430.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM56 m cn s VNW P12LL W=650.00n L=60.00n
MM54 net0255 SE VDD VNW P12LL W=200.00n L=60.00n
MM53 net0267 E VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM63 net_0157 c pm VNW P12LL W=600.00n L=60.00n
MM37 net_0157 SE net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 s net0267 VNW P12LL W=500.00n L=60.00n
MM39 net_0157 RN net0255 VNW P12LL W=200.00n L=60.00n
MM57 net0279 en VDD VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD sp net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c s VNW P12LL W=300.00n L=60.00n
MM21 Q sp VDD VNW P12LL W=1.3u L=60.00n
MM18 sp s VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 SE net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 D net0279 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDGRNQHSV4
****Sub-Circuit for SEDHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDHSV1 CK D E Q QN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=300.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=300.00n L=60.00n
MM68 QN s VSS VPW N12LL W=290.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=420.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=420.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=420.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=300.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=420.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=420.00n L=60.00n
MM0 m pm VSS VPW N12LL W=400.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=300.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=300.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM69 QN s VDD VNW P12LL W=440.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=500.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=500.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=500.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=500.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=500.00n L=60.00n
MM1 m pm VDD VNW P12LL W=600.00n L=60.00n
.ENDS SEDHSV1
****Sub-Circuit for SEDHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDHSV2 CK D E Q QN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 QN s VSS VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=400.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=400.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM69 QN s VDD VNW P12LL W=650.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=420.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDHSV2
****Sub-Circuit for SEDHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDHSV4 CK D E Q QN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 QN s VSS VPW N12LL W=860.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=390.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=440.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=440.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM69 QN s VDD VNW P12LL W=1.3u L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=500.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDHSV4
****Sub-Circuit for SEDQHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDQHSV1 CK D E Q SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=300.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=300.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=300.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=300.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDQHSV1
****Sub-Circuit for SEDQHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDQHSV2 CK D E Q SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=400.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=400.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDQHSV2
****Sub-Circuit for SEDQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDQHSV4 CK D E Q SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=400.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SI VSS VPW N12LL W=200.00n L=60.00n
MM45 net0171 SE net_0152 VPW N12LL W=200.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=400.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=400.00n L=60.00n
MM58 net_0164 sen VSS VPW N12LL W=400.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=400.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=400.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=420.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=420.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=570.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=570.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 sen net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 SI VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=570.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=570.00n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=570.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=570.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDQHSV4
****Sub-Circuit for SEDRNHSV1, Fri May 27 10:36:55 CST 2011****
.SUBCKT SEDRNHSV1 CK D E Q QN RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=390.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM73 QN s VSS VPW N12LL W=290.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=250.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=250.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=275.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=250.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=270.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM74 QN s VDD VNW P12LL W=440.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=355.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=390.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=390.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=380.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=400.00n L=60.00n
.ENDS SEDRNHSV1
****Sub-Circuit for SEDRNHSV2, Thu May 26 17:37:04 CST 2011****
.SUBCKT SEDRNHSV2 CK D E Q QN RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=390.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM73 QN s VSS VPW N12LL W=430.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=250.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=250.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=275.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=290.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=360.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM74 QN s VDD VNW P12LL W=650.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=355.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=390.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=390.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=440.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=540.00n L=60.00n
.ENDS SEDRNHSV2
****Sub-Circuit for SEDRNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDRNHSV4 CK D E Q QN RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=360.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=360.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM73 QN s VSS VPW N12LL W=860.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=250.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=250.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=275.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=430.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=400.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=400.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=470.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=470.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM74 QN s VDD VNW P12LL W=1.3u L=60.00n
MM53 net0267 SE VDD VNW P12LL W=355.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=390.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=390.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=650.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=440.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=600.00n L=60.00n
.ENDS SEDRNHSV4
****Sub-Circuit for SEDRNQHSV1, Thu May 26 14:31:08 CST 2011****
.SUBCKT SEDRNQHSV1 CK D E Q RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=390.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=240.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=240.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=300.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=385.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=385.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=370.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=380.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=380.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDRNQHSV1
****Sub-Circuit for SEDRNQHSV2, Thu May 26 13:48:52 CST 2011****
.SUBCKT SEDRNQHSV2 CK D E Q RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=240.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=240.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=290.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=310.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=380.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=380.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=380.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDRNQHSV2
****Sub-Circuit for SEDRNQHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SEDRNQHSV4 CK D E Q RDN SE SI VDD VSS
MM39 ps c net_0155 VPW N12LL W=390.00n L=60.00n
MM65 net_0155 m VSS VPW N12LL W=400.00n L=60.00n
MM68 net0157 RDN VSS VPW N12LL W=310.00n L=60.00n
MM60 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM70 VSS RDN net0183 VPW N12LL W=200.00n L=60.00n
MM46 net_0152 SE net0157 VPW N12LL W=240.00n L=60.00n
MM45 net0171 SI net_0152 VPW N12LL W=240.00n L=60.00n
MM40 net0171 s net_0149 VPW N12LL W=310.00n L=60.00n
MM41 net_0149 en net_0164 VPW N12LL W=310.00n L=60.00n
MM71 VSS RDN net0163 VPW N12LL W=200.00n L=60.00n
MM58 net_0164 sen net0157 VPW N12LL W=300.00n L=60.00n
MM63 pm cn net0171 VPW N12LL W=400.00n L=60.00n
MM31 en E VSS VPW N12LL W=200.00n L=60.00n
MM30 c cn VSS VPW N12LL W=300.00n L=60.00n
MM27 cn CK VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 net0163 s net48 VPW N12LL W=200.00n L=60.00n
MM22 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=200.00n L=60.00n
MM12 net52 c pm VPW N12LL W=200.00n L=60.00n
MM11 net0183 m net52 VPW N12LL W=200.00n L=60.00n
MM9 net0171 D net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 E net_0164 VPW N12LL W=310.00n L=60.00n
MM0 m pm VSS VPW N12LL W=430.00n L=60.00n
MM66 ps cn net_0153 VNW P12LL W=415.00n L=60.00n
MM67 net_0153 m VDD VNW P12LL W=415.00n L=60.00n
MM64 pm c net_0157 VNW P12LL W=520.00n L=60.00n
MM53 net0267 SE VDD VNW P12LL W=390.00n L=60.00n
MM61 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM51 net_0157 SI net_0247 VNW P12LL W=300.00n L=60.00n
MM50 net_0247 sen VDD VNW P12LL W=300.00n L=60.00n
MM37 net_0157 s net_0228 VNW P12LL W=380.00n L=60.00n
MM38 net_0228 E net0267 VNW P12LL W=380.00n L=60.00n
MM69 pm RDN VDD VNW P12LL W=300.0n L=60.00n
MM72 ps RDN VDD VNW P12LL W=300.0n L=60.00n
MM32 en E VDD VNW P12LL W=300.00n L=60.00n
MM29 c cn VDD VNW P12LL W=450.00n L=60.00n
MM28 cn CK VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM21 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=300.00n L=60.00n
MM14 net117 cn pm VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0157 D net128 VNW P12LL W=390.00n L=60.00n
MM8 net128 en net0267 VNW P12LL W=390.00n L=60.00n
MM1 m pm VDD VNW P12LL W=650.00n L=60.00n
.ENDS SEDRNQHSV4
****Sub-Circuit for SNDHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDHSV1 CKN D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=290.00n L=60.00n
MM46 net_0107 SE VSS VPW N12LL W=250.00n L=60.00n
MM45 net_0163 SI net_0107 VPW N12LL W=250.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=230.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=230.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=250.00n L=60.00n
MM30 cn c VSS VPW N12LL W=250.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=290.00n L=60.00n
MM17 s ps VSS VPW N12LL W=240.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=250.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=250.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=270.00n L=60.00n
MM53 QN s VDD VNW P12LL W=440.00n L=60.00n
MM51 net128 SI net_0174 VNW P12LL W=650.00n L=60.00n
MM50 net_0174 SEN VDD VNW P12LL W=650.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=380.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=440.00n L=60.00n
MM18 s ps VDD VNW P12LL W=360.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=650.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=650.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=650.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=400.00n L=60.00n
.ENDS SNDHSV1
****Sub-Circuit for SNDHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDHSV2 CKN D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=430.00n L=60.00n
MM46 net_0107 SE VSS VPW N12LL W=250.00n L=60.00n
MM45 net_0163 SI net_0107 VPW N12LL W=250.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=230.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=230.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=250.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=430.00n L=60.00n
MM17 s ps VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=250.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=250.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=390.00n L=60.00n
MM53 QN s VDD VNW P12LL W=650.00n L=60.00n
MM51 net128 SI net_0174 VNW P12LL W=650.00n L=60.00n
MM50 net_0174 SEN VDD VNW P12LL W=650.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=650.00n L=60.00n
MM18 s ps VDD VNW P12LL W=440.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=650.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=650.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=650.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=580.00n L=60.00n
.ENDS SNDHSV2
****Sub-Circuit for SNDHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDHSV4 CKN D Q QN SE SI VDD VSS
MM52 QN s VSS VPW N12LL W=860.00n L=60.00n
MM46 net_0107 SE VSS VPW N12LL W=260.00n L=60.00n
MM45 net_0163 SI net_0107 VPW N12LL W=260.00n L=60.00n
MM39 ps c net_099 VPW N12LL W=250.00n L=60.00n
MM48 SEN SE VSS VPW N12LL W=200.00n L=60.00n
MM40 net_099 m VSS VPW N12LL W=250.00n L=60.00n
MM43 net_0123 SEN VSS VPW N12LL W=260.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=290.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q ps VSS VPW N12LL W=860.00n L=60.00n
MM17 s ps VSS VPW N12LL W=360.00n L=60.00n
MM12 net52 c net_0159 VPW N12LL W=200.00n L=60.00n
MM11 VSS m net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0159 cn net_0163 VPW N12LL W=260.00n L=60.00n
MM42 net_0163 D net_0123 VPW N12LL W=260.00n L=60.00n
MM0 m net_0159 VSS VPW N12LL W=430.00n L=60.00n
MM53 QN s VDD VNW P12LL W=1.3u L=60.00n
MM51 net128 SI net_0174 VNW P12LL W=650.00n L=60.00n
MM50 net_0174 SEN VDD VNW P12LL W=650.00n L=60.00n
MM38 ps cn net_0158 VNW P12LL W=650.00n L=60.00n
MM41 net_0158 m VDD VNW P12LL W=650.00n L=60.00n
MM49 SEN SE VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q ps VDD VNW P12LL W=1.3u L=60.00n
MM18 s ps VDD VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0159 VNW P12LL W=300.00n L=60.00n
MM13 VDD m net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0159 c net128 VNW P12LL W=650.00n L=60.00n
MM44 net_0230 SE VDD VNW P12LL W=650.00n L=60.00n
MM47 net128 D net_0230 VNW P12LL W=650.00n L=60.00n
MM1 m net_0159 VDD VNW P12LL W=650.00n L=60.00n
.ENDS SNDHSV4
****Sub-Circuit for SNDRNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRNHSV1 CKN D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=290.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=300.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=300.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=300.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=300.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=300.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM39 s ps net_099 VPW N12LL W=360.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=360.00n L=60.00n
MM30 cn c VSS VPW N12LL W=300.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=300.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=440.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=500.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM38 s ps VDD VNW P12LL W=390.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=390.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=450.00n L=60.00n
MM29 cn c VDD VNW P12LL W=450.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=450.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=450.00n L=60.00n
.ENDS SNDRNHSV1
****Sub-Circuit for SNDRNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRNHSV2 CKN D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=430.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=350.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=350.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=300.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=290.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=300.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=190.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM39 s ps net_099 VPW N12LL W=360.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=360.00n L=60.00n
MM30 cn c VSS VPW N12LL W=300.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=190.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=190.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=300.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=650.00n L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=450.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=450.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM38 s ps VDD VNW P12LL W=390.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=390.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=445.00n L=60.00n
MM29 cn c VDD VNW P12LL W=450.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn ps VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=450.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=450.00n L=60.00n
.ENDS SNDRNHSV2
****Sub-Circuit for SNDRNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRNHSV4 CKN D Q QN RDN SE SI VDD VSS
MM53 QN ps VSS VPW N12LL W=860.00n L=60.00n
MM45 net_0137 sen net_0133 VPW N12LL W=350.00n L=60.00n
MM46 net_0133 D net_0104 VPW N12LL W=350.00n L=60.00n
MM3 net_0154 c ps VPW N12LL W=300.00n L=60.00n
MM49 net_0137 cn net_0132 VPW N12LL W=300.00n L=60.00n
MM44 net_0104 RDN VSS VPW N12LL W=300.00n L=60.00n
MM42 VSS RDN net_0119 VPW N12LL W=200.00n L=60.00n
MM51 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM39 s ps net_099 VPW N12LL W=380.00n L=60.00n
MM40 net_099 RDN VSS VPW N12LL W=380.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=300.00n L=60.00n
MM24 net48 cn ps VPW N12LL W=200.00n L=60.00n
MM23 VSS s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0132 VPW N12LL W=200.00n L=60.00n
MM11 net_0119 net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0137 SE net69 VPW N12LL W=300.00n L=60.00n
MM7 net69 SI net_0104 VPW N12LL W=300.00n L=60.00n
MM0 net_0154 net_0132 VSS VPW N12LL W=300.00n L=60.00n
MM54 QN ps VDD VNW P12LL W=1.3u L=60.00n
MM47 net_0137 SE net_0212 VNW P12LL W=500.00n L=60.00n
MM48 net_0212 D VDD VNW P12LL W=500.00n L=60.00n
MM43 net_0132 RDN VDD VNW P12LL W=300.00n L=60.00n
MM52 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM38 s ps VDD VNW P12LL W=350.00n L=60.00n
MM41 s RDN VDD VNW P12LL W=300.00n L=60.00n
MM50 net_0137 c net_0132 VNW P12LL W=450.00n L=60.00n
MM29 cn c VDD VNW P12LL W=530.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=450.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c ps VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn ps VNW P12LL W=450.00n L=60.00n
MM14 net117 cn net_0132 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0137 sen net128 VNW P12LL W=450.00n L=60.00n
MM8 net128 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0132 VDD VNW P12LL W=450.00n L=60.00n
.ENDS SNDRNHSV4
****Sub-Circuit for SNDRSNHSV1, Mon May 30 19:16:43 CST 2011****
.SUBCKT SNDRSNHSV1 CKN D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=270.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=340.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=300.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=300.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=300.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=300.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=450.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=450.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=500.00n L=60.00n
MM29 cn c VDD VNW P12LL W=540.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=540.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=540.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=500.00n L=60.00n
.ENDS SNDRSNHSV1
****Sub-Circuit for SNDRSNHSV2, Mon May 30 17:13:17 CST 2011****
.SUBCKT SNDRSNHSV2 CKN D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=270.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=340.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=340.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=300.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=300.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=300.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=300.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=450.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=450.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=500.00n L=60.00n
MM29 cn c VDD VNW P12LL W=540.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=540.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=540.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=500.00n L=60.00n
.ENDS SNDRSNHSV2
****Sub-Circuit for SNDRSNHSV4, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDRSNHSV4 CKN D Q QN RDN SDN SE SI VDD VSS
MM58 sen SE VSS VPW N12LL W=300.00n L=60.00n
MM45 R RDN VSS VPW N12LL W=270.00n L=60.00n
MM47 net_0154 R L VPW N12LL W=200.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=350.00n L=60.00n
MM48 L SDN VSS VPW N12LL W=360.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 net_0140 cn net_0139 VPW N12LL W=300.00n L=60.00n
MM51 net_0140 sen net_0144 VPW N12LL W=320.00n L=60.00n
MM40 net43 R L VPW N12LL W=200.00n L=60.00n
MM52 net_0144 D VSS VPW N12LL W=320.00n L=60.00n
MM9 net_0140 SE net_0156 VPW N12LL W=300.00n L=60.00n
MM7 net_0156 SI VSS VPW N12LL W=300.00n L=60.00n
MM30 cn c VSS VPW N12LL W=360.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 L s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0139 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM0 net_0154 net_0139 L VPW N12LL W=360.00n L=60.00n
MM59 sen SE VDD VNW P12LL W=450.00n L=60.00n
MM46 R RDN VDD VNW P12LL W=430.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM10 net_0140 sen net_0223 VNW P12LL W=450.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM57 net_0140 c net_0139 VNW P12LL W=450.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=390.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM44 H R VDD VNW P12LL W=540.00n L=60.00n
MM29 cn c VDD VNW P12LL W=540.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 H s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=540.00n L=60.00n
MM14 net117 cn net_0139 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM54 net_0140 SE net_0231 VNW P12LL W=540.00n L=60.00n
MM55 net_0231 D VDD VNW P12LL W=540.00n L=60.00n
MM8 net_0223 SI VDD VNW P12LL W=450.00n L=60.00n
MM1 net_0154 net_0139 H VNW P12LL W=540.00n L=60.00n
.ENDS SNDRSNHSV4
****Sub-Circuit for SNDSNHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDSNHSV1 CKN D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=220.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=220.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=220.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=220.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=200.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=290.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=240.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=250.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=290.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=220.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=430.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=480.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=480.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=480.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=480.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=440.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=360.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=380.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=440.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=480.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=500.00n L=60.00n
.ENDS SNDSNHSV1
****Sub-Circuit for SNDSNHSV2, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT SNDSNHSV2 CKN D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=220.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=220.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=220.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=220.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=250.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=430.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=290.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=290.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=200.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=430.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=220.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=430.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=480.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=480.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=480.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=480.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=650.00n L=60.00n
MM38 s net43 VDD VNW P12LL W=440.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=440.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=300.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=650.00n L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=480.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=500.00n L=60.00n
.ENDS SNDSNHSV2
****Sub-Circuit for SNDSNHSV4, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT SNDSNHSV4 CKN D Q QN SDN SE SI VDD VSS
MM51 N11 sen net_0129 VPW N12LL W=250.00n L=60.00n
MM52 net_0129 D VSS VPW N12LL W=250.00n L=60.00n
MM54 N11 SE net_0121 VPW N12LL W=250.00n L=60.00n
MM55 net_0121 SI VSS VPW N12LL W=250.00n L=60.00n
MM3 net_0154 c net43 VPW N12LL W=430.00n L=60.00n
MM48 net_0132 SDN VSS VPW N12LL W=430.00n L=60.00n
MM49 QN net43 VSS VPW N12LL W=860.00n L=60.00n
MM39 s net43 VSS VPW N12LL W=380.00n L=60.00n
MM56 sen SE VSS VPW N12LL W=200.00n L=60.00n
MM30 cn c VSS VPW N12LL W=390.00n L=60.00n
MM27 c CKN VSS VPW N12LL W=270.00n L=60.00n
MM24 net48 cn net43 VPW N12LL W=200.00n L=60.00n
MM23 net_0132 s net48 VPW N12LL W=200.00n L=60.00n
MM19 Q s VSS VPW N12LL W=860.00n L=60.00n
MM12 net52 c net_0181 VPW N12LL W=200.00n L=60.00n
MM11 VSS net_0154 net52 VPW N12LL W=200.00n L=60.00n
MM9 net_0181 cn N11 VPW N12LL W=250.00n L=60.00n
MM0 net_0154 net_0181 net_0132 VPW N12LL W=430.00n L=60.00n
MM57 N7 sen net_0204 VNW P12LL W=480.00n L=60.00n
MM59 N7 SE net_0200 VNW P12LL W=480.00n L=60.00n
MM60 net_0200 D VDD VNW P12LL W=480.00n L=60.00n
MM61 net_0204 SI VDD VNW P12LL W=480.00n L=60.00n
MM43 net_0154 SDN VDD VNW P12LL W=300.00n L=60.00n
MM62 sen SE VDD VNW P12LL W=300.00n L=60.00n
MM50 QN net43 VDD VNW P12LL W=1.3u L=60.00n
MM38 s net43 VDD VNW P12LL W=540.00n L=60.00n
MM41 net43 SDN VDD VNW P12LL W=300.00n L=60.00n
MM29 cn c VDD VNW P12LL W=470.00n L=60.00n
MM28 c CKN VDD VNW P12LL W=430.00n L=60.00n
MM26 VDD s net109 VNW P12LL W=300.00n L=60.00n
MM25 net109 c net43 VNW P12LL W=300.00n L=60.00n
MM20 Q s VDD VNW P12LL W=1.3u L=60.00n
MM4 net_0154 cn net43 VNW P12LL W=500.00n L=60.00n
MM14 net117 cn net_0181 VNW P12LL W=300.00n L=60.00n
MM13 VDD net_0154 net117 VNW P12LL W=300.00n L=60.00n
MM10 net_0181 c N7 VNW P12LL W=480.00n L=60.00n
MM1 net_0154 net_0181 VDD VNW P12LL W=500.00n L=60.00n
.ENDS SNDSNHSV4
****Sub-Circuit for TBUFHSV0, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT TBUFHSV0 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=200.00n L=60.00n
MM44 net080 oen VSS VPW N12LL W=200.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=200.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=200.00n L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=200.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=200.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=300.00n L=60.00n
MM28 oen OE VDD VNW P12LL W=300.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=300.00n L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=300.00n L=60.00n
.ENDS TBUFHSV0
****Sub-Circuit for TBUFHSV1, Wed Dec  8 11:21:18 CST 2010****
.SUBCKT TBUFHSV1 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=200.00n L=60.00n
MM44 net080 oen VSS VPW N12LL W=200.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=200.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=300.00n L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=200.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=200.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=300.00n L=60.00n
MM28 oen OE VDD VNW P12LL W=300.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=450.00n L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=300.00n L=60.00n
.ENDS TBUFHSV1
****Sub-Circuit for TBUFHSV12, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT TBUFHSV12 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=830.00n L=60.00n
MM44 net080 oen VSS VPW N12LL W=300.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=260.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=2.49u L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=430.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=450.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=1.27u L=60.00n
MM28 oen OE VDD VNW P12LL W=400.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=3.81u L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=650.00n L=60.00n
.ENDS TBUFHSV12
****Sub-Circuit for TBUFHSV16, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT TBUFHSV16 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=1.14u L=60.00n
MM44 net080 oen VSS VPW N12LL W=350.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=400.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=3.32u L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=830.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=520.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=1.68u L=60.00n
MM28 oen OE VDD VNW P12LL W=600.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=5.08u L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=1.27u L=60.00n
.ENDS TBUFHSV16
****Sub-Circuit for TBUFHSV2, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT TBUFHSV2 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=200.00n L=60.00n
MM44 net080 oen VSS VPW N12LL W=200.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=200.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=430.00n L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=200.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=200.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=300.00n L=60.00n
MM28 oen OE VDD VNW P12LL W=300.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=650.00n L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=300.00n L=60.00n
.ENDS TBUFHSV2
****Sub-Circuit for TBUFHSV20, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT TBUFHSV20 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=1.6u L=60.00n
MM44 net080 oen VSS VPW N12LL W=415.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=415.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=4.15u L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=830.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=635.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=2.4u L=60.00n
MM28 oen OE VDD VNW P12LL W=635.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=6.35u L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=1.27u L=60.00n
.ENDS TBUFHSV20
****Sub-Circuit for TBUFHSV24, Fri Dec 10 10:21:29 CST 2010****
.SUBCKT TBUFHSV24 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=1.68u L=60.00n
MM44 net080 oen VSS VPW N12LL W=415.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=415.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=4.98u L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=830.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=635.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=2.52u L=60.00n
MM28 oen OE VDD VNW P12LL W=635.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=7.62u L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=1.27u L=60.00n
.ENDS TBUFHSV24
****Sub-Circuit for TBUFHSV3, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT TBUFHSV3 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=200.00n L=60.00n
MM44 net080 oen VSS VPW N12LL W=200.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=200.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=660.00n L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=200.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=200.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=300.00n L=60.00n
MM28 oen OE VDD VNW P12LL W=300.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=1u L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=300.00n L=60.00n
.ENDS TBUFHSV3
****Sub-Circuit for TBUFHSV4, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT TBUFHSV4 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=520.00n L=60.00n
MM44 net080 oen VSS VPW N12LL W=200.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=200.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=860.00n L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=520.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=200.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=520.00n L=60.00n
MM28 oen OE VDD VNW P12LL W=300.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=1.3u L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=520.00n L=60.00n
.ENDS TBUFHSV4
****Sub-Circuit for TBUFHSV6, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT TBUFHSV6 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=415.00n L=60.00n
MM44 net080 oen VSS VPW N12LL W=200.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=200.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=1.245u L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=420.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=205.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=635.00n L=60.00n
MM28 oen OE VDD VNW P12LL W=305.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=1.905u L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=650.00n L=60.00n
.ENDS TBUFHSV6
****Sub-Circuit for TBUFHSV8, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT TBUFHSV8 I OE Z VDD VSS
MM43 net080 I VSS VPW N12LL W=680.00n L=60.00n
MM44 net080 oen VSS VPW N12LL W=200.00n L=60.00n
MM27 oen OE VSS VPW N12LL W=200.00n L=60.00n
MM22 Z net080 VSS VPW N12LL W=1.66u L=60.00n
MM36 net080 OE net_0163 VPW N12LL W=430.00n L=60.00n
MM45 net_0163 OE VDD VNW P12LL W=300.00n L=60.00n
MM46 net_0163 I VDD VNW P12LL W=1.04u L=60.00n
MM28 oen OE VDD VNW P12LL W=300.00n L=60.00n
MM21 Z net_0163 VDD VNW P12LL W=2.54u L=60.00n
MM39 net080 oen net_0163 VNW P12LL W=650.00n L=60.00n
.ENDS TBUFHSV8
****Sub-Circuit for XNOR2HSV0, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR2HSV0 A1 A2 ZN VDD VSS
MM57 ZN xa1a2 VSS VPW N12LL W=200.00n L=60.00n
MM47 a2n A1 xa1a2 VPW N12LL W=200.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM55 a2nn a2n VSS VPW N12LL W=200.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=260.00n L=60.00n
MM36 a2nn a1n xa1a2 VPW N12LL W=200.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=300.00n L=60.00n
MM58 ZN xa1a2 VDD VNW P12LL W=300.00n L=60.00n
MM48 a2n a1n xa1a2 VNW P12LL W=300.00n L=60.00n
MM56 a2nn a2n VDD VNW P12LL W=300.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=400.0n L=60.00n
MM39 a2nn A1 xa1a2 VNW P12LL W=300.00n L=60.00n
.ENDS XNOR2HSV0
****Sub-Circuit for XNOR2HSV1, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR2HSV1 A1 A2 ZN VDD VSS
MM57 ZN xa1a2 VSS VPW N12LL W=290.00n L=60.00n
MM47 a2n A1 xa1a2 VPW N12LL W=250.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=210.00n L=60.00n
MM55 a2nn a2n VSS VPW N12LL W=260.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=350.00n L=60.00n
MM36 a2nn a1n xa1a2 VPW N12LL W=250.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=320.00n L=60.00n
MM58 ZN xa1a2 VDD VNW P12LL W=440.00n L=60.00n
MM48 a2n a1n xa1a2 VNW P12LL W=400.00n L=60.00n
MM56 a2nn a2n VDD VNW P12LL W=400.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=540.0n L=60.00n
MM39 a2nn A1 xa1a2 VNW P12LL W=400.00n L=60.00n
.ENDS XNOR2HSV1
****Sub-Circuit for XNOR2HSV2, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR2HSV2 A1 A2 ZN VDD VSS
MM57 ZN xa1a2 VSS VPW N12LL W=430.00n L=60.00n
MM47 a2n A1 xa1a2 VPW N12LL W=300.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=240.00n L=60.00n
MM55 a2nn a2n VSS VPW N12LL W=300.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=400.00n L=60.00n
MM36 a2nn a1n xa1a2 VPW N12LL W=300.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=360.00n L=60.00n
MM58 ZN xa1a2 VDD VNW P12LL W=650.00n L=60.00n
MM48 a2n a1n xa1a2 VNW P12LL W=450.00n L=60.00n
MM56 a2nn a2n VDD VNW P12LL W=450.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=600.0n L=60.00n
MM39 a2nn A1 xa1a2 VNW P12LL W=450.00n L=60.00n
.ENDS XNOR2HSV2
****Sub-Circuit for XNOR2HSV4, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR2HSV4 A1 A2 ZN VDD VSS
MM57 ZN xa1a2 VSS VPW N12LL W=860.00n L=60.00n
MM47 a2n A1 xa1a2 VPW N12LL W=390.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=340.00n L=60.00n
MM55 a2nn a2n VSS VPW N12LL W=430.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=580.00n L=60.00n
MM36 a2nn a1n xa1a2 VPW N12LL W=390.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=520.00n L=60.00n
MM58 ZN xa1a2 VDD VNW P12LL W=1.3u L=60.00n
MM48 a2n a1n xa1a2 VNW P12LL W=600.00n L=60.00n
MM56 a2nn a2n VDD VNW P12LL W=650.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=860.0n L=60.00n
MM39 a2nn A1 xa1a2 VNW P12LL W=600.00n L=60.00n
.ENDS XNOR2HSV4
****Sub-Circuit for XNOR3HSV0, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR3HSV0 A1 A2 A3 ZN VDD VSS
MM47 xa1a2 a3n xa1a2a3 VPW N12LL W=200.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=260.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=200.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=260.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=260.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=200.00n L=60.00n
MM67 ZN xa1a2a3 VSS VPW N12LL W=200.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=200.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=200.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=320.00n L=60.00n
MM36 xna1a2 A3 xa1a2a3 VPW N12LL W=200.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=400.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=300.00n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=300.00n L=60.00n
MM48 xa1a2 A3 xa1a2a3 VNW P12LL W=300.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=400.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=400.00n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=300.00n L=60.00n
MM68 ZN xa1a2a3 VDD VNW P12LL W=300.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=300.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=470.00n L=60.00n
MM39 xna1a2 a3n xa1a2a3 VNW P12LL W=300.00n L=60.00n
.ENDS XNOR3HSV0
****Sub-Circuit for XNOR3HSV1, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR3HSV1 A1 A2 A3 ZN VDD VSS
MM47 xa1a2 a3n xa1a2a3 VPW N12LL W=240.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=320.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=240.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=320.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=320.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=240.00n L=60.00n
MM67 ZN xa1a2a3 VSS VPW N12LL W=300.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=210.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=240.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=380.00n L=60.00n
MM36 xna1a2 A3 xa1a2a3 VPW N12LL W=240.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=480.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=320.00n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=360.00n L=60.00n
MM48 xa1a2 A3 xa1a2a3 VNW P12LL W=360.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=480.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=480.00n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=360.00n L=60.00n
MM68 ZN xa1a2a3 VDD VNW P12LL W=450.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=360.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=560.00n L=60.00n
MM39 xna1a2 a3n xa1a2a3 VNW P12LL W=360.00n L=60.00n
.ENDS XNOR3HSV1
****Sub-Circuit for XNOR3HSV2, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR3HSV2 A1 A2 A3 ZN VDD VSS
MM47 xa1a2 a3n xa1a2a3 VPW N12LL W=300.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=400.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=300.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=400.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=400.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=300.00n L=60.00n
MM67 ZN xa1a2a3 VSS VPW N12LL W=430.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=240.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=300.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=400.00n L=60.00n
MM36 xna1a2 A3 xa1a2a3 VPW N12LL W=300.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=600.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=360.00n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=450.00n L=60.00n
MM48 xa1a2 A3 xa1a2a3 VNW P12LL W=450.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=600.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=600.00n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=450.00n L=60.00n
MM68 ZN xa1a2a3 VDD VNW P12LL W=650.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=450.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=620.00n L=60.00n
MM39 xna1a2 a3n xa1a2a3 VNW P12LL W=450.00n L=60.00n
.ENDS XNOR3HSV2
****Sub-Circuit for XNOR3HSV4, Mon May 30 15:54:44 CST 2011****
.SUBCKT XNOR3HSV4 A1 A2 A3 ZN VDD VSS
MM47 xa1a2 a3n xa1a2a3 VPW N12LL W=400.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=540.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=400.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=540.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=490.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=350.00n L=60.00n
MM67 ZN xa1a2a3 VSS VPW N12LL W=760.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=340.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=370.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=620.00n L=60.00n
MM36 xna1a2 A3 xa1a2a3 VPW N12LL W=400.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=800.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=500.00n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=600.00n L=60.00n
MM48 xa1a2 A3 xa1a2a3 VNW P12LL W=600.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=800.0n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=750.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=550.00n L=60.00n
MM68 ZN xa1a2a3 VDD VNW P12LL W=1.2u L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=600.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=930.00n L=60.00n
MM39 xna1a2 a3n xa1a2a3 VNW P12LL W=600.00n L=60.00n
.ENDS XNOR3HSV4
****Sub-Circuit for XNOR4HSV0, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR4HSV0 A1 A2 A3 A4 ZN VDD VSS
MM47 xa1a2 xna3a4 xa1a2a3a4 VPW N12LL W=200.00n L=60.00n
MM69 a4n A4 VSS VPW N12LL W=320.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=260.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=200.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=260.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=260.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=200.00n L=60.00n
MM67 ZN xa1a2a3a4 VSS VPW N12LL W=200.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=260.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=200.00n L=60.00n
MM71 a3nn a3n VSS VPW N12LL W=200.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=320.00n L=60.00n
MM73 a3n a4n xna3a4 VPW N12LL W=260.00n L=60.00n
MM74 a3nn A4 xna3a4 VPW N12LL W=200.00n L=60.00n
MM75 a3n A4 xa3a4 VPW N12LL W=260.00n L=60.00n
MM76 a3nn a4n xa3a4 VPW N12LL W=200.00n L=60.00n
MM36 xna1a2 xa3a4 xa1a2a3a4 VPW N12LL W=200.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=400.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=400.0n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=300.00n L=60.00n
MM48 xa1a2 xa3a4 xa1a2a3a4 VNW P12LL W=300.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=400.0n L=60.00n
MM70 a4n A4 VDD VNW P12LL W=470.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=400.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=300.00n L=60.00n
MM68 ZN xa1a2a3a4 VDD VNW P12LL W=300.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=300.00n L=60.00n
MM72 a3nn a3n VDD VNW P12LL W=300.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=470.00n L=60.00n
MM77 a3n A4 xna3a4 VNW P12LL W=400.0n L=60.00n
MM78 a3nn a4n xna3a4 VNW P12LL W=300.00n L=60.00n
MM79 a3n a4n xa3a4 VNW P12LL W=400.0n L=60.00n
MM80 a3nn A4 xa3a4 VNW P12LL W=300.00n L=60.00n
MM39 xna1a2 xna3a4 xa1a2a3a4 VNW P12LL W=300.00n L=60.00n
.ENDS XNOR4HSV0
****Sub-Circuit for XNOR4HSV1, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR4HSV1 A1 A2 A3 A4 ZN VDD VSS
MM47 xa1a2 xna3a4 xa1a2a3a4 VPW N12LL W=240.00n L=60.00n
MM69 a4n A4 VSS VPW N12LL W=380.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=320.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=240.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=320.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=320.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=240.00n L=60.00n
MM67 ZN xa1a2a3a4 VSS VPW N12LL W=300.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=320.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=240.00n L=60.00n
MM71 a3nn a3n VSS VPW N12LL W=240.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=380.00n L=60.00n
MM73 a3n a4n xna3a4 VPW N12LL W=320.00n L=60.00n
MM74 a3nn A4 xna3a4 VPW N12LL W=240.00n L=60.00n
MM75 a3n A4 xa3a4 VPW N12LL W=320.00n L=60.00n
MM76 a3nn a4n xa3a4 VPW N12LL W=200.00n L=60.00n
MM36 xna1a2 xa3a4 xa1a2a3a4 VPW N12LL W=240.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=480.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=480.0n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=360.00n L=60.00n
MM48 xa1a2 xa3a4 xa1a2a3a4 VNW P12LL W=360.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=480.0n L=60.00n
MM70 a4n A4 VDD VNW P12LL W=560.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=480.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=360.00n L=60.00n
MM68 ZN xa1a2a3a4 VDD VNW P12LL W=450.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=360.00n L=60.00n
MM72 a3nn a3n VDD VNW P12LL W=360.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=560.00n L=60.00n
MM77 a3n A4 xna3a4 VNW P12LL W=480.0n L=60.00n
MM78 a3nn a4n xna3a4 VNW P12LL W=360.00n L=60.00n
MM79 a3n a4n xa3a4 VNW P12LL W=440.0n L=60.00n
MM80 a3nn A4 xa3a4 VNW P12LL W=360.00n L=60.00n
MM39 xna1a2 xna3a4 xa1a2a3a4 VNW P12LL W=360.00n L=60.00n
.ENDS XNOR4HSV1
****Sub-Circuit for XNOR4HSV2, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR4HSV2 A1 A2 A3 A4 ZN VDD VSS
MM47 xa1a2 xna3a4 xa1a2a3a4 VPW N12LL W=300.00n L=60.00n
MM69 a4n A4 VSS VPW N12LL W=400.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=400.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=300.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=400.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=380.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=300.00n L=60.00n
MM67 ZN xa1a2a3a4 VSS VPW N12LL W=430.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=400.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=300.00n L=60.00n
MM71 a3nn a3n VSS VPW N12LL W=300.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=400.00n L=60.00n
MM73 a3n a4n xna3a4 VPW N12LL W=400.00n L=60.00n
MM74 a3nn A4 xna3a4 VPW N12LL W=300.00n L=60.00n
MM75 a3n A4 xa3a4 VPW N12LL W=400.00n L=60.00n
MM76 a3nn a4n xa3a4 VPW N12LL W=295.00n L=60.00n
MM36 xna1a2 xa3a4 xa1a2a3a4 VPW N12LL W=300.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=600.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=600.0n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=450.00n L=60.00n
MM48 xa1a2 xa3a4 xa1a2a3a4 VNW P12LL W=450.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=600.0n L=60.00n
MM70 a4n A4 VDD VNW P12LL W=620.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=600.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=450.00n L=60.00n
MM68 ZN xa1a2a3a4 VDD VNW P12LL W=650.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=450.00n L=60.00n
MM72 a3nn a3n VDD VNW P12LL W=450.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=600.00n L=60.00n
MM77 a3n A4 xna3a4 VNW P12LL W=600.0n L=60.00n
MM78 a3nn a4n xna3a4 VNW P12LL W=450.00n L=60.00n
MM79 a3n a4n xa3a4 VNW P12LL W=595.0n L=60.00n
MM80 a3nn A4 xa3a4 VNW P12LL W=450.00n L=60.00n
MM39 xna1a2 xna3a4 xa1a2a3a4 VNW P12LL W=450.00n L=60.00n
.ENDS XNOR4HSV2
****Sub-Circuit for XNOR4HSV4, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XNOR4HSV4 A1 A2 A3 A4 ZN VDD VSS
MM47 xa1a2 xna3a4 xa1a2a3a4 VPW N12LL W=400.00n L=60.00n
MM69 a4n A4 VSS VPW N12LL W=620.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=540.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=400.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=540.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=400.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=400.00n L=60.00n
MM67 ZN xa1a2a3a4 VSS VPW N12LL W=860.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=540.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=400.00n L=60.00n
MM71 a3nn a3n VSS VPW N12LL W=400.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=620.00n L=60.00n
MM73 a3n a4n xna3a4 VPW N12LL W=540.00n L=60.00n
MM74 a3nn A4 xna3a4 VPW N12LL W=400.00n L=60.00n
MM75 a3n A4 xa3a4 VPW N12LL W=540.00n L=60.00n
MM76 a3nn a4n xa3a4 VPW N12LL W=370.00n L=60.00n
MM36 xna1a2 xa3a4 xa1a2a3a4 VPW N12LL W=400.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=800.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=800.0n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=600.00n L=60.00n
MM48 xa1a2 xa3a4 xa1a2a3a4 VNW P12LL W=600.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=800.0n L=60.00n
MM70 a4n A4 VDD VNW P12LL W=930.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=800.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=600.00n L=60.00n
MM68 ZN xa1a2a3a4 VDD VNW P12LL W=1.3u L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=600.00n L=60.00n
MM72 a3nn a3n VDD VNW P12LL W=600.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=790.00n L=60.00n
MM77 a3n A4 xna3a4 VNW P12LL W=800.0n L=60.00n
MM78 a3nn a4n xna3a4 VNW P12LL W=600.00n L=60.00n
MM79 a3n a4n xa3a4 VNW P12LL W=800.0n L=60.00n
MM80 a3nn A4 xa3a4 VNW P12LL W=600.00n L=60.00n
MM39 xna1a2 xna3a4 xa1a2a3a4 VNW P12LL W=600.00n L=60.00n
.ENDS XNOR4HSV4
****Sub-Circuit for XOR2HSV0, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR2HSV0 A1 A2 Z VDD VSS
MM57 Z xna1a2 VSS VPW N12LL W=200.00n L=60.00n
MM47 a2n a1n xna1a2 VPW N12LL W=200.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=200.00n L=60.00n
MM55 a2nn a2n VSS VPW N12LL W=200.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=250.00n L=60.00n
MM36 a2nn A1 xna1a2 VPW N12LL W=200.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=300.00n L=60.00n
MM58 Z xna1a2 VDD VNW P12LL W=300.00n L=60.00n
MM48 a2n A1 xna1a2 VNW P12LL W=300.00n L=60.00n
MM56 a2nn a2n VDD VNW P12LL W=300.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=450.0n L=60.00n
MM39 a2nn a1n xna1a2 VNW P12LL W=300.00n L=60.00n
.ENDS XOR2HSV0
****Sub-Circuit for XOR2HSV1, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR2HSV1 A1 A2 Z VDD VSS
MM57 Z xna1a2 VSS VPW N12LL W=290.00n L=60.00n
MM47 a2n a1n xna1a2 VPW N12LL W=220.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=210.00n L=60.00n
MM55 a2nn a2n VSS VPW N12LL W=260.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=350.00n L=60.00n
MM36 a2nn A1 xna1a2 VPW N12LL W=260.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=320.00n L=60.00n
MM58 Z xna1a2 VDD VNW P12LL W=440.00n L=60.00n
MM48 a2n A1 xna1a2 VNW P12LL W=400.00n L=60.00n
MM56 a2nn a2n VDD VNW P12LL W=400.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=540.0n L=60.00n
MM39 a2nn a1n xna1a2 VNW P12LL W=400.00n L=60.00n
.ENDS XOR2HSV1
****Sub-Circuit for XOR2HSV2, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR2HSV2 A1 A2 Z VDD VSS
MM57 Z xna1a2 VSS VPW N12LL W=430.00n L=60.00n
MM47 a2n a1n xna1a2 VPW N12LL W=280.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=240.00n L=60.00n
MM55 a2nn a2n VSS VPW N12LL W=270.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=400.00n L=60.00n
MM36 a2nn A1 xna1a2 VPW N12LL W=270.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=360.00n L=60.00n
MM58 Z xna1a2 VDD VNW P12LL W=650.00n L=60.00n
MM48 a2n A1 xna1a2 VNW P12LL W=450.00n L=60.00n
MM56 a2nn a2n VDD VNW P12LL W=450.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=600.0n L=60.00n
MM39 a2nn a1n xna1a2 VNW P12LL W=450.00n L=60.00n
.ENDS XOR2HSV2
****Sub-Circuit for XOR2HSV4, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR2HSV4 A1 A2 Z VDD VSS
MM57 Z xna1a2 VSS VPW N12LL W=860.00n L=60.00n
MM47 a2n a1n xna1a2 VPW N12LL W=360.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=340.00n L=60.00n
MM55 a2nn a2n VSS VPW N12LL W=430.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=550.00n L=60.00n
MM36 a2nn A1 xna1a2 VPW N12LL W=360.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=520.00n L=60.00n
MM58 Z xna1a2 VDD VNW P12LL W=1.3u L=60.00n
MM48 a2n A1 xna1a2 VNW P12LL W=635.00n L=60.00n
MM56 a2nn a2n VDD VNW P12LL W=635.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=860.0n L=60.00n
MM39 a2nn a1n xna1a2 VNW P12LL W=565.00n L=60.00n
.ENDS XOR2HSV4
****Sub-Circuit for XOR3HSV0, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR3HSV0 A1 A2 A3 Z VDD VSS
MM47 xa1a2 A3 xna1a2a3 VPW N12LL W=200.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=260.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=200.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=260.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=260.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=200.00n L=60.00n
MM67 Z xna1a2a3 VSS VPW N12LL W=200.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=200.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=200.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=320.00n L=60.00n
MM36 xna1a2 a3n xna1a2a3 VPW N12LL W=200.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=400.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=300.00n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=300.00n L=60.00n
MM48 xa1a2 a3n xna1a2a3 VNW P12LL W=300.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=400.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=400.00n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=300.00n L=60.00n
MM68 Z xna1a2a3 VDD VNW P12LL W=300.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=300.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=470.00n L=60.00n
MM39 xna1a2 A3 xna1a2a3 VNW P12LL W=300.00n L=60.00n
.ENDS XOR3HSV0
****Sub-Circuit for XOR3HSV1, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR3HSV1 A1 A2 A3 Z VDD VSS
MM47 xa1a2 A3 xna1a2a3 VPW N12LL W=240.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=320.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=240.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=320.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=320.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=240.00n L=60.00n
MM67 Z xna1a2a3 VSS VPW N12LL W=300.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=210.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=240.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=380.00n L=60.00n
MM36 xna1a2 a3n xna1a2a3 VPW N12LL W=240.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=480.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=320.00n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=360.00n L=60.00n
MM48 xa1a2 a3n xna1a2a3 VNW P12LL W=360.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=480.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=480.00n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=360.00n L=60.00n
MM68 Z xna1a2a3 VDD VNW P12LL W=450.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=360.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=560.00n L=60.00n
MM39 xna1a2 A3 xna1a2a3 VNW P12LL W=360.00n L=60.00n
.ENDS XOR3HSV1
****Sub-Circuit for XOR3HSV2, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR3HSV2 A1 A2 A3 Z VDD VSS
MM47 xa1a2 A3 xna1a2a3 VPW N12LL W=300.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=400.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=300.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=400.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=400.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=300.00n L=60.00n
MM67 Z xna1a2a3 VSS VPW N12LL W=430.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=240.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=300.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=400.00n L=60.00n
MM36 xna1a2 a3n xna1a2a3 VPW N12LL W=300.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=600.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=360.00n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=450.00n L=60.00n
MM48 xa1a2 a3n xna1a2a3 VNW P12LL W=450.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=600.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=600.00n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=450.00n L=60.00n
MM68 Z xna1a2a3 VDD VNW P12LL W=650.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=450.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=620.00n L=60.00n
MM39 xna1a2 A3 xna1a2a3 VNW P12LL W=450.00n L=60.00n
.ENDS XOR3HSV2
****Sub-Circuit for XOR3HSV4, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR3HSV4 A1 A2 A3 Z VDD VSS
MM47 xa1a2 A3 xna1a2a3 VPW N12LL W=400.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=540.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=400.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=540.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=510.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=400.00n L=60.00n
MM67 Z xna1a2a3 VSS VPW N12LL W=860.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=340.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=370.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=620.00n L=60.00n
MM36 xna1a2 a3n xna1a2a3 VPW N12LL W=400.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=800.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=500.00n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=600.00n L=60.00n
MM48 xa1a2 a3n xna1a2a3 VNW P12LL W=600.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=800.0n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=770.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=600.00n L=60.00n
MM68 Z xna1a2a3 VDD VNW P12LL W=1.3u L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=600.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=930.00n L=60.00n
MM39 xna1a2 A3 xna1a2a3 VNW P12LL W=600.00n L=60.00n
.ENDS XOR3HSV4
****Sub-Circuit for XOR4HSV0, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR4HSV0 A1 A2 A3 A4 Z VDD VSS
MM47 xa1a2 xa3a4 xna1a2a3a4 VPW N12LL W=200.00n L=60.00n
MM69 a4n A4 VSS VPW N12LL W=320.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=260.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=200.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=260.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=260.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=200.00n L=60.00n
MM67 Z xna1a2a3a4 VSS VPW N12LL W=200.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=260.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=200.00n L=60.00n
MM71 a3nn a3n VSS VPW N12LL W=200.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=320.00n L=60.00n
MM73 a3n a4n xna3a4 VPW N12LL W=260.00n L=60.00n
MM74 a3nn A4 xna3a4 VPW N12LL W=200.00n L=60.00n
MM75 a3n A4 xa3a4 VPW N12LL W=260.00n L=60.00n
MM76 a3nn a4n xa3a4 VPW N12LL W=200.00n L=60.00n
MM36 xna1a2 xna3a4 xna1a2a3a4 VPW N12LL W=200.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=400.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=400.0n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=300.00n L=60.00n
MM48 xa1a2 xna3a4 xna1a2a3a4 VNW P12LL W=300.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=400.0n L=60.00n
MM70 a4n A4 VDD VNW P12LL W=470.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=400.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=300.00n L=60.00n
MM68 Z xna1a2a3a4 VDD VNW P12LL W=300.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=300.00n L=60.00n
MM72 a3nn a3n VDD VNW P12LL W=300.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=470.00n L=60.00n
MM77 a3n A4 xna3a4 VNW P12LL W=400.0n L=60.00n
MM78 a3nn a4n xna3a4 VNW P12LL W=300.00n L=60.00n
MM79 a3n a4n xa3a4 VNW P12LL W=400.0n L=60.00n
MM80 a3nn A4 xa3a4 VNW P12LL W=300.00n L=60.00n
MM39 xna1a2 xa3a4 xna1a2a3a4 VNW P12LL W=300.00n L=60.00n
.ENDS XOR4HSV0
****Sub-Circuit for XOR4HSV1, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR4HSV1 A1 A2 A3 A4 Z VDD VSS
MM47 xa1a2 xa3a4 xna1a2a3a4 VPW N12LL W=240.00n L=60.00n
MM69 a4n A4 VSS VPW N12LL W=380.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=320.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=240.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=320.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=320.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=240.00n L=60.00n
MM67 Z xna1a2a3a4 VSS VPW N12LL W=300.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=320.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=240.00n L=60.00n
MM71 a3nn a3n VSS VPW N12LL W=240.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=380.00n L=60.00n
MM73 a3n a4n xna3a4 VPW N12LL W=320.00n L=60.00n
MM74 a3nn A4 xna3a4 VPW N12LL W=240.00n L=60.00n
MM75 a3n A4 xa3a4 VPW N12LL W=320.00n L=60.00n
MM76 a3nn a4n xa3a4 VPW N12LL W=240.00n L=60.00n
MM36 xna1a2 xna3a4 xna1a2a3a4 VPW N12LL W=240.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=480.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=480.0n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=360.00n L=60.00n
MM48 xa1a2 xna3a4 xna1a2a3a4 VNW P12LL W=360.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=480.0n L=60.00n
MM70 a4n A4 VDD VNW P12LL W=560.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=480.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=360.00n L=60.00n
MM68 Z xna1a2a3a4 VDD VNW P12LL W=450.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=360.00n L=60.00n
MM72 a3nn a3n VDD VNW P12LL W=360.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=560.00n L=60.00n
MM77 a3n A4 xna3a4 VNW P12LL W=480.0n L=60.00n
MM78 a3nn a4n xna3a4 VNW P12LL W=360.00n L=60.00n
MM79 a3n a4n xa3a4 VNW P12LL W=480.0n L=60.00n
MM80 a3nn A4 xa3a4 VNW P12LL W=360.00n L=60.00n
MM39 xna1a2 xa3a4 xna1a2a3a4 VNW P12LL W=360.00n L=60.00n
.ENDS XOR4HSV1
****Sub-Circuit for XOR4HSV2, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR4HSV2 A1 A2 A3 A4 Z VDD VSS
MM47 xa1a2 xa3a4 xna1a2a3a4 VPW N12LL W=300.00n L=60.00n
MM69 a4n A4 VSS VPW N12LL W=400.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=400.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=300.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=400.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=400.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=300.00n L=60.00n
MM67 Z xna1a2a3a4 VSS VPW N12LL W=430.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=400.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=300.00n L=60.00n
MM71 a3nn a3n VSS VPW N12LL W=300.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=400.00n L=60.00n
MM73 a3n a4n xna3a4 VPW N12LL W=400.00n L=60.00n
MM74 a3nn A4 xna3a4 VPW N12LL W=300.00n L=60.00n
MM75 a3n A4 xa3a4 VPW N12LL W=400.00n L=60.00n
MM76 a3nn a4n xa3a4 VPW N12LL W=295.00n L=60.00n
MM36 xna1a2 xna3a4 xna1a2a3a4 VPW N12LL W=300.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=600.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=600.0n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=450.00n L=60.00n
MM48 xa1a2 xna3a4 xna1a2a3a4 VNW P12LL W=450.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=600.0n L=60.00n
MM70 a4n A4 VDD VNW P12LL W=620.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=600.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=450.00n L=60.00n
MM68 Z xna1a2a3a4 VDD VNW P12LL W=650.00n L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=450.00n L=60.00n
MM72 a3nn a3n VDD VNW P12LL W=450.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=620.00n L=60.00n
MM77 a3n A4 xna3a4 VNW P12LL W=600.0n L=60.00n
MM78 a3nn a4n xna3a4 VNW P12LL W=450.00n L=60.00n
MM79 a3n a4n xa3a4 VNW P12LL W=595.0n L=60.00n
MM80 a3nn A4 xa3a4 VNW P12LL W=450.00n L=60.00n
MM39 xna1a2 xa3a4 xna1a2a3a4 VNW P12LL W=450.00n L=60.00n
.ENDS XOR4HSV2
****Sub-Circuit for XOR4HSV4, Wed Dec  8 11:21:19 CST 2010****
.SUBCKT XOR4HSV4 A1 A2 A3 A4 Z VDD VSS
MM47 xa1a2 xa3a4 xna1a2a3a4 VPW N12LL W=400.00n L=60.00n
MM69 a4n A4 VSS VPW N12LL W=620.00n L=60.00n
MM49 a1n A1 VSS VPW N12LL W=540.00n L=60.00n
MM60 a1nn A2 xna1a2 VPW N12LL W=400.00n L=60.00n
MM59 a1n a2n xna1a2 VPW N12LL W=540.00n L=60.00n
MM65 a1n A2 xa1a2 VPW N12LL W=510.00n L=60.00n
MM66 a1nn a2n xa1a2 VPW N12LL W=400.00n L=60.00n
MM67 Z xna1a2a3a4 VSS VPW N12LL W=860.00n L=60.00n
MM57 a3n A3 VSS VPW N12LL W=540.00n L=60.00n
MM55 a1nn a1n VSS VPW N12LL W=400.00n L=60.00n
MM71 a3nn a3n VSS VPW N12LL W=400.00n L=60.00n
MM53 a2n A2 VSS VPW N12LL W=620.00n L=60.00n
MM73 a3n a4n xna3a4 VPW N12LL W=540.00n L=60.00n
MM74 a3nn A4 xna3a4 VPW N12LL W=400.00n L=60.00n
MM75 a3n A4 xa3a4 VPW N12LL W=540.00n L=60.00n
MM76 a3nn a4n xa3a4 VPW N12LL W=400.00n L=60.00n
MM36 xna1a2 xna3a4 xna1a2a3a4 VPW N12LL W=400.00n L=60.00n
MM50 a1n A1 VDD VNW P12LL W=800.0n L=60.00n
MM58 a3n A3 VDD VNW P12LL W=800.0n L=60.00n
MM62 a1nn a2n xna1a2 VNW P12LL W=600.00n L=60.00n
MM48 xa1a2 xna3a4 xna1a2a3a4 VNW P12LL W=600.00n L=60.00n
MM61 a1n A2 xna1a2 VNW P12LL W=800.0n L=60.00n
MM70 a4n A4 VDD VNW P12LL W=930.00n L=60.00n
MM63 a1n a2n xa1a2 VNW P12LL W=770.0n L=60.00n
MM64 a1nn A2 xa1a2 VNW P12LL W=600.00n L=60.00n
MM68 Z xna1a2a3a4 VDD VNW P12LL W=1.3u L=60.00n
MM56 a1nn a1n VDD VNW P12LL W=600.00n L=60.00n
MM72 a3nn a3n VDD VNW P12LL W=600.00n L=60.00n
MM54 a2n A2 VDD VNW P12LL W=930.00n L=60.00n
MM77 a3n A4 xna3a4 VNW P12LL W=800.0n L=60.00n
MM78 a3nn a4n xna3a4 VNW P12LL W=600.00n L=60.00n
MM79 a3n a4n xa3a4 VNW P12LL W=800.0n L=60.00n
MM80 a3nn A4 xa3a4 VNW P12LL W=600.00n L=60.00n
MM39 xna1a2 xa3a4 xna1a2a3a4 VNW P12LL W=600.00n L=60.00n
.ENDS XOR4HSV4
