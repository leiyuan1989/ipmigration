* SPICE INPUT		Mon Sep 24 12:03:06 2018	ad01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d0
.subckt ad01d0 S VDD CO GND B CI A
M1 N_4 N_13 N_2 GND mn5  l=0.5u w=0.6u m=1
M2 N_2 CI N_3 GND mn5  l=0.5u w=0.6u m=1
M3 GND N_2 S GND mn5  l=0.5u w=0.6u m=1
M4 N_12 B GND GND mn5  l=0.5u w=0.6u m=1
M5 N_19 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_19 N_11 N_3 GND mn5  l=0.5u w=0.6u m=1
M7 N_3 N_19 N_11 GND mn5  l=0.5u w=0.6u m=1
M8 N_11 A GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 N_12 N_11 GND mn5  l=0.5u w=0.6u m=1
M10 N_12 N_11 N_4 GND mn5  l=0.5u w=0.6u m=1
M11 N_12 N_4 N_14 GND mn5  l=0.5u w=0.6u m=1
M12 N_13 N_3 N_14 GND mn5  l=0.5u w=0.6u m=1
M13 N_13 CI GND GND mn5  l=0.5u w=0.6u m=1
M14 CO N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_3 N_13 N_2 VDD mp5  l=0.42u w=0.62u m=1
M16 N_4 CI N_2 VDD mp5  l=0.42u w=0.62u m=1
M17 VDD N_2 S VDD mp5  l=0.42u w=0.62u m=1
M18 N_11 A VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_11 N_12 N_3 VDD mp5  l=0.42u w=0.62u m=1
M20 N_12 N_11 N_3 VDD mp5  l=0.42u w=0.62u m=1
M21 N_14 N_3 N_12 VDD mp5  l=0.42u w=0.62u m=1
M22 N_14 N_4 N_13 VDD mp5  l=0.42u w=0.62u m=1
M23 N_13 CI VDD VDD mp5  l=0.42u w=0.62u m=1
M24 VDD N_14 CO VDD mp5  l=0.42u w=0.62u m=1
M25 N_12 B VDD VDD mp5  l=0.42u w=0.62u m=1
M26 N_19 N_12 VDD VDD mp5  l=0.42u w=0.62u m=1
M27 N_19 N_11 N_4 VDD mp5  l=0.42u w=0.62u m=1
M28 N_11 N_19 N_4 VDD mp5  l=0.42u w=0.62u m=1
.ends ad01d0
* SPICE INPUT		Mon Sep 24 12:03:14 2018	ad01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d1
.subckt ad01d1 VDD CO S GND B A CI
M1 N_5 N_14 N_6 GND mn5  l=0.5u w=0.6u m=1
M2 N_14 N_6 N_5 GND mn5  l=0.5u w=0.6u m=1
M3 N_14 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_7 B GND GND mn5  l=0.5u w=0.6u m=1
M5 CO N_9 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_8 CI GND GND mn5  l=0.5u w=0.6u m=1
M7 N_8 N_5 N_9 GND mn5  l=0.5u w=0.6u m=1
M8 N_7 N_10 N_9 GND mn5  l=0.5u w=0.6u m=1
M9 N_7 N_6 N_10 GND mn5  l=0.5u w=0.6u m=1
M10 N_10 N_7 N_6 GND mn5  l=0.5u w=0.6u m=1
M11 N_6 A GND GND mn5  l=0.5u w=0.6u m=1
M12 GND N_17 S GND mn5  l=0.5u w=0.72u m=1
M13 N_17 CI N_5 GND mn5  l=0.5u w=0.6u m=1
M14 N_10 N_8 N_17 GND mn5  l=0.5u w=0.6u m=1
M15 CO N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_8 CI VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_9 N_10 N_8 VDD mp5  l=0.42u w=0.62u m=1
M18 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.62u m=1
M19 N_7 N_6 N_5 VDD mp5  l=0.42u w=0.62u m=1
M20 N_6 N_7 N_5 VDD mp5  l=0.42u w=0.62u m=1
M21 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_6 N_14 N_10 VDD mp5  l=0.42u w=0.62u m=1
M23 N_14 N_6 N_10 VDD mp5  l=0.42u w=0.62u m=1
M24 N_14 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_7 B VDD VDD mp5  l=0.42u w=0.62u m=1
M26 VDD N_17 S VDD mp5  l=0.42u w=0.96u m=1
M27 N_10 CI N_17 VDD mp5  l=0.42u w=0.62u m=1
M28 N_5 N_8 N_17 VDD mp5  l=0.42u w=0.62u m=1
.ends ad01d1
* SPICE INPUT		Mon Sep 24 12:03:23 2018	ad01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d2
.subckt ad01d2 VDD CO S GND B A CI
M1 N_5 N_14 N_6 GND mn5  l=0.5u w=0.6u m=1
M2 N_14 N_6 N_5 GND mn5  l=0.5u w=0.6u m=1
M3 N_14 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_7 B GND GND mn5  l=0.5u w=0.6u m=1
M5 CO N_9 GND GND mn5  l=0.5u w=0.98u m=1
M6 N_8 CI GND GND mn5  l=0.5u w=0.6u m=1
M7 N_8 N_5 N_9 GND mn5  l=0.5u w=0.6u m=1
M8 N_7 N_10 N_9 GND mn5  l=0.5u w=0.6u m=1
M9 N_7 N_6 N_10 GND mn5  l=0.5u w=0.6u m=1
M10 N_10 N_7 N_6 GND mn5  l=0.5u w=0.6u m=1
M11 N_6 A GND GND mn5  l=0.5u w=0.6u m=1
M12 GND N_17 S GND mn5  l=0.5u w=0.98u m=1
M13 N_17 CI N_5 GND mn5  l=0.5u w=0.6u m=1
M14 N_10 N_8 N_17 GND mn5  l=0.5u w=0.6u m=1
M15 CO N_9 VDD VDD mp5  l=0.42u w=1.28u m=1
M16 N_8 CI VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_9 N_10 N_8 VDD mp5  l=0.42u w=0.62u m=1
M18 N_9 N_5 N_7 VDD mp5  l=0.42u w=0.62u m=1
M19 N_7 N_6 N_5 VDD mp5  l=0.42u w=0.62u m=1
M20 N_6 N_7 N_5 VDD mp5  l=0.42u w=0.62u m=1
M21 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_6 N_14 N_10 VDD mp5  l=0.42u w=0.62u m=1
M23 N_14 N_6 N_10 VDD mp5  l=0.42u w=0.62u m=1
M24 N_14 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_7 B VDD VDD mp5  l=0.42u w=0.62u m=1
M26 VDD N_17 S VDD mp5  l=0.42u w=1.28u m=1
M27 N_10 CI N_17 VDD mp5  l=0.42u w=0.62u m=1
M28 N_5 N_8 N_17 VDD mp5  l=0.42u w=0.62u m=1
.ends ad01d2
* SPICE INPUT		Mon Sep 24 12:03:31 2018	ah01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d0
.subckt ah01d0 B A GND S CO VDD
M1 N_26 B GND GND mn5  l=0.5u w=0.6u m=1
M2 N_26 A N_7 GND mn5  l=0.5u w=0.6u m=1
M3 CO N_7 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_2 B GND GND mn5  l=0.5u w=0.6u m=1
M5 N_4 A GND GND mn5  l=0.5u w=0.6u m=1
M6 N_12 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_4 B S GND mn5  l=0.5u w=0.6u m=1
M8 S N_2 N_12 GND mn5  l=0.5u w=0.6u m=1
M9 N_2 B VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_4 A VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_4 N_2 S VDD mp5  l=0.42u w=0.62u m=1
M12 N_12 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 S B N_12 VDD mp5  l=0.42u w=0.62u m=1
M14 N_7 B VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_7 A VDD VDD mp5  l=0.42u w=0.62u m=1
M16 CO N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends ah01d0
* SPICE INPUT		Mon Sep 24 12:03:40 2018	ah01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d1
.subckt ah01d1 A B CO GND VDD S
M1 S N_9 N_14 GND mn5  l=0.5u w=0.72u m=1
M2 S B N_7 GND mn5  l=0.5u w=0.72u m=1
M3 N_14 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_9 B GND GND mn5  l=0.5u w=0.6u m=1
M5 N_7 A GND GND mn5  l=0.5u w=0.6u m=1
M6 N_16 B GND GND mn5  l=0.5u w=0.6u m=1
M7 CO N_3 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_16 A N_3 GND mn5  l=0.5u w=0.6u m=1
M9 N_14 B S VDD mp5  l=0.42u w=0.96u m=1
M10 N_7 N_9 S VDD mp5  l=0.42u w=0.96u m=1
M11 N_14 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_9 B VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_7 A VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_3 B VDD VDD mp5  l=0.42u w=0.62u m=1
M15 CO N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_3 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends ah01d1
* SPICE INPUT		Mon Sep 24 12:03:49 2018	ah01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d2
.subckt ah01d2 A B GND VDD CO S
M1 CO N_8 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_25 A N_8 GND mn5  l=0.5u w=0.6u m=1
M3 N_25 B GND GND mn5  l=0.5u w=0.6u m=1
M4 N_4 B GND GND mn5  l=0.5u w=0.6u m=1
M5 N_14 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M6 S N_4 N_14 GND mn5  l=0.5u w=0.98u m=1
M7 S B N_5 GND mn5  l=0.5u w=0.98u m=1
M8 N_5 A GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 B VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_14 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 S B N_14 VDD mp5  l=0.42u w=1.28u m=1
M12 S N_4 N_5 VDD mp5  l=0.42u w=1.28u m=1
M13 CO N_8 VDD VDD mp5  l=0.42u w=1.28u m=1
M14 N_8 A VDD VDD mp5  l=0.42u w=0.62u m=1
M15 VDD A N_5 VDD mp5  l=0.42u w=0.62u m=1
M16 N_8 B VDD VDD mp5  l=0.42u w=0.62u m=1
.ends ah01d2
* SPICE INPUT		Mon Sep 24 12:03:58 2018	an02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d0
.subckt an02d0 A B GND Y VDD
M1 Y N_4 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_12 B GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 A N_4 GND mn5  l=0.5u w=0.6u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M5 N_4 B VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an02d0
* SPICE INPUT		Mon Sep 24 12:04:07 2018	an02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d1
.subckt an02d1 A B GND Y VDD
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.6u m=1
M3 N_8 A N_4 GND mn5  l=0.5u w=0.6u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M5 N_4 B VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an02d1
* SPICE INPUT		Mon Sep 24 12:04:15 2018	an02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d2
.subckt an02d2 A B GND Y VDD
M1 Y N_4 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_8 B GND GND mn5  l=0.5u w=0.6u m=1
M3 N_8 A N_4 GND mn5  l=0.5u w=0.6u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
M5 N_4 B VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_4 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an02d2
* SPICE INPUT		Mon Sep 24 12:04:24 2018	an03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d0
.subckt an03d0 C A B VDD GND Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.6u m=1
M3 N_9 A N_5 GND mn5  l=0.5u w=0.6u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_5 B VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_5 A VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 C VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an03d0
* SPICE INPUT		Mon Sep 24 12:04:32 2018	an03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d1
.subckt an03d1 C A B VDD GND Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.6u m=1
M3 N_9 A N_5 GND mn5  l=0.5u w=0.6u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_5 B VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_5 A VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 C VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an03d1
* SPICE INPUT		Mon Sep 24 12:04:41 2018	an03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d2
.subckt an03d2 C A B VDD GND Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_10 B N_9 GND mn5  l=0.5u w=0.6u m=1
M3 N_9 A N_5 GND mn5  l=0.5u w=0.6u m=1
M4 N_10 C GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M6 N_5 B VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_5 A VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 C VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an03d2
* SPICE INPUT		Mon Sep 24 12:04:50 2018	an04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d0
.subckt an04d0 A B C D VDD Y GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_12 D GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 C N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A N_6 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_6 D VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 C VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an04d0
* SPICE INPUT		Mon Sep 24 12:04:58 2018	an04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d1
.subckt an04d1 A B C D VDD Y GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_12 D GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 C N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A N_6 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_6 D VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 C VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an04d1
* SPICE INPUT		Mon Sep 24 12:05:07 2018	an04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d2
.subckt an04d2 A B C D VDD Y GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_12 D GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 C N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A N_6 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_6 D VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 C VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 B VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an04d2
* SPICE INPUT		Mon Sep 24 12:05:15 2018	an12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an12d0
.subckt an12d0 B AN VDD GND Y
M1 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_15 B GND GND mn5  l=0.5u w=0.6u m=1
M4 N_15 N_2 N_4 GND mn5  l=0.5u w=0.6u m=1
M5 N_2 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_4 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an12d0
* SPICE INPUT		Mon Sep 24 12:05:24 2018	an12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an12d1
.subckt an12d1 AN B VDD GND Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_15 B GND GND mn5  l=0.5u w=0.6u m=1
M3 N_15 N_3 N_5 GND mn5  l=0.5u w=0.6u m=1
M4 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M6 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_5 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an12d1
* SPICE INPUT		Mon Sep 24 12:05:32 2018	an12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an12d2
.subckt an12d2 AN B VDD GND Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_15 B GND GND mn5  l=0.5u w=0.6u m=1
M3 N_15 N_3 N_5 GND mn5  l=0.5u w=0.6u m=1
M4 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M6 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_5 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an12d2
* SPICE INPUT		Mon Sep 24 12:05:42 2018	an13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an13d0
.subckt an13d0 B C AN Y GND VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 GND C N_10 GND mn5  l=0.5u w=0.6u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_11 N_2 N_6 GND mn5  l=0.5u w=0.6u m=1
M6 N_6 C VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_6 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_2 AN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an13d0
* SPICE INPUT		Mon Sep 24 12:05:50 2018	an13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an13d1
.subckt an13d1 AN B C Y GND VDD
M1 GND C N_16 GND mn5  l=0.5u w=0.6u m=1
M2 N_17 B N_16 GND mn5  l=0.5u w=0.6u m=1
M3 N_17 N_4 N_3 GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_4 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_3 C VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_4 AN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an13d1
* SPICE INPUT		Mon Sep 24 12:05:59 2018	an13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an13d2
.subckt an13d2 B C AN VDD GND Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_10 C GND GND mn5  l=0.5u w=0.6u m=1
M4 N_11 B N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_6 N_2 N_11 GND mn5  l=0.5u w=0.6u m=1
M6 N_6 C VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_6 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M10 N_2 AN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an13d2
* SPICE INPUT		Mon Sep 24 12:06:07 2018	an23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an23d0
.subckt an23d0 C AN BN Y VDD GND
M1 N_5 BN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 N_5 N_11 GND mn5  l=0.5u w=0.6u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_11 N_3 N_4 GND mn5  l=0.5u w=0.6u m=1
M6 N_12 C GND GND mn5  l=0.5u w=0.6u m=1
M7 N_5 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_4 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_4 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_4 C VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an23d0
* SPICE INPUT		Mon Sep 24 12:06:16 2018	an23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an23d1
.subckt an23d1 BN AN C GND VDD Y
M1 N_11 N_7 N_4 GND mn5  l=0.5u w=0.6u m=1
M2 N_12 N_6 N_11 GND mn5  l=0.5u w=0.6u m=1
M3 N_12 C GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_7 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_6 BN GND GND mn5  l=0.5u w=0.6u m=1
M7 N_4 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_4 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_4 C VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 N_7 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_6 BN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an23d1
* SPICE INPUT		Mon Sep 24 12:06:24 2018	an23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an23d2
.subckt an23d2 C AN BN Y VDD GND
M1 N_5 BN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 N_5 N_11 GND mn5  l=0.5u w=0.6u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.98u m=1
M5 N_11 N_3 N_4 GND mn5  l=0.5u w=0.6u m=1
M6 N_12 C GND GND mn5  l=0.5u w=0.6u m=1
M7 N_5 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_4 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
M11 N_4 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_4 C VDD VDD mp5  l=0.42u w=0.62u m=1
.ends an23d2
* SPICE INPUT		Mon Sep 24 14:01:53 2018	antenna
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=antenna
.subckt antenna GND VDD A
D1 A VDD dppnw_5  area=0.5375p pj=3.36u
D2 GND A dnppw_5  area=0.4386p pj=2.9u
.ends antenna
* SPICE INPUT		Mon Sep 24 12:06:38 2018	aoi211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d0
.subckt aoi211d0 C0 A1 A0 B0 VDD Y GND
M1 Y B0 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_16 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 Y A1 N_16 GND mn5  l=0.5u w=0.6u m=1
M4 Y C0 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_8 B0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M6 N_8 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_8 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y C0 N_10 VDD mp5  l=0.42u w=0.62u m=1
.ends aoi211d0
* SPICE INPUT		Mon Sep 24 12:06:47 2018	aoi211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d1
.subckt aoi211d1 C0 A1 A0 B0 VDD Y GND
M1 Y B0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_16 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y A1 N_16 GND mn5  l=0.5u w=0.72u m=1
M4 Y C0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_8 B0 N_10 VDD mp5  l=0.42u w=0.96u m=1
M6 VDD A0 N_8 VDD mp5  l=0.42u w=0.96u m=1
M7 N_8 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y C0 N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends aoi211d1
* SPICE INPUT		Mon Sep 24 12:06:55 2018	aoi211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d2
.subckt aoi211d2 A1 B0 C0 A0 Y VDD GND
M1 N_16 A0 GND GND mn5  l=0.5u w=0.98u m=1
M2 Y C0 GND GND mn5  l=0.5u w=0.98u m=1
M3 Y B0 GND GND mn5  l=0.5u w=0.98u m=1
M4 Y A1 N_16 GND mn5  l=0.5u w=0.98u m=1
M5 VDD A0 N_8 VDD mp5  l=0.42u w=1.28u m=1
M6 Y C0 N_10 VDD mp5  l=0.42u w=1.28u m=1
M7 N_8 B0 N_10 VDD mp5  l=0.42u w=1.28u m=1
M8 N_8 A1 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends aoi211d2
* SPICE INPUT		Mon Sep 24 12:07:03 2018	aoi21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d0
.subckt aoi21d0 A0 A1 B0 VDD GND Y
M1 GND B0 Y GND mn5  l=0.5u w=0.6u m=1
M2 N_13 A1 Y GND mn5  l=0.5u w=0.6u m=1
M3 N_13 A0 GND GND mn5  l=0.5u w=0.6u m=1
M4 Y B0 N_8 VDD mp5  l=0.42u w=0.62u m=1
M5 VDD A1 N_8 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD A0 N_8 VDD mp5  l=0.42u w=0.62u m=1
.ends aoi21d0
* SPICE INPUT		Mon Sep 24 12:07:12 2018	aoi21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d1
.subckt aoi21d1 A0 A1 B0 VDD GND Y
M1 GND B0 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_13 A1 Y GND mn5  l=0.5u w=0.72u m=1
M3 N_13 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 N_8 VDD mp5  l=0.42u w=0.96u m=1
M5 VDD A1 N_8 VDD mp5  l=0.42u w=0.96u m=1
M6 VDD A0 N_8 VDD mp5  l=0.42u w=0.96u m=1
.ends aoi21d1
* SPICE INPUT		Mon Sep 24 12:07:20 2018	aoi21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d2
.subckt aoi21d2 A0 A1 B0 GND Y VDD
M1 GND B0 Y GND mn5  l=0.5u w=0.96u m=1
M2 N_13 A1 Y GND mn5  l=0.5u w=0.96u m=1
M3 N_13 A0 GND GND mn5  l=0.5u w=0.96u m=1
M4 Y B0 N_6 VDD mp5  l=0.42u w=1.28u m=1
M5 VDD A1 N_6 VDD mp5  l=0.42u w=1.28u m=1
M6 VDD A0 N_6 VDD mp5  l=0.42u w=1.28u m=1
.ends aoi21d2
* SPICE INPUT		Mon Sep 24 12:07:29 2018	aoi221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d0
.subckt aoi221d0 A0 B1 A1 B0 C0 Y GND VDD
M1 Y C0 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_12 B0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_13 A1 Y GND mn5  l=0.5u w=0.6u m=1
M4 Y B1 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_13 A0 GND GND mn5  l=0.5u w=0.6u m=1
M6 Y C0 N_7 VDD mp5  l=0.42u w=0.62u m=1
M7 N_9 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_9 A1 N_7 VDD mp5  l=0.42u w=0.62u m=1
M9 N_9 B1 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_7 A0 N_9 VDD mp5  l=0.42u w=0.62u m=1
.ends aoi221d0
* SPICE INPUT		Mon Sep 24 12:07:38 2018	aoi221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d1
.subckt aoi221d1 B0 B1 A1 A0 C0 Y VDD GND
M1 Y C0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_13 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_13 A1 Y GND mn5  l=0.5u w=0.72u m=1
M4 Y B1 N_12 GND mn5  l=0.5u w=0.72u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y C0 N_8 VDD mp5  l=0.42u w=0.96u m=1
M7 N_7 A0 N_8 VDD mp5  l=0.42u w=0.96u m=1
M8 N_7 A1 N_8 VDD mp5  l=0.42u w=0.96u m=1
M9 N_7 B1 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 VDD B0 N_7 VDD mp5  l=0.42u w=0.96u m=1
.ends aoi221d1
* SPICE INPUT		Mon Sep 24 12:07:46 2018	aoi221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d2
.subckt aoi221d2 A1 B1 B0 C0 A0 GND VDD Y
M1 N_13 A0 GND GND mn5  l=0.5u w=0.98u m=1
M2 Y C0 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_12 B0 GND GND mn5  l=0.5u w=0.98u m=1
M4 Y B1 N_12 GND mn5  l=0.5u w=0.98u m=1
M5 N_13 A1 Y GND mn5  l=0.5u w=0.98u m=1
M6 N_9 A0 N_11 VDD mp5  l=0.42u w=1.28u m=1
M7 VDD B0 N_9 VDD mp5  l=0.42u w=1.28u m=1
M8 N_9 B1 VDD VDD mp5  l=0.42u w=1.28u m=1
M9 N_9 A1 N_11 VDD mp5  l=0.42u w=1.28u m=1
M10 Y C0 N_11 VDD mp5  l=0.42u w=1.28u m=1
.ends aoi221d2
* SPICE INPUT		Mon Sep 24 12:07:55 2018	aoi22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d0
.subckt aoi22d0 B0 B1 A1 A0 GND VDD Y
M1 N_15 A0 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y A1 N_15 GND mn5  l=0.5u w=0.6u m=1
M3 Y B1 N_14 GND mn5  l=0.5u w=0.6u m=1
M4 GND B0 N_14 GND mn5  l=0.5u w=0.6u m=1
M5 N_8 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_8 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_8 B1 Y VDD mp5  l=0.42u w=0.62u m=1
M8 N_8 B0 Y VDD mp5  l=0.42u w=0.62u m=1
.ends aoi22d0
* SPICE INPUT		Mon Sep 24 12:08:03 2018	aoi22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d1
.subckt aoi22d1 B0 B1 A1 A0 GND VDD Y
M1 N_11 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A1 N_11 GND mn5  l=0.5u w=0.72u m=1
M3 Y B1 N_10 GND mn5  l=0.5u w=0.72u m=1
M4 GND B0 N_10 GND mn5  l=0.5u w=0.72u m=1
M5 VDD A0 N_8 VDD mp5  l=0.42u w=0.96u m=1
M6 N_8 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_8 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M8 N_8 B0 Y VDD mp5  l=0.42u w=0.96u m=1
.ends aoi22d1
* SPICE INPUT		Mon Sep 24 12:08:12 2018	aoi22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d2
.subckt aoi22d2 B0 B1 A1 A0 GND VDD Y
M1 N_11 A0 GND GND mn5  l=0.5u w=0.98u m=1
M2 Y A1 N_11 GND mn5  l=0.5u w=0.98u m=1
M3 Y B1 N_10 GND mn5  l=0.5u w=0.98u m=1
M4 GND B0 N_10 GND mn5  l=0.5u w=0.98u m=1
M5 VDD A0 N_7 VDD mp5  l=0.42u w=1.28u m=1
M6 N_7 A1 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_7 B1 Y VDD mp5  l=0.42u w=1.28u m=1
M8 N_7 B0 Y VDD mp5  l=0.42u w=1.28u m=1
.ends aoi22d2
* SPICE INPUT		Mon Sep 24 12:08:21 2018	aoi31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d0
.subckt aoi31d0 B0 A2 A0 A1 Y VDD GND
M1 N_11 A1 N_10 GND mn5  l=0.5u w=0.6u m=1
M2 N_10 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_11 A2 Y GND mn5  l=0.5u w=0.6u m=1
M4 GND B0 Y GND mn5  l=0.5u w=0.6u m=1
M5 VDD A1 N_9 VDD mp5  l=0.42u w=0.62u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 VDD A2 N_9 VDD mp5  l=0.42u w=0.62u m=1
M8 Y B0 N_9 VDD mp5  l=0.42u w=0.62u m=1
.ends aoi31d0
* SPICE INPUT		Mon Sep 24 12:08:30 2018	aoi31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d1
.subckt aoi31d1 B0 A2 A0 A1 Y VDD GND
M1 N_11 A1 N_10 GND mn5  l=0.5u w=0.72u m=1
M2 N_10 A0 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 A2 Y GND mn5  l=0.5u w=0.72u m=1
M4 GND B0 Y GND mn5  l=0.5u w=0.72u m=1
M5 VDD A1 N_9 VDD mp5  l=0.42u w=0.96u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 VDD A2 N_9 VDD mp5  l=0.42u w=0.96u m=1
M8 Y B0 N_9 VDD mp5  l=0.42u w=0.96u m=1
.ends aoi31d1
* SPICE INPUT		Mon Sep 24 12:08:39 2018	aoi31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d2
.subckt aoi31d2 B0 A2 A1 A0 Y GND VDD
M1 N_10 A0 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_11 A1 N_10 GND mn5  l=0.5u w=0.98u m=1
M3 N_11 A2 Y GND mn5  l=0.5u w=0.98u m=1
M4 GND B0 Y GND mn5  l=0.5u w=0.98u m=1
M5 N_6 A0 VDD VDD mp5  l=0.42u w=1.28u m=1
M6 VDD A1 N_6 VDD mp5  l=0.42u w=1.28u m=1
M7 VDD A2 N_6 VDD mp5  l=0.42u w=1.28u m=1
M8 Y B0 N_6 VDD mp5  l=0.42u w=1.28u m=1
.ends aoi31d2
* SPICE INPUT		Mon Sep 24 12:08:47 2018	aoi32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d0
.subckt aoi32d0 B0 B1 A2 A0 A1 Y GND VDD
M1 N_13 A1 N_12 GND mn5  l=0.5u w=0.6u m=1
M2 N_12 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 Y A2 N_13 GND mn5  l=0.5u w=0.6u m=1
M4 Y B1 N_11 GND mn5  l=0.5u w=0.6u m=1
M5 GND B0 N_11 GND mn5  l=0.5u w=0.6u m=1
M6 N_7 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_7 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_7 A2 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_7 B1 Y VDD mp5  l=0.42u w=0.62u m=1
M10 N_7 B0 Y VDD mp5  l=0.42u w=0.62u m=1
.ends aoi32d0
* SPICE INPUT		Mon Sep 24 12:08:56 2018	aoi32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d1
.subckt aoi32d1 B0 B1 A2 A1 A0 VDD GND Y
M1 N_12 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_13 A1 N_12 GND mn5  l=0.5u w=0.72u m=1
M3 Y A2 N_13 GND mn5  l=0.5u w=0.72u m=1
M4 Y B1 N_11 GND mn5  l=0.5u w=0.72u m=1
M5 GND B0 N_11 GND mn5  l=0.5u w=0.72u m=1
M6 N_7 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_7 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_7 A2 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_7 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M10 N_7 B0 Y VDD mp5  l=0.42u w=0.96u m=1
.ends aoi32d1
* SPICE INPUT		Mon Sep 24 12:09:05 2018	aoi32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d2
.subckt aoi32d2 GND Y VDD A1 B1 B0 A2 A0
M1 GND B0 N_6 GND mn5  l=0.5u w=0.98u m=1
M2 Y B1 N_6 GND mn5  l=0.5u w=0.98u m=1
M3 Y A2 N_8 GND mn5  l=0.5u w=0.98u m=1
M4 N_8 A1 N_7 GND mn5  l=0.5u w=0.98u m=1
M5 N_7 A0 GND GND mn5  l=0.5u w=0.98u m=1
M6 N_12 B0 Y VDD mp5  l=0.42u w=1.28u m=1
M7 N_12 B1 Y VDD mp5  l=0.42u w=1.28u m=1
M8 N_12 A2 VDD VDD mp5  l=0.42u w=1.28u m=1
M9 VDD A1 N_12 VDD mp5  l=0.42u w=1.28u m=1
M10 N_12 A0 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends aoi32d2
* SPICE INPUT		Mon Sep 24 12:09:14 2018	aoi33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d0
.subckt aoi33d0 A0 B0 B1 B2 A2 A1 VDD GND Y
M1 N_14 A1 N_13 GND mn5  l=0.5u w=0.6u m=1
M2 Y A2 N_14 GND mn5  l=0.5u w=0.6u m=1
M3 N_15 B2 Y GND mn5  l=0.5u w=0.6u m=1
M4 N_15 B1 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 GND B0 N_12 GND mn5  l=0.5u w=0.6u m=1
M6 N_13 A0 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_10 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_10 A2 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y B2 N_10 VDD mp5  l=0.42u w=0.62u m=1
M10 Y B1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M11 Y B0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M12 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends aoi33d0
* SPICE INPUT		Mon Sep 24 12:09:22 2018	aoi33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d1
.subckt aoi33d1 B0 B1 B2 A2 A1 A0 Y VDD GND
M1 N_13 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_14 A1 N_13 GND mn5  l=0.5u w=0.72u m=1
M3 Y A2 N_14 GND mn5  l=0.5u w=0.72u m=1
M4 N_15 B2 Y GND mn5  l=0.5u w=0.72u m=1
M5 N_15 B1 N_12 GND mn5  l=0.5u w=0.72u m=1
M6 GND B0 N_12 GND mn5  l=0.5u w=0.72u m=1
M7 N_11 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_11 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_11 A2 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y B2 N_11 VDD mp5  l=0.42u w=0.96u m=1
M11 Y B1 N_11 VDD mp5  l=0.42u w=0.96u m=1
M12 Y B0 N_11 VDD mp5  l=0.42u w=0.96u m=1
.ends aoi33d1
* SPICE INPUT		Mon Sep 24 12:09:31 2018	aoi33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d2
.subckt aoi33d2 GND Y VDD A1 B2 B1 A2 B0 A0
M1 GND B0 N_6 GND mn5  l=0.5u w=0.98u m=1
M2 N_9 B1 N_6 GND mn5  l=0.5u w=0.98u m=1
M3 N_9 B2 Y GND mn5  l=0.5u w=0.98u m=1
M4 Y A2 N_8 GND mn5  l=0.5u w=0.98u m=1
M5 N_8 A1 N_7 GND mn5  l=0.5u w=0.98u m=1
M6 N_7 A0 GND GND mn5  l=0.5u w=0.98u m=1
M7 Y B0 N_13 VDD mp5  l=0.42u w=1.28u m=1
M8 Y B1 N_13 VDD mp5  l=0.42u w=1.28u m=1
M9 Y B2 N_13 VDD mp5  l=0.42u w=1.28u m=1
M10 N_13 A2 VDD VDD mp5  l=0.42u w=1.28u m=1
M11 VDD A1 N_13 VDD mp5  l=0.42u w=1.28u m=1
M12 N_13 A0 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends aoi33d2
* SPICE INPUT		Mon Sep 24 12:09:41 2018	aoim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d0
.subckt aoim21d0 A0N A1N B0 GND Y VDD
M1 GND N_5 Y GND mn5  l=0.5u w=0.6u m=1
M2 Y B0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 A1N GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 A0N GND GND mn5  l=0.5u w=0.6u m=1
M5 VDD N_5 N_9 VDD mp5  l=0.42u w=0.62u m=1
M6 Y B0 N_9 VDD mp5  l=0.42u w=0.62u m=1
M7 N_5 A1N N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 VDD A0N N_10 VDD mp5  l=0.42u w=0.62u m=1
.ends aoim21d0
* SPICE INPUT		Mon Sep 24 12:09:50 2018	aoim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d1
.subckt aoim21d1 A1N A0N B0 GND VDD Y
M1 GND B0 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_2 A0N GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 A1N GND GND mn5  l=0.5u w=0.6u m=1
M4 GND N_2 Y GND mn5  l=0.5u w=0.72u m=1
M5 VDD A0N N_9 VDD mp5  l=0.42u w=0.62u m=1
M6 N_2 A1N N_9 VDD mp5  l=0.42u w=0.62u m=1
M7 Y B0 N_10 VDD mp5  l=0.42u w=0.96u m=1
M8 VDD N_2 N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends aoim21d1
* SPICE INPUT		Mon Sep 24 12:09:58 2018	aoim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d2
.subckt aoim21d2 B0 A0N A1N GND VDD Y
M1 N_4 A1N GND GND mn5  l=0.5u w=0.6u m=1
M2 GND N_4 Y GND mn5  l=0.5u w=0.98u m=1
M3 N_4 A0N GND GND mn5  l=0.5u w=0.6u m=1
M4 GND B0 Y GND mn5  l=0.5u w=0.98u m=1
M5 N_4 A1N N_9 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD A0N N_9 VDD mp5  l=0.42u w=0.62u m=1
M7 VDD N_4 N_10 VDD mp5  l=0.42u w=1.28u m=1
M8 Y B0 N_10 VDD mp5  l=0.42u w=1.28u m=1
.ends aoim21d2
* SPICE INPUT		Mon Sep 24 12:10:07 2018	aoim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d0
.subckt aoim22d0 B0 A1N B1 A0N Y GND VDD
M1 GND N_6 Y GND mn5  l=0.5u w=0.6u m=1
M2 N_6 A0N GND GND mn5  l=0.5u w=0.6u m=1
M3 N_18 B1 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 A1N GND GND mn5  l=0.5u w=0.6u m=1
M5 N_18 B0 Y GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 N_9 VDD mp5  l=0.42u w=0.62u m=1
M7 VDD B1 N_9 VDD mp5  l=0.42u w=0.62u m=1
M8 VDD B0 N_9 VDD mp5  l=0.42u w=0.62u m=1
M9 VDD A0N N_11 VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 A1N N_11 VDD mp5  l=0.42u w=0.62u m=1
.ends aoim22d0
* SPICE INPUT		Mon Sep 24 12:10:16 2018	aoim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d1
.subckt aoim22d1 B0 A1N B1 A0N Y GND VDD
M1 GND N_6 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_6 A0N GND GND mn5  l=0.5u w=0.6u m=1
M3 N_18 B1 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_6 A1N GND GND mn5  l=0.5u w=0.6u m=1
M5 N_18 B0 Y GND mn5  l=0.5u w=0.72u m=1
M6 Y N_6 N_9 VDD mp5  l=0.42u w=0.96u m=1
M7 VDD B1 N_9 VDD mp5  l=0.42u w=0.96u m=1
M8 VDD B0 N_9 VDD mp5  l=0.42u w=0.96u m=1
M9 VDD A0N N_11 VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 A1N N_11 VDD mp5  l=0.42u w=0.62u m=1
.ends aoim22d1
* SPICE INPUT		Mon Sep 24 12:10:25 2018	aoim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d2
.subckt aoim22d2 B0 B1 A1N A0N GND VDD Y
M1 N_2 A0N GND GND mn5  l=0.5u w=0.6u m=1
M2 N_2 A1N GND GND mn5  l=0.5u w=0.6u m=1
M3 N_11 B1 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_11 B0 Y GND mn5  l=0.5u w=0.98u m=1
M5 GND N_2 Y GND mn5  l=0.5u w=0.98u m=1
M6 VDD B1 N_10 VDD mp5  l=0.42u w=1.28u m=1
M7 VDD B0 N_10 VDD mp5  l=0.42u w=1.28u m=1
M8 Y N_2 N_10 VDD mp5  l=0.42u w=1.28u m=1
M9 VDD A0N N_19 VDD mp5  l=0.42u w=0.62u m=1
M10 N_2 A1N N_19 VDD mp5  l=0.42u w=0.62u m=1
.ends aoim22d2
* SPICE INPUT		Mon Sep 24 12:10:33 2018	aoim31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim31d0
.subckt aoim31d0 A0N A1N A2N B0 Y VDD GND
M1 GND B0 Y GND mn5  l=0.5u w=0.6u m=1
M2 GND N_5 Y GND mn5  l=0.5u w=0.6u m=1
M3 N_5 A2N GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 A1N GND GND mn5  l=0.5u w=0.6u m=1
M5 N_5 A0N GND GND mn5  l=0.5u w=0.6u m=1
M6 Y B0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 VDD N_5 N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 A2N N_5 VDD mp5  l=0.42u w=0.62u m=1
M9 N_12 A1N N_11 VDD mp5  l=0.42u w=0.62u m=1
M10 N_12 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
.ends aoim31d0
* SPICE INPUT		Mon Sep 24 12:10:42 2018	aoim31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim31d1
.subckt aoim31d1 B0 A0N A1N A2N Y VDD GND
M1 GND N_6 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_6 A2N GND GND mn5  l=0.5u w=0.6u m=1
M3 N_6 A1N GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 A0N GND GND mn5  l=0.5u w=0.6u m=1
M5 GND B0 Y GND mn5  l=0.5u w=0.72u m=1
M6 N_10 A2N N_6 VDD mp5  l=0.42u w=0.62u m=1
M7 N_11 A1N N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M9 VDD N_6 N_12 VDD mp5  l=0.42u w=0.96u m=1
M10 Y B0 N_12 VDD mp5  l=0.42u w=0.96u m=1
.ends aoim31d1
* SPICE INPUT		Mon Sep 24 12:10:50 2018	aoim31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim31d2
.subckt aoim31d2 B0 A0N A1N A2N Y VDD GND
M1 GND N_6 Y GND mn5  l=0.5u w=0.98u m=1
M2 N_6 A2N GND GND mn5  l=0.5u w=0.6u m=1
M3 N_6 A1N GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 A0N GND GND mn5  l=0.5u w=0.6u m=1
M5 GND B0 Y GND mn5  l=0.5u w=0.98u m=1
M6 N_10 A2N N_6 VDD mp5  l=0.42u w=0.62u m=1
M7 N_11 A1N N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M9 VDD N_6 N_12 VDD mp5  l=0.42u w=1.28u m=1
M10 Y B0 N_12 VDD mp5  l=0.42u w=1.28u m=1
.ends aoim31d2
* SPICE INPUT		Mon Sep 24 12:11:00 2018	aor211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d0
.subckt aor211d0 C0 B0 A0 A1 VDD GND Y
M1 N_18 A1 N_2 GND mn5  l=0.5u w=0.6u m=1
M2 N_18 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_2 C0 GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.6u m=1
M6 VDD A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_10 B0 N_11 VDD mp5  l=0.42u w=0.62u m=1
M9 N_11 C0 N_2 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends aor211d0
* SPICE INPUT		Mon Sep 24 12:11:08 2018	aor211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d1
.subckt aor211d1 C0 B0 A0 A1 VDD GND Y
M1 N_11 A1 N_2 GND mn5  l=0.5u w=0.6u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_2 C0 GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 VDD A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_10 B0 N_19 VDD mp5  l=0.42u w=0.62u m=1
M9 N_19 C0 N_2 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aor211d1
* SPICE INPUT		Mon Sep 24 12:11:17 2018	aor211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d2
.subckt aor211d2 C0 B0 A0 A1 GND VDD Y
M1 N_11 A1 N_2 GND mn5  l=0.5u w=0.6u m=1
M2 N_11 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 B0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_2 C0 GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.98u m=1
M6 VDD A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_10 B0 N_19 VDD mp5  l=0.42u w=0.62u m=1
M9 N_19 C0 N_2 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends aor211d2
* SPICE INPUT		Mon Sep 24 12:11:25 2018	aor21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d0
.subckt aor21d0 A1 A0 B0 GND VDD Y
M1 N_4 B0 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_10 A0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_4 A1 N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_6 B0 N_4 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD A0 N_6 VDD mp5  l=0.42u w=0.62u m=1
M7 VDD A1 N_6 VDD mp5  l=0.42u w=0.62u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends aor21d0
* SPICE INPUT		Mon Sep 24 12:11:34 2018	aor21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d1
.subckt aor21d1 A1 A0 B0 GND VDD Y
M1 N_4 B0 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_10 A0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_4 A1 N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_6 B0 N_4 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD A0 N_6 VDD mp5  l=0.42u w=0.62u m=1
M7 VDD A1 N_6 VDD mp5  l=0.42u w=0.62u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aor21d1
* SPICE INPUT		Mon Sep 24 12:11:43 2018	aor21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d2
.subckt aor21d2 A1 A0 B0 GND VDD Y
M1 N_4 B0 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_10 A0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_4 A1 N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_6 B0 N_4 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD A0 N_6 VDD mp5  l=0.42u w=0.62u m=1
M7 VDD A1 N_6 VDD mp5  l=0.42u w=0.62u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends aor21d2
* SPICE INPUT		Mon Sep 24 12:11:52 2018	aor221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d0
.subckt aor221d0 B1 B0 C0 A0 A1 GND Y VDD
M1 N_14 A1 N_2 GND mn5  l=0.5u w=0.6u m=1
M2 N_14 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 C0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 B0 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 B1 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 GND N_2 Y GND mn5  l=0.5u w=0.6u m=1
M7 N_9 A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_9 A0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M9 N_2 C0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M10 VDD B0 N_9 VDD mp5  l=0.42u w=0.62u m=1
M11 N_9 B1 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 VDD N_2 Y VDD mp5  l=0.42u w=0.62u m=1
.ends aor221d0
* SPICE INPUT		Mon Sep 24 12:12:00 2018	aor221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d1
.subckt aor221d1 B1 B0 C0 A0 A1 GND Y VDD
M1 N_14 A1 N_2 GND mn5  l=0.5u w=0.6u m=1
M2 N_14 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 C0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 B0 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 B1 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_9 A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_9 A0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M9 N_2 C0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M10 VDD B0 N_9 VDD mp5  l=0.42u w=0.62u m=1
M11 N_9 B1 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aor221d1
* SPICE INPUT		Mon Sep 24 12:12:09 2018	aor221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d2
.subckt aor221d2 B1 B0 C0 A0 A1 GND Y VDD
M1 N_14 A1 N_2 GND mn5  l=0.5u w=0.6u m=1
M2 N_14 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 C0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 B0 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 B1 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.98u m=1
M7 N_9 A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_9 A0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M9 N_2 C0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M10 VDD B0 N_9 VDD mp5  l=0.42u w=0.62u m=1
M11 N_9 B1 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends aor221d2
* SPICE INPUT		Mon Sep 24 12:12:17 2018	aor22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d0
.subckt aor22d0 B0 B1 A1 A0 Y VDD GND
M1 N_11 A0 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 A1 N_11 GND mn5  l=0.5u w=0.6u m=1
M3 N_12 B1 N_3 GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.6u m=1
M6 VDD A0 N_9 VDD mp5  l=0.42u w=0.62u m=1
M7 N_9 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_9 B1 N_3 VDD mp5  l=0.42u w=0.62u m=1
M9 N_3 B0 N_9 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends aor22d0
* SPICE INPUT		Mon Sep 24 12:12:26 2018	aor22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d1
.subckt aor22d1 B0 B1 A1 A0 Y VDD GND
M1 N_11 A0 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 A1 N_11 GND mn5  l=0.5u w=0.6u m=1
M3 N_12 B1 N_3 GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.6u m=1
M6 VDD A0 N_9 VDD mp5  l=0.42u w=0.62u m=1
M7 N_9 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_9 B1 N_3 VDD mp5  l=0.42u w=0.62u m=1
M9 N_3 B0 N_9 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aor22d1
* SPICE INPUT		Mon Sep 24 12:12:35 2018	aor22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d2
.subckt aor22d2 B0 B1 A1 A0 GND VDD Y
M1 N_11 A0 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 A1 N_11 GND mn5  l=0.5u w=0.6u m=1
M3 N_12 B1 N_3 GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.98u m=1
M5 N_12 B0 GND GND mn5  l=0.5u w=0.6u m=1
M6 VDD A0 N_8 VDD mp5  l=0.42u w=0.62u m=1
M7 N_8 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_8 B1 N_3 VDD mp5  l=0.42u w=0.62u m=1
M9 N_3 B0 N_8 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends aor22d2
* SPICE INPUT		Mon Sep 24 12:12:43 2018	aor311d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor311d0
.subckt aor311d0 B0 C0 A0 A2 A1 GND VDD Y
M1 N_6 A1 N_20 GND mn5  l=0.5u w=0.6u m=1
M2 GND N_6 Y GND mn5  l=0.5u w=0.6u m=1
M3 N_19 A2 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_20 A0 N_19 GND mn5  l=0.5u w=0.6u m=1
M5 N_6 C0 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_6 B0 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_8 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 VDD N_6 Y VDD mp5  l=0.42u w=0.62u m=1
M9 N_8 A2 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_8 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_6 C0 N_12 VDD mp5  l=0.42u w=0.62u m=1
M12 N_8 B0 N_12 VDD mp5  l=0.42u w=0.62u m=1
.ends aor311d0
* SPICE INPUT		Mon Sep 24 12:12:52 2018	aor311d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor311d1
.subckt aor311d1 C0 B0 A1 A0 A2 VDD Y GND
M1 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_19 A2 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_20 A0 N_19 GND mn5  l=0.5u w=0.6u m=1
M4 N_7 A1 N_20 GND mn5  l=0.5u w=0.6u m=1
M5 N_7 B0 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 C0 GND GND mn5  l=0.5u w=0.6u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_9 A2 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_9 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_9 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_9 B0 N_12 VDD mp5  l=0.42u w=0.62u m=1
M12 N_7 C0 N_12 VDD mp5  l=0.42u w=0.62u m=1
.ends aor311d1
* SPICE INPUT		Mon Sep 24 12:13:00 2018	aor311d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor311d2
.subckt aor311d2 C0 B0 A1 A0 A2 VDD Y GND
M1 Y N_7 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_19 A2 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_20 A0 N_19 GND mn5  l=0.5u w=0.6u m=1
M4 N_7 A1 N_20 GND mn5  l=0.5u w=0.6u m=1
M5 N_7 B0 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 C0 GND GND mn5  l=0.5u w=0.6u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 N_9 A2 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_9 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_9 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_9 B0 N_12 VDD mp5  l=0.42u w=0.62u m=1
M12 N_7 C0 N_12 VDD mp5  l=0.42u w=0.62u m=1
.ends aor311d2
* SPICE INPUT		Mon Sep 24 12:13:09 2018	aor31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d0
.subckt aor31d0 B0 A2 A1 A0 VDD Y GND
M1 N_11 A0 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 A1 N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_5 A2 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_5 B0 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 VDD A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 VDD A2 N_10 VDD mp5  l=0.42u w=0.62u m=1
M9 N_10 B0 N_5 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends aor31d0
* SPICE INPUT		Mon Sep 24 12:13:17 2018	aor31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d1
.subckt aor31d1 B0 A2 A1 A0 VDD Y GND
M1 N_11 A0 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_12 A1 N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_5 A2 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_5 B0 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 VDD A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 VDD A2 N_10 VDD mp5  l=0.42u w=0.62u m=1
M9 N_10 B0 N_5 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends aor31d1
* SPICE INPUT		Mon Sep 24 12:13:27 2018	aor31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d2
.subckt aor31d2 A0 A2 A1 B0 VDD Y GND
M1 N_5 B0 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_12 A1 N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_5 A2 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_11 A0 GND GND mn5  l=0.5u w=0.6u m=1
M6 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_9 B0 N_5 VDD mp5  l=0.42u w=0.62u m=1
M8 VDD A1 N_9 VDD mp5  l=0.42u w=0.62u m=1
M9 VDD A2 N_9 VDD mp5  l=0.42u w=0.62u m=1
M10 N_9 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends aor31d2
* SPICE INPUT		Mon Sep 24 12:13:36 2018	buffd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd0
.subckt buffd0 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends buffd0
* SPICE INPUT		Mon Sep 24 12:13:45 2018	buffd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd1
.subckt buffd1 VDD Y GND A
M1 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends buffd1
* SPICE INPUT		Mon Sep 24 12:13:54 2018	buffd10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd10
.subckt buffd10 GND Y VDD A
M1 GND A N_5 GND mn5  l=0.5u w=0.98u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.98u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M4 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M5 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M6 GND N_5 Y GND mn5  l=0.5u w=0.98u m=1
M7 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M8 VDD A N_5 VDD mp5  l=0.42u w=1.28u m=1
M9 N_5 A VDD VDD mp5  l=0.42u w=1.28u m=1
M10 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M11 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M13 VDD N_5 Y VDD mp5  l=0.42u w=1.28u m=1
M14 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends buffd10
* SPICE INPUT		Mon Sep 24 12:14:03 2018	buffd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd2
.subckt buffd2 GND Y VDD A
M1 Y N_4 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
M4 N_4 A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buffd2
* SPICE INPUT		Mon Sep 24 12:14:11 2018	buffd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd3
.subckt buffd3 VDD A GND Y
M1 N_6 A GND GND mn5  l=0.5u w=0.72u m=1
M2 GND N_6 Y GND mn5  l=0.5u w=0.766u m=1
M3 Y N_6 GND GND mn5  l=0.5u w=0.704u m=1
M4 VDD A N_6 VDD mp5  l=0.42u w=0.96u m=1
M5 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M6 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
.ends buffd3
* SPICE INPUT		Mon Sep 24 12:14:21 2018	buffd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd4
.subckt buffd4 Y GND VDD A
M1 GND N_4 Y GND mn5  l=0.5u w=0.98u m=1
M2 GND N_4 Y GND mn5  l=0.5u w=0.98u m=1
M3 GND A N_4 GND mn5  l=0.5u w=0.98u m=1
M4 VDD N_4 Y VDD mp5  l=0.42u w=1.28u m=1
M5 VDD N_4 Y VDD mp5  l=0.42u w=1.28u m=1
M6 VDD A N_4 VDD mp5  l=0.42u w=1.28u m=1
.ends buffd4
* SPICE INPUT		Mon Sep 24 12:14:32 2018	buffd5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd5
.subckt buffd5 GND Y VDD A
M1 GND N_4 Y GND mn5  l=0.5u w=0.98u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.735u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.735u m=1
M4 GND A N_4 GND mn5  l=0.5u w=0.98u m=1
M5 VDD N_4 Y VDD mp5  l=0.42u w=1.28u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 VDD A N_4 VDD mp5  l=0.42u w=1.28u m=1
.ends buffd5
* SPICE INPUT		Mon Sep 24 12:14:42 2018	buffd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd6
.subckt buffd6 GND Y VDD A
M1 GND A N_4 GND mn5  l=0.5u w=0.98u m=1
M2 Y N_4 GND GND mn5  l=0.5u w=0.98u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.98u m=1
M4 Y N_4 GND GND mn5  l=0.5u w=0.98u m=1
M5 VDD A N_4 VDD mp5  l=0.42u w=1.28u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 Y N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends buffd6
* SPICE INPUT		Mon Sep 24 12:14:51 2018	buffd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd8
.subckt buffd8 Y GND VDD A
M1 GND A N_5 GND mn5  l=0.5u w=0.98u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.49u m=1
M3 GND N_5 Y GND mn5  l=0.5u w=0.98u m=1
M4 GND N_5 Y GND mn5  l=0.5u w=0.98u m=1
M5 GND N_5 Y GND mn5  l=0.5u w=0.98u m=1
M6 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M7 VDD A N_5 VDD mp5  l=0.42u w=0.96u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.96u m=1
M9 VDD N_5 Y VDD mp5  l=0.42u w=1.28u m=1
M10 VDD N_5 Y VDD mp5  l=0.42u w=1.28u m=1
M11 VDD N_5 Y VDD mp5  l=0.42u w=1.28u m=1
M12 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends buffd8
* SPICE INPUT		Mon Sep 24 12:15:00 2018	buftd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd0
.subckt buftd0 A OE Y GND VDD
M1 N_3 OE GND GND mn5  l=0.5u w=0.6u m=1
M2 N_4 OE GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 N_4 GND mn5  l=0.5u w=0.6u m=1
M5 N_4 A GND GND mn5  l=0.5u w=0.6u m=1
M6 N_6 OE N_4 VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends buftd0
* SPICE INPUT		Mon Sep 24 12:15:08 2018	buftd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd1
.subckt buftd1 A OE Y GND VDD
M1 N_3 OE GND GND mn5  l=0.5u w=0.6u m=1
M2 N_4 OE GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_6 N_3 N_4 GND mn5  l=0.5u w=0.6u m=1
M5 N_4 A GND GND mn5  l=0.5u w=0.6u m=1
M6 N_6 OE N_4 VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends buftd1
* SPICE INPUT		Mon Sep 24 12:15:17 2018	buftd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd2
.subckt buftd2 A OE VDD Y GND
M1 N_3 OE GND GND mn5  l=0.5u w=0.6u m=1
M2 N_4 OE GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.96u m=1
M4 N_6 N_3 N_4 GND mn5  l=0.5u w=0.6u m=1
M5 N_4 A GND GND mn5  l=0.5u w=0.6u m=1
M6 N_6 OE N_4 VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M10 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends buftd2
* SPICE INPUT		Mon Sep 24 12:15:25 2018	buftld0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld0
.subckt buftld0 A OE VDD GND Y
M1 N_2 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 OE GND GND mn5  l=0.5u w=0.6u m=1
M3 N_6 OE N_2 GND mn5  l=0.5u w=0.6u m=1
M4 N_2 A GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_6 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M7 N_6 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends buftld0
* SPICE INPUT		Mon Sep 24 12:15:34 2018	buftld1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld1
.subckt buftld1 A OE GND VDD Y
M1 N_2 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 OE GND GND mn5  l=0.5u w=0.6u m=1
M3 N_6 OE N_2 GND mn5  l=0.5u w=0.6u m=1
M4 N_2 A GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_6 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_5 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_6 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
.ends buftld1
* SPICE INPUT		Mon Sep 24 12:15:43 2018	buftld2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftld2
.subckt buftld2 OE A GND VDD Y
M1 N_3 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 OE GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 A GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.98u m=1
M5 N_6 OE N_3 GND mn5  l=0.5u w=0.6u m=1
M6 N_6 A VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 N_6 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_5 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 N_5 N_3 VDD mp5  l=0.42u w=0.62u m=1
.ends buftld2
* SPICE INPUT		Mon Sep 24 12:15:52 2018	dfbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb1
.subckt dfbfb1 CKN D SN RN GND QN VDD Q
M1 N_9 RN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_19 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_57 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_10 N_5 N_57 GND mn5  l=0.5u w=0.6u m=1
M6 N_58 N_4 N_10 GND mn5  l=0.5u w=0.6u m=1
M7 N_58 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_4 CKN GND GND mn5  l=0.5u w=0.6u m=1
M9 N_59 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_11 N_4 N_59 GND mn5  l=0.5u w=0.6u m=1
M11 N_60 N_5 N_11 GND mn5  l=0.5u w=0.6u m=1
M12 N_60 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_26 SN GND GND mn5  l=0.5u w=0.6u m=1
M14 N_26 N_9 N_14 GND mn5  l=0.5u w=0.6u m=1
M15 N_26 N_11 N_14 GND mn5  l=0.5u w=0.6u m=1
M16 N_25 N_10 N_3 GND mn5  l=0.5u w=0.6u m=1
M17 N_25 N_9 N_3 GND mn5  l=0.5u w=0.6u m=1
M18 N_25 SN GND GND mn5  l=0.5u w=0.6u m=1
M19 Q N_19 GND GND mn5  l=0.5u w=0.72u m=1
M20 QN N_14 GND GND mn5  l=0.5u w=0.72u m=1
M21 N_9 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_19 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 Q N_19 VDD VDD mp5  l=0.42u w=0.96u m=1
M24 QN N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M25 N_32 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M26 N_32 N_5 N_11 VDD mp5  l=0.42u w=0.62u m=1
M27 N_33 N_4 N_11 VDD mp5  l=0.42u w=0.6u m=1
M28 N_33 N_14 VDD VDD mp5  l=0.42u w=0.6u m=1
M29 N_14 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_14 N_9 N_30 VDD mp5  l=0.42u w=0.62u m=1
M31 N_30 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_31 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_31 N_9 N_3 VDD mp5  l=0.42u w=0.62u m=1
M34 VDD SN N_3 VDD mp5  l=0.42u w=0.62u m=1
M35 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_34 D VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_35 N_5 N_10 VDD mp5  l=0.42u w=0.6u m=1
M38 N_34 N_4 N_10 VDD mp5  l=0.42u w=0.62u m=1
M39 N_35 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M40 N_4 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
.ends dfbfb1
* SPICE INPUT		Mon Sep 24 12:16:00 2018	dfbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb2
.subckt dfbfb2 SN D CKN RN QN VDD GND Q
M1 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_8 CKN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_58 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_58 N_8 N_4 GND mn5  l=0.5u w=0.6u m=1
M6 N_4 N_9 N_57 GND mn5  l=0.5u w=0.6u m=1
M7 N_9 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_57 D GND GND mn5  l=0.5u w=0.6u m=1
M9 N_25 N_13 N_3 GND mn5  l=0.5u w=0.6u m=1
M10 N_25 N_5 N_3 GND mn5  l=0.5u w=0.6u m=1
M11 N_25 SN GND GND mn5  l=0.5u w=0.6u m=1
M12 N_60 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_60 N_9 N_13 GND mn5  l=0.5u w=0.6u m=1
M14 N_13 N_8 N_59 GND mn5  l=0.5u w=0.6u m=1
M15 N_59 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_24 SN GND GND mn5  l=0.5u w=0.6u m=1
M17 N_24 N_5 N_7 GND mn5  l=0.5u w=0.6u m=1
M18 N_24 N_4 N_7 GND mn5  l=0.5u w=0.6u m=1
M19 QN N_3 GND GND mn5  l=0.5u w=0.96u m=1
M20 Q N_2 GND GND mn5  l=0.5u w=0.96u m=1
M21 N_30 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_3 N_5 N_30 VDD mp5  l=0.42u w=0.62u m=1
M23 N_3 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_33 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 N_33 N_8 N_13 VDD mp5  l=0.42u w=0.6u m=1
M26 N_32 N_9 N_13 VDD mp5  l=0.42u w=0.62u m=1
M27 N_32 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 VDD SN N_7 VDD mp5  l=0.42u w=0.62u m=1
M29 N_31 N_5 N_7 VDD mp5  l=0.42u w=0.62u m=1
M30 N_31 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_8 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_35 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M33 N_34 N_8 N_4 VDD mp5  l=0.42u w=0.62u m=1
M34 N_35 N_9 N_4 VDD mp5  l=0.42u w=0.6u m=1
M35 N_9 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_34 D VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_2 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M38 N_5 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M39 QN N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M40 Q N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends dfbfb2
* SPICE INPUT		Mon Sep 24 12:16:09 2018	dfbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb1
.subckt dfbrb1 SN D CK RN Q QN VDD GND
M1 QN N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_20 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_20 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_3 RN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_7 CK GND GND mn5  l=0.5u w=0.6u m=1
M6 N_31 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_31 N_6 N_2 GND mn5  l=0.5u w=0.6u m=1
M8 N_2 N_7 N_30 GND mn5  l=0.5u w=0.6u m=1
M9 N_6 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_30 D GND GND mn5  l=0.5u w=0.6u m=1
M11 N_25 N_11 N_8 GND mn5  l=0.5u w=0.6u m=1
M12 N_25 N_3 N_8 GND mn5  l=0.5u w=0.6u m=1
M13 N_25 SN GND GND mn5  l=0.5u w=0.6u m=1
M14 N_33 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_33 N_7 N_11 GND mn5  l=0.5u w=0.6u m=1
M16 N_11 N_6 N_32 GND mn5  l=0.5u w=0.6u m=1
M17 N_32 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M18 N_24 SN GND GND mn5  l=0.5u w=0.6u m=1
M19 N_24 N_3 N_5 GND mn5  l=0.5u w=0.6u m=1
M20 N_24 N_2 N_5 GND mn5  l=0.5u w=0.6u m=1
M21 N_53 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_8 N_3 N_53 VDD mp5  l=0.42u w=0.62u m=1
M23 N_8 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_56 N_8 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 N_56 N_6 N_11 VDD mp5  l=0.42u w=0.6u m=1
M26 N_55 N_7 N_11 VDD mp5  l=0.42u w=0.62u m=1
M27 N_55 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 VDD SN N_5 VDD mp5  l=0.42u w=0.62u m=1
M29 N_54 N_3 N_5 VDD mp5  l=0.42u w=0.62u m=1
M30 N_54 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_7 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_58 N_5 VDD VDD mp5  l=0.42u w=0.6u m=1
M33 N_57 N_6 N_2 VDD mp5  l=0.42u w=0.62u m=1
M34 N_58 N_7 N_2 VDD mp5  l=0.42u w=0.6u m=1
M35 N_6 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_57 D VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_20 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M38 N_3 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M39 QN N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M40 Q N_20 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfbrb1
* SPICE INPUT		Mon Sep 24 12:16:17 2018	dfbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb2
.subckt dfbrb2 SN D CK RN Q QN VDD GND
M1 QN N_8 GND GND mn5  l=0.5u w=0.98u m=1
M2 Q N_20 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_20 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_3 RN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_7 CK GND GND mn5  l=0.5u w=0.6u m=1
M6 N_58 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_58 N_6 N_2 GND mn5  l=0.5u w=0.6u m=1
M8 N_2 N_7 N_57 GND mn5  l=0.5u w=0.6u m=1
M9 N_6 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_57 D GND GND mn5  l=0.5u w=0.6u m=1
M11 N_25 N_11 N_8 GND mn5  l=0.5u w=0.6u m=1
M12 N_25 N_3 N_8 GND mn5  l=0.5u w=0.6u m=1
M13 N_25 SN GND GND mn5  l=0.5u w=0.6u m=1
M14 N_60 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_60 N_7 N_11 GND mn5  l=0.5u w=0.6u m=1
M16 N_11 N_6 N_59 GND mn5  l=0.5u w=0.6u m=1
M17 N_59 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M18 N_24 SN GND GND mn5  l=0.5u w=0.6u m=1
M19 N_24 N_3 N_5 GND mn5  l=0.5u w=0.6u m=1
M20 N_24 N_2 N_5 GND mn5  l=0.5u w=0.6u m=1
M21 N_30 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_8 N_3 N_30 VDD mp5  l=0.42u w=0.62u m=1
M23 N_8 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_33 N_8 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 N_33 N_6 N_11 VDD mp5  l=0.42u w=0.6u m=1
M26 N_32 N_7 N_11 VDD mp5  l=0.42u w=0.62u m=1
M27 N_32 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 VDD SN N_5 VDD mp5  l=0.42u w=0.62u m=1
M29 N_31 N_3 N_5 VDD mp5  l=0.42u w=0.62u m=1
M30 N_31 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_7 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_35 N_5 VDD VDD mp5  l=0.42u w=0.6u m=1
M33 N_34 N_6 N_2 VDD mp5  l=0.42u w=0.62u m=1
M34 N_35 N_7 N_2 VDD mp5  l=0.42u w=0.6u m=1
M35 N_6 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_34 D VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_20 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M38 N_3 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M39 QN N_8 VDD VDD mp5  l=0.42u w=1.28u m=1
M40 Q N_20 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends dfbrb2
* SPICE INPUT		Mon Sep 24 12:16:26 2018	dfbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq1
.subckt dfbrq1 VDD Q GND SN D RN CK
M1 N_4 N_16 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_55 D GND GND mn5  l=0.5u w=0.6u m=1
M3 N_6 N_16 N_55 GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_4 N_54 GND mn5  l=0.5u w=0.6u m=1
M5 N_54 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_10 N_4 N_56 GND mn5  l=0.5u w=0.6u m=1
M7 N_12 N_10 N_29 GND mn5  l=0.5u w=0.6u m=1
M8 N_29 SN GND GND mn5  l=0.5u w=0.6u m=1
M9 N_29 N_3 N_12 GND mn5  l=0.5u w=0.6u m=1
M10 N_57 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_28 N_6 N_9 GND mn5  l=0.5u w=0.6u m=1
M12 N_56 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_28 N_3 N_9 GND mn5  l=0.5u w=0.6u m=1
M14 N_57 N_16 N_10 GND mn5  l=0.5u w=0.6u m=1
M15 GND SN N_28 GND mn5  l=0.5u w=0.6u m=1
M16 N_25 SN GND GND mn5  l=0.5u w=0.72u m=1
M17 N_3 RN GND GND mn5  l=0.5u w=0.6u m=1
M18 N_25 N_3 Q GND mn5  l=0.5u w=0.72u m=1
M19 Q N_10 N_25 GND mn5  l=0.5u w=0.72u m=1
M20 N_16 CK GND GND mn5  l=0.5u w=0.6u m=1
M21 N_22 N_4 N_10 VDD mp5  l=0.42u w=0.6u m=1
M22 VDD N_16 N_4 VDD mp5  l=0.42u w=0.62u m=1
M23 N_18 D VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_23 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 N_12 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M26 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_3 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_23 N_3 N_12 VDD mp5  l=0.42u w=0.6u m=1
M29 N_22 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M30 N_18 N_4 N_6 VDD mp5  l=0.42u w=0.62u m=1
M31 N_19 N_16 N_6 VDD mp5  l=0.42u w=0.6u m=1
M32 N_19 N_9 VDD VDD mp5  l=0.42u w=0.6u m=1
M33 N_20 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M34 Q N_3 N_24 VDD mp5  l=0.42u w=0.96u m=1
M35 N_10 N_16 N_21 VDD mp5  l=0.42u w=0.62u m=1
M36 N_21 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_9 N_3 N_20 VDD mp5  l=0.42u w=0.62u m=1
M38 N_24 N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
M39 N_9 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M40 N_16 CK VDD VDD mp5  l=0.42u w=0.6u m=1
.ends dfbrq1
* SPICE INPUT		Mon Sep 24 12:16:35 2018	dfbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq2
.subckt dfbrq2 VDD Q GND SN D RN CK
M1 N_4 N_16 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_55 D GND GND mn5  l=0.5u w=0.6u m=1
M3 N_6 N_16 N_55 GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_4 N_54 GND mn5  l=0.5u w=0.6u m=1
M5 N_54 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_10 N_4 N_56 GND mn5  l=0.5u w=0.6u m=1
M7 N_12 N_10 N_29 GND mn5  l=0.5u w=0.6u m=1
M8 N_29 SN GND GND mn5  l=0.5u w=0.6u m=1
M9 N_29 N_3 N_12 GND mn5  l=0.5u w=0.6u m=1
M10 N_57 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_28 N_6 N_9 GND mn5  l=0.5u w=0.6u m=1
M12 N_56 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_28 N_3 N_9 GND mn5  l=0.5u w=0.6u m=1
M14 N_57 N_16 N_10 GND mn5  l=0.5u w=0.6u m=1
M15 GND SN N_28 GND mn5  l=0.5u w=0.6u m=1
M16 N_25 SN GND GND mn5  l=0.5u w=0.98u m=1
M17 N_3 RN GND GND mn5  l=0.5u w=0.6u m=1
M18 N_25 N_3 Q GND mn5  l=0.5u w=0.98u m=1
M19 Q N_10 N_25 GND mn5  l=0.5u w=0.98u m=1
M20 N_16 CK GND GND mn5  l=0.5u w=0.6u m=1
M21 N_22 N_4 N_10 VDD mp5  l=0.42u w=0.6u m=1
M22 VDD N_16 N_4 VDD mp5  l=0.42u w=0.62u m=1
M23 N_18 D VDD VDD mp5  l=0.42u w=0.62u m=1
M24 VDD N_10 N_23 VDD mp5  l=0.42u w=0.6u m=1
M25 N_12 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M26 Q SN VDD VDD mp5  l=0.42u w=1.28u m=1
M27 N_3 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_23 N_3 N_12 VDD mp5  l=0.42u w=0.6u m=1
M29 N_22 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M30 N_18 N_4 N_6 VDD mp5  l=0.42u w=0.62u m=1
M31 N_19 N_16 N_6 VDD mp5  l=0.42u w=0.6u m=1
M32 N_19 N_9 VDD VDD mp5  l=0.42u w=0.6u m=1
M33 N_20 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M34 Q N_3 N_24 VDD mp5  l=0.42u w=1.28u m=1
M35 N_10 N_16 N_21 VDD mp5  l=0.42u w=0.62u m=1
M36 N_21 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_9 N_3 N_20 VDD mp5  l=0.42u w=0.62u m=1
M38 N_24 N_10 VDD VDD mp5  l=0.42u w=1.28u m=1
M39 N_9 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M40 N_16 CK VDD VDD mp5  l=0.42u w=0.6u m=1
.ends dfbrq2
* SPICE INPUT		Mon Sep 24 12:16:43 2018	dfcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb1
.subckt dfcfb1 VDD QN Q GND D RN CKN
M1 N_13 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_14 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 CKN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_48 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_6 N_48 GND mn5  l=0.5u w=0.6u m=1
M7 N_49 N_3 N_7 GND mn5  l=0.5u w=0.6u m=1
M8 N_49 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_50 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_51 N_6 N_17 GND mn5  l=0.5u w=0.6u m=1
M13 N_17 N_3 N_50 GND mn5  l=0.5u w=0.6u m=1
M14 N_51 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M15 GND N_17 N_15 GND mn5  l=0.5u w=0.6u m=1
M16 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M17 QN N_15 GND GND mn5  l=0.5u w=0.72u m=1
M18 Q N_13 GND GND mn5  l=0.5u w=0.72u m=1
M19 N_3 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
M20 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_3 N_7 VDD mp5  l=0.42u w=0.62u m=1
M23 N_22 N_6 N_7 VDD mp5  l=0.42u w=0.6u m=1
M24 N_22 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_7 N_20 VDD mp5  l=0.42u w=0.62u m=1
M26 N_20 N_14 N_4 VDD mp5  l=0.42u w=0.62u m=1
M27 QN N_15 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 Q N_13 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_13 N_15 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_14 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_24 N_6 N_17 VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 N_3 N_17 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD N_15 N_25 VDD mp5  l=0.42u w=0.6u m=1
M35 VDD N_17 N_23 VDD mp5  l=0.42u w=0.62u m=1
M36 N_15 N_14 N_23 VDD mp5  l=0.42u w=0.62u m=1
.ends dfcfb1
* SPICE INPUT		Mon Sep 24 12:16:52 2018	dfcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb2
.subckt dfcfb2 VDD QN Q GND D RN CKN
M1 N_13 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_14 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 CKN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_48 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_6 N_48 GND mn5  l=0.5u w=0.6u m=1
M7 N_49 N_3 N_7 GND mn5  l=0.5u w=0.6u m=1
M8 N_49 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_50 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_51 N_6 N_17 GND mn5  l=0.5u w=0.6u m=1
M13 N_17 N_3 N_50 GND mn5  l=0.5u w=0.6u m=1
M14 N_51 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M15 GND N_17 N_15 GND mn5  l=0.5u w=0.6u m=1
M16 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M17 QN N_15 GND GND mn5  l=0.5u w=0.98u m=1
M18 Q N_13 GND GND mn5  l=0.5u w=0.98u m=1
M19 N_3 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
M20 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_3 N_7 VDD mp5  l=0.42u w=0.62u m=1
M23 N_22 N_6 N_7 VDD mp5  l=0.42u w=0.6u m=1
M24 N_22 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_7 N_20 VDD mp5  l=0.42u w=0.62u m=1
M26 N_20 N_14 N_4 VDD mp5  l=0.42u w=0.62u m=1
M27 QN N_15 VDD VDD mp5  l=0.42u w=1.28u m=1
M28 Q N_13 VDD VDD mp5  l=0.42u w=1.28u m=1
M29 N_13 N_15 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_14 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_24 N_6 N_17 VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 N_3 N_17 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD N_15 N_25 VDD mp5  l=0.42u w=0.6u m=1
M35 VDD N_17 N_23 VDD mp5  l=0.42u w=0.62u m=1
M36 N_15 N_14 N_23 VDD mp5  l=0.42u w=0.62u m=1
.ends dfcfb2
* SPICE INPUT		Mon Sep 24 12:17:01 2018	dfcfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfq1
.subckt dfcfq1 VDD Q GND D RN CKN
M1 N_12 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_13 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 CKN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_46 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_6 N_46 GND mn5  l=0.5u w=0.6u m=1
M7 N_47 N_3 N_7 GND mn5  l=0.5u w=0.6u m=1
M8 N_47 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_48 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_49 N_6 N_16 GND mn5  l=0.5u w=0.6u m=1
M13 N_16 N_3 N_48 GND mn5  l=0.5u w=0.6u m=1
M14 N_49 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 GND N_16 N_14 GND mn5  l=0.5u w=0.6u m=1
M16 N_14 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M17 Q N_12 GND GND mn5  l=0.5u w=0.72u m=1
M18 N_3 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
M19 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_20 D VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_20 N_3 N_7 VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_6 N_7 VDD mp5  l=0.42u w=0.6u m=1
M23 N_21 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M24 VDD N_7 N_19 VDD mp5  l=0.42u w=0.62u m=1
M25 N_19 N_13 N_4 VDD mp5  l=0.42u w=0.62u m=1
M26 Q N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 N_12 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_13 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_23 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_23 N_6 N_16 VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 N_3 N_16 VDD mp5  l=0.42u w=0.6u m=1
M32 VDD N_14 N_24 VDD mp5  l=0.42u w=0.6u m=1
M33 VDD N_16 N_22 VDD mp5  l=0.42u w=0.62u m=1
M34 N_14 N_13 N_22 VDD mp5  l=0.42u w=0.62u m=1
.ends dfcfq1
* SPICE INPUT		Mon Sep 24 12:17:09 2018	dfcfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfq2
.subckt dfcfq2 VDD Q GND D RN CKN
M1 N_12 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_13 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 CKN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_46 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_6 N_46 GND mn5  l=0.5u w=0.6u m=1
M7 N_47 N_3 N_7 GND mn5  l=0.5u w=0.6u m=1
M8 N_47 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_48 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_49 N_6 N_16 GND mn5  l=0.5u w=0.6u m=1
M13 N_16 N_3 N_48 GND mn5  l=0.5u w=0.6u m=1
M14 N_49 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 GND N_16 N_14 GND mn5  l=0.5u w=0.6u m=1
M16 N_14 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M17 Q N_12 GND GND mn5  l=0.5u w=0.98u m=1
M18 N_3 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
M19 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_20 D VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_20 N_3 N_7 VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_6 N_7 VDD mp5  l=0.42u w=0.6u m=1
M23 N_21 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M24 VDD N_7 N_19 VDD mp5  l=0.42u w=0.62u m=1
M25 N_19 N_13 N_4 VDD mp5  l=0.42u w=0.62u m=1
M26 Q N_12 VDD VDD mp5  l=0.42u w=1.28u m=1
M27 N_12 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_13 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_23 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_23 N_6 N_16 VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 N_3 N_16 VDD mp5  l=0.42u w=0.6u m=1
M32 VDD N_14 N_24 VDD mp5  l=0.42u w=0.6u m=1
M33 VDD N_16 N_22 VDD mp5  l=0.42u w=0.62u m=1
M34 N_14 N_13 N_22 VDD mp5  l=0.42u w=0.62u m=1
.ends dfcfq2
* SPICE INPUT		Mon Sep 24 12:17:17 2018	dfcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb1
.subckt dfcrb1 VDD QN Q GND D RN CK
M1 N_13 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_14 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_48 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_3 N_48 GND mn5  l=0.5u w=0.6u m=1
M7 N_49 N_6 N_7 GND mn5  l=0.5u w=0.6u m=1
M8 N_49 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_50 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_51 N_3 N_17 GND mn5  l=0.5u w=0.6u m=1
M13 N_17 N_6 N_50 GND mn5  l=0.5u w=0.6u m=1
M14 N_51 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M15 GND N_17 N_15 GND mn5  l=0.5u w=0.6u m=1
M16 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M17 QN N_15 GND GND mn5  l=0.5u w=0.72u m=1
M18 Q N_13 GND GND mn5  l=0.5u w=0.72u m=1
M19 N_3 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M20 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_6 N_7 VDD mp5  l=0.42u w=0.62u m=1
M23 N_22 N_3 N_7 VDD mp5  l=0.42u w=0.6u m=1
M24 N_22 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_7 N_20 VDD mp5  l=0.42u w=0.62u m=1
M26 N_20 N_14 N_4 VDD mp5  l=0.42u w=0.62u m=1
M27 QN N_15 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 Q N_13 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_13 N_15 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_14 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_24 N_3 N_17 VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 N_6 N_17 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD N_15 N_25 VDD mp5  l=0.42u w=0.6u m=1
M35 VDD N_17 N_23 VDD mp5  l=0.42u w=0.62u m=1
M36 N_15 N_14 N_23 VDD mp5  l=0.42u w=0.62u m=1
.ends dfcrb1
* SPICE INPUT		Mon Sep 24 12:17:26 2018	dfcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb2
.subckt dfcrb2 VDD QN Q GND D RN CK
M1 N_13 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_14 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_48 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_3 N_48 GND mn5  l=0.5u w=0.6u m=1
M7 N_49 N_6 N_7 GND mn5  l=0.5u w=0.6u m=1
M8 N_49 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_50 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_51 N_3 N_17 GND mn5  l=0.5u w=0.6u m=1
M13 N_17 N_6 N_50 GND mn5  l=0.5u w=0.6u m=1
M14 N_51 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M15 GND N_17 N_15 GND mn5  l=0.5u w=0.6u m=1
M16 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M17 QN N_15 GND GND mn5  l=0.5u w=0.98u m=1
M18 Q N_13 GND GND mn5  l=0.5u w=0.98u m=1
M19 N_3 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M20 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_21 D VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_6 N_7 VDD mp5  l=0.42u w=0.62u m=1
M23 N_22 N_3 N_7 VDD mp5  l=0.42u w=0.6u m=1
M24 N_22 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_7 N_20 VDD mp5  l=0.42u w=0.62u m=1
M26 N_20 N_14 N_4 VDD mp5  l=0.42u w=0.62u m=1
M27 QN N_15 VDD VDD mp5  l=0.42u w=1.28u m=1
M28 Q N_13 VDD VDD mp5  l=0.42u w=1.28u m=1
M29 N_13 N_15 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_14 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_24 N_3 N_17 VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 N_6 N_17 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD N_15 N_25 VDD mp5  l=0.42u w=0.6u m=1
M35 VDD N_17 N_23 VDD mp5  l=0.42u w=0.62u m=1
M36 N_15 N_14 N_23 VDD mp5  l=0.42u w=0.62u m=1
.ends dfcrb2
* SPICE INPUT		Mon Sep 24 12:17:35 2018	dfcrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrn1
.subckt dfcrn1 VDD QN GND D CK RN
M1 N_15 RN GND GND mn5  l=0.5u w=0.6u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M4 N_9 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M5 GND N_11 N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_45 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_11 N_6 N_44 GND mn5  l=0.5u w=0.6u m=1
M8 N_45 N_3 N_11 GND mn5  l=0.5u w=0.6u m=1
M9 N_44 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_4 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_43 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_43 N_6 N_7 GND mn5  l=0.5u w=0.6u m=1
M15 N_7 N_3 N_42 GND mn5  l=0.5u w=0.6u m=1
M16 N_42 D GND GND mn5  l=0.5u w=0.6u m=1
M17 N_3 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M18 N_17 N_15 N_4 VDD mp5  l=0.42u w=0.62u m=1
M19 VDD N_7 N_17 VDD mp5  l=0.42u w=0.62u m=1
M20 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_19 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_19 N_3 N_7 VDD mp5  l=0.42u w=0.6u m=1
M23 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.62u m=1
M24 N_18 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_9 N_15 N_20 VDD mp5  l=0.42u w=0.62u m=1
M26 VDD N_11 N_20 VDD mp5  l=0.42u w=0.62u m=1
M27 VDD N_9 N_22 VDD mp5  l=0.42u w=0.6u m=1
M28 N_22 N_6 N_11 VDD mp5  l=0.42u w=0.6u m=1
M29 N_21 N_3 N_11 VDD mp5  l=0.42u w=0.62u m=1
M30 N_21 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_15 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M32 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfcrn1
* SPICE INPUT		Mon Sep 24 12:17:43 2018	dfcrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrn2
.subckt dfcrn2 VDD QN GND D RN CK
M1 QN N_12 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_11 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_42 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_3 N_42 GND mn5  l=0.5u w=0.6u m=1
M7 N_43 N_6 N_7 GND mn5  l=0.5u w=0.6u m=1
M8 N_43 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_44 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_45 N_3 N_14 GND mn5  l=0.5u w=0.6u m=1
M13 N_14 N_6 N_44 GND mn5  l=0.5u w=0.6u m=1
M14 N_45 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M15 GND N_14 N_12 GND mn5  l=0.5u w=0.6u m=1
M16 N_12 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M17 N_3 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M18 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_18 D VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_18 N_6 N_7 VDD mp5  l=0.42u w=0.62u m=1
M21 N_19 N_3 N_7 VDD mp5  l=0.42u w=0.6u m=1
M22 N_19 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M23 VDD N_7 N_17 VDD mp5  l=0.42u w=0.62u m=1
M24 N_17 N_11 N_4 VDD mp5  l=0.42u w=0.62u m=1
M25 QN N_12 VDD VDD mp5  l=0.42u w=1.28u m=1
M26 N_11 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M27 N_21 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_21 N_3 N_14 VDD mp5  l=0.42u w=0.62u m=1
M29 N_22 N_6 N_14 VDD mp5  l=0.42u w=0.6u m=1
M30 VDD N_12 N_22 VDD mp5  l=0.42u w=0.6u m=1
M31 VDD N_14 N_20 VDD mp5  l=0.42u w=0.62u m=1
M32 N_12 N_11 N_20 VDD mp5  l=0.42u w=0.62u m=1
.ends dfcrn2
* SPICE INPUT		Mon Sep 24 12:17:52 2018	dfcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq1
.subckt dfcrq1 VDD Q GND D CK RN
M1 N_11 CK GND GND mn5  l=0.5u w=0.6u m=1
M2 Q N_14 GND GND mn5  l=0.5u w=0.72u m=1
M3 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_12 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_12 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_30 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_14 N_4 N_29 GND mn5  l=0.5u w=0.6u m=1
M8 N_30 N_11 N_14 GND mn5  l=0.5u w=0.6u m=1
M9 N_29 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_2 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_2 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_28 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_8 RN GND GND mn5  l=0.5u w=0.6u m=1
M14 N_28 N_4 N_5 GND mn5  l=0.5u w=0.6u m=1
M15 N_5 N_11 N_27 GND mn5  l=0.5u w=0.6u m=1
M16 N_27 D GND GND mn5  l=0.5u w=0.6u m=1
M17 N_4 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M18 N_17 N_8 N_2 VDD mp5  l=0.42u w=0.62u m=1
M19 VDD N_5 N_17 VDD mp5  l=0.42u w=0.62u m=1
M20 N_19 N_2 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_19 N_11 N_5 VDD mp5  l=0.42u w=0.6u m=1
M22 N_18 N_4 N_5 VDD mp5  l=0.42u w=0.62u m=1
M23 N_18 D VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_4 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_20 N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 N_20 N_8 Q VDD mp5  l=0.42u w=0.96u m=1
M27 N_8 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_11 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M29 N_12 N_8 N_21 VDD mp5  l=0.42u w=0.62u m=1
M30 VDD N_14 N_21 VDD mp5  l=0.42u w=0.62u m=1
M31 N_23 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_23 N_4 N_14 VDD mp5  l=0.42u w=0.6u m=1
M33 N_22 N_11 N_14 VDD mp5  l=0.42u w=0.62u m=1
M34 N_22 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends dfcrq1
* SPICE INPUT		Mon Sep 24 12:18:01 2018	dfcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq2
.subckt dfcrq2 VDD Q GND D CK RN
M1 N_11 CK GND GND mn5  l=0.5u w=0.6u m=1
M2 Q N_14 GND GND mn5  l=0.5u w=0.98u m=1
M3 Q N_8 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_12 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_12 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_30 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_14 N_4 N_29 GND mn5  l=0.5u w=0.6u m=1
M8 N_30 N_11 N_14 GND mn5  l=0.5u w=0.6u m=1
M9 N_29 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_2 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_2 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_28 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_8 RN GND GND mn5  l=0.5u w=0.6u m=1
M14 N_28 N_4 N_5 GND mn5  l=0.5u w=0.6u m=1
M15 N_5 N_11 N_27 GND mn5  l=0.5u w=0.6u m=1
M16 N_27 D GND GND mn5  l=0.5u w=0.6u m=1
M17 N_4 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M18 N_17 N_8 N_2 VDD mp5  l=0.42u w=0.62u m=1
M19 VDD N_5 N_17 VDD mp5  l=0.42u w=0.62u m=1
M20 N_19 N_2 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_19 N_11 N_5 VDD mp5  l=0.42u w=0.6u m=1
M22 N_18 N_4 N_5 VDD mp5  l=0.42u w=0.62u m=1
M23 N_18 D VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_4 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_20 N_14 VDD VDD mp5  l=0.42u w=1.28u m=1
M26 N_20 N_8 Q VDD mp5  l=0.42u w=1.28u m=1
M27 N_8 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_11 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M29 N_12 N_8 N_21 VDD mp5  l=0.42u w=0.62u m=1
M30 VDD N_14 N_21 VDD mp5  l=0.42u w=0.62u m=1
M31 N_23 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_23 N_4 N_14 VDD mp5  l=0.42u w=0.6u m=1
M33 N_22 N_11 N_14 VDD mp5  l=0.42u w=0.62u m=1
M34 N_22 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends dfcrq2
* SPICE INPUT		Mon Sep 24 12:18:09 2018	dfnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb1
.subckt dfnfb1 D CKN GND Q QN VDD
M1 N_22 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_22 N_6 N_3 GND mn5  l=0.5u w=0.6u m=1
M3 N_3 N_4 N_21 GND mn5  l=0.5u w=0.6u m=1
M4 N_21 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_4 CKN GND GND mn5  l=0.5u w=0.6u m=1
M7 N_8 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_24 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_24 N_4 N_9 GND mn5  l=0.5u w=0.6u m=1
M10 N_9 N_6 N_23 GND mn5  l=0.5u w=0.6u m=1
M11 N_23 D GND GND mn5  l=0.5u w=0.6u m=1
M12 N_6 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M13 Q N_3 GND GND mn5  l=0.5u w=0.72u m=1
M14 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M15 N_41 N_2 VDD VDD mp5  l=0.42u w=0.6u m=1
M16 N_41 N_4 N_3 VDD mp5  l=0.42u w=0.6u m=1
M17 N_40 N_6 N_3 VDD mp5  l=0.42u w=0.62u m=1
M18 N_40 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_2 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_8 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_43 N_8 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_43 N_6 N_9 VDD mp5  l=0.42u w=0.6u m=1
M23 N_42 N_4 N_9 VDD mp5  l=0.42u w=0.62u m=1
M24 N_42 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_6 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M26 N_4 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
M27 Q N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfnfb1
* SPICE INPUT		Mon Sep 24 12:18:18 2018	dfnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb2
.subckt dfnfb2 D CKN GND Q QN VDD
M1 N_41 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_41 N_6 N_3 GND mn5  l=0.5u w=0.6u m=1
M3 N_3 N_4 N_40 GND mn5  l=0.5u w=0.6u m=1
M4 N_40 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_4 CKN GND GND mn5  l=0.5u w=0.6u m=1
M7 N_8 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_43 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_43 N_4 N_9 GND mn5  l=0.5u w=0.6u m=1
M10 N_9 N_6 N_42 GND mn5  l=0.5u w=0.6u m=1
M11 N_42 D GND GND mn5  l=0.5u w=0.6u m=1
M12 N_6 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M13 Q N_3 GND GND mn5  l=0.5u w=0.98u m=1
M14 QN N_2 GND GND mn5  l=0.5u w=0.98u m=1
M15 N_22 N_2 VDD VDD mp5  l=0.42u w=0.6u m=1
M16 N_22 N_4 N_3 VDD mp5  l=0.42u w=0.6u m=1
M17 N_21 N_6 N_3 VDD mp5  l=0.42u w=0.62u m=1
M18 N_21 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_2 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_8 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_24 N_8 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_24 N_6 N_9 VDD mp5  l=0.42u w=0.6u m=1
M23 N_23 N_4 N_9 VDD mp5  l=0.42u w=0.62u m=1
M24 N_23 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_6 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M26 N_4 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
M27 Q N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M28 QN N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends dfnfb2
* SPICE INPUT		Mon Sep 24 12:18:27 2018	dfnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb1
.subckt dfnrb1 CK D GND Q QN VDD
M1 N_41 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_41 N_5 N_3 GND mn5  l=0.5u w=0.6u m=1
M3 N_3 N_8 N_40 GND mn5  l=0.5u w=0.6u m=1
M4 N_40 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_9 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_43 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_43 N_8 N_10 GND mn5  l=0.5u w=0.6u m=1
M9 N_10 N_5 N_42 GND mn5  l=0.5u w=0.6u m=1
M10 N_42 D GND GND mn5  l=0.5u w=0.6u m=1
M11 GND N_5 N_8 GND mn5  l=0.5u w=0.6u m=1
M12 N_5 CK GND GND mn5  l=0.5u w=0.6u m=1
M13 Q N_3 GND GND mn5  l=0.5u w=0.72u m=1
M14 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M15 N_22 N_2 VDD VDD mp5  l=0.42u w=0.6u m=1
M16 N_22 N_8 N_3 VDD mp5  l=0.42u w=0.6u m=1
M17 N_21 N_5 N_3 VDD mp5  l=0.42u w=0.62u m=1
M18 N_21 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_2 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_9 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_24 N_9 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_24 N_5 N_10 VDD mp5  l=0.42u w=0.6u m=1
M23 N_23 N_8 N_10 VDD mp5  l=0.42u w=0.62u m=1
M24 N_23 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_8 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M26 N_5 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M27 Q N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfnrb1
* SPICE INPUT		Mon Sep 24 12:18:35 2018	dfnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb2
.subckt dfnrb2 CK D GND Q QN VDD
M1 N_41 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_41 N_5 N_3 GND mn5  l=0.5u w=0.6u m=1
M3 N_3 N_8 N_40 GND mn5  l=0.5u w=0.6u m=1
M4 N_40 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_9 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_43 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_43 N_8 N_10 GND mn5  l=0.5u w=0.6u m=1
M9 N_10 N_5 N_42 GND mn5  l=0.5u w=0.6u m=1
M10 N_42 D GND GND mn5  l=0.5u w=0.6u m=1
M11 GND N_5 N_8 GND mn5  l=0.5u w=0.6u m=1
M12 N_5 CK GND GND mn5  l=0.5u w=0.6u m=1
M13 Q N_3 GND GND mn5  l=0.5u w=0.98u m=1
M14 QN N_2 GND GND mn5  l=0.5u w=0.98u m=1
M15 N_22 N_2 VDD VDD mp5  l=0.42u w=0.6u m=1
M16 N_22 N_8 N_3 VDD mp5  l=0.42u w=0.6u m=1
M17 N_21 N_5 N_3 VDD mp5  l=0.42u w=0.62u m=1
M18 N_21 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_2 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_9 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_24 N_9 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_24 N_5 N_10 VDD mp5  l=0.42u w=0.6u m=1
M23 N_23 N_8 N_10 VDD mp5  l=0.42u w=0.62u m=1
M24 N_23 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_8 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M26 N_5 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M27 Q N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M28 QN N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends dfnrb2
* SPICE INPUT		Mon Sep 24 12:18:44 2018	dfnrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrn1
.subckt dfnrn1 CK D GND VDD QN
M1 N_38 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_11 N_6 N_38 GND mn5  l=0.5u w=0.6u m=1
M3 N_39 N_7 N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_2 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_39 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M6 GND N_7 N_6 GND mn5  l=0.5u w=0.6u m=1
M7 N_40 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_4 N_7 N_40 GND mn5  l=0.5u w=0.6u m=1
M9 N_41 N_6 N_4 GND mn5  l=0.5u w=0.6u m=1
M10 N_41 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_7 CK GND GND mn5  l=0.5u w=0.6u m=1
M13 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M14 N_20 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_20 N_7 N_11 VDD mp5  l=0.42u w=0.62u m=1
M16 N_2 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_21 N_6 N_11 VDD mp5  l=0.42u w=0.6u m=1
M18 N_21 N_2 VDD VDD mp5  l=0.42u w=0.6u m=1
M19 N_7 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M20 N_6 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_22 D VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_22 N_6 N_4 VDD mp5  l=0.42u w=0.62u m=1
M23 N_23 N_7 N_4 VDD mp5  l=0.42u w=0.6u m=1
M24 N_23 N_5 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M26 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfnrn1
* SPICE INPUT		Mon Sep 24 12:18:54 2018	dfnrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrn2
.subckt dfnrn2 CK D GND VDD QN
M1 N_38 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_11 N_6 N_38 GND mn5  l=0.5u w=0.6u m=1
M3 N_39 N_7 N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_2 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_39 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M6 GND N_7 N_6 GND mn5  l=0.5u w=0.6u m=1
M7 N_40 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_4 N_7 N_40 GND mn5  l=0.5u w=0.6u m=1
M9 N_41 N_6 N_4 GND mn5  l=0.5u w=0.6u m=1
M10 N_41 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_7 CK GND GND mn5  l=0.5u w=0.6u m=1
M13 QN N_2 GND GND mn5  l=0.5u w=0.98u m=1
M14 N_20 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_20 N_7 N_11 VDD mp5  l=0.42u w=0.62u m=1
M16 N_2 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_21 N_6 N_11 VDD mp5  l=0.42u w=0.6u m=1
M18 N_21 N_2 VDD VDD mp5  l=0.42u w=0.6u m=1
M19 N_7 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M20 N_6 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_22 D VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_22 N_6 N_4 VDD mp5  l=0.42u w=0.62u m=1
M23 N_23 N_7 N_4 VDD mp5  l=0.42u w=0.6u m=1
M24 N_23 N_5 VDD VDD mp5  l=0.42u w=0.6u m=1
M25 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M26 QN N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends dfnrn2
* SPICE INPUT		Mon Sep 24 12:19:04 2018	dfnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq1
.subckt dfnrq1 CK D VDD GND Q
M1 Q N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_38 N_3 N_9 GND mn5  l=0.5u w=0.6u m=1
M3 N_9 N_6 N_37 GND mn5  l=0.5u w=0.6u m=1
M4 N_37 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_38 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_10 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_40 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_40 N_6 N_8 GND mn5  l=0.5u w=0.6u m=1
M10 N_8 N_3 N_39 GND mn5  l=0.5u w=0.6u m=1
M11 N_39 D GND GND mn5  l=0.5u w=0.6u m=1
M12 GND N_3 N_6 GND mn5  l=0.5u w=0.6u m=1
M13 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M14 N_20 N_6 N_9 VDD mp5  l=0.42u w=0.6u m=1
M15 N_19 N_3 N_9 VDD mp5  l=0.42u w=0.62u m=1
M16 N_19 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_20 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M18 N_10 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_3 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M20 N_7 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_22 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_22 N_3 N_8 VDD mp5  l=0.42u w=0.6u m=1
M23 N_21 N_6 N_8 VDD mp5  l=0.42u w=0.62u m=1
M24 N_21 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_6 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M26 Q N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends dfnrq1
* SPICE INPUT		Mon Sep 24 12:19:14 2018	dfnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq2
.subckt dfnrq2 CK D VDD GND Q
M1 Q N_9 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_38 N_3 N_9 GND mn5  l=0.5u w=0.6u m=1
M3 N_9 N_6 N_37 GND mn5  l=0.5u w=0.6u m=1
M4 N_37 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_38 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_10 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_40 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_40 N_6 N_8 GND mn5  l=0.5u w=0.6u m=1
M10 N_8 N_3 N_39 GND mn5  l=0.5u w=0.6u m=1
M11 N_39 D GND GND mn5  l=0.5u w=0.6u m=1
M12 GND N_3 N_6 GND mn5  l=0.5u w=0.6u m=1
M13 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M14 N_20 N_6 N_9 VDD mp5  l=0.42u w=0.6u m=1
M15 N_19 N_3 N_9 VDD mp5  l=0.42u w=0.62u m=1
M16 N_19 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_20 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M18 N_10 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_3 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M20 N_7 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_22 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_22 N_3 N_8 VDD mp5  l=0.42u w=0.6u m=1
M23 N_21 N_6 N_8 VDD mp5  l=0.42u w=0.62u m=1
M24 N_21 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_6 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M26 Q N_9 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends dfnrq2
* SPICE INPUT		Mon Sep 24 12:19:23 2018	dfpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb1
.subckt dfpfb1 GND QN Q VDD SN CKN D
M1 QN N_14 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.6u m=1
M3 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_8 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_19 SN N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_11 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_20 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_12 N_11 N_20 GND mn5  l=0.5u w=0.6u m=1
M9 N_21 N_5 N_12 GND mn5  l=0.5u w=0.6u m=1
M10 GND N_12 N_19 GND mn5  l=0.5u w=0.6u m=1
M11 N_21 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_23 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M13 GND SN N_22 GND mn5  l=0.5u w=0.6u m=1
M14 N_24 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_22 N_16 N_14 GND mn5  l=0.5u w=0.6u m=1
M16 N_16 N_5 N_23 GND mn5  l=0.5u w=0.6u m=1
M17 N_24 N_11 N_16 GND mn5  l=0.5u w=0.6u m=1
M18 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_8 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_5 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_9 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_47 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 VDD N_5 N_11 VDD mp5  l=0.42u w=0.6u m=1
M24 N_45 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_46 N_11 N_12 VDD mp5  l=0.42u w=0.6u m=1
M26 N_45 N_5 N_12 VDD mp5  l=0.42u w=0.62u m=1
M27 N_9 N_12 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 QN N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_14 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M30 VDD N_14 N_48 VDD mp5  l=0.42u w=0.6u m=1
M31 N_46 N_9 VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_14 N_16 VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_48 N_5 N_16 VDD mp5  l=0.42u w=0.6u m=1
M34 N_16 N_11 N_47 VDD mp5  l=0.42u w=0.62u m=1
.ends dfpfb1
* SPICE INPUT		Mon Sep 24 12:19:32 2018	dfpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb2
.subckt dfpfb2 GND QN Q VDD SN CKN D
M1 QN N_14 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_5 CKN GND GND mn5  l=0.5u w=0.6u m=1
M3 Q N_8 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_8 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_19 SN N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_11 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_20 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_12 N_11 N_20 GND mn5  l=0.5u w=0.6u m=1
M9 N_21 N_5 N_12 GND mn5  l=0.5u w=0.6u m=1
M10 GND N_12 N_19 GND mn5  l=0.5u w=0.6u m=1
M11 N_21 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_23 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M13 GND SN N_22 GND mn5  l=0.5u w=0.6u m=1
M14 N_24 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_22 N_16 N_14 GND mn5  l=0.5u w=0.6u m=1
M16 N_16 N_5 N_23 GND mn5  l=0.5u w=0.6u m=1
M17 N_24 N_11 N_16 GND mn5  l=0.5u w=0.6u m=1
M18 Q N_8 VDD VDD mp5  l=0.42u w=1.28u m=1
M19 N_8 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_5 CKN VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_9 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_47 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 VDD N_5 N_11 VDD mp5  l=0.42u w=0.6u m=1
M24 N_45 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_46 N_11 N_12 VDD mp5  l=0.42u w=0.6u m=1
M26 N_45 N_5 N_12 VDD mp5  l=0.42u w=0.62u m=1
M27 N_9 N_12 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 QN N_14 VDD VDD mp5  l=0.42u w=1.28u m=1
M29 N_14 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M30 VDD N_14 N_48 VDD mp5  l=0.42u w=0.6u m=1
M31 N_46 N_9 VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_14 N_16 VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_48 N_5 N_16 VDD mp5  l=0.42u w=0.6u m=1
M34 N_16 N_11 N_47 VDD mp5  l=0.42u w=0.62u m=1
.ends dfpfb2
* SPICE INPUT		Mon Sep 24 12:19:41 2018	dfprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb1
.subckt dfprb1 GND QN Q VDD D SN CK
M1 QN N_14 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.6u m=1
M3 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_8 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_19 SN N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_11 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_20 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_12 N_5 N_20 GND mn5  l=0.5u w=0.6u m=1
M9 N_21 N_11 N_12 GND mn5  l=0.5u w=0.6u m=1
M10 GND N_12 N_19 GND mn5  l=0.5u w=0.6u m=1
M11 N_21 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_23 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M13 GND SN N_22 GND mn5  l=0.5u w=0.6u m=1
M14 N_24 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_22 N_16 N_14 GND mn5  l=0.5u w=0.6u m=1
M16 N_16 N_11 N_23 GND mn5  l=0.5u w=0.6u m=1
M17 N_24 N_5 N_16 GND mn5  l=0.5u w=0.6u m=1
M18 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_8 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_5 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_9 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_47 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 VDD N_5 N_11 VDD mp5  l=0.42u w=0.6u m=1
M24 N_45 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_46 N_5 N_12 VDD mp5  l=0.42u w=0.6u m=1
M26 N_45 N_11 N_12 VDD mp5  l=0.42u w=0.62u m=1
M27 N_9 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M28 QN N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 N_14 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M30 VDD N_14 N_48 VDD mp5  l=0.42u w=0.6u m=1
M31 N_46 N_9 VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_14 N_16 VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_48 N_11 N_16 VDD mp5  l=0.42u w=0.6u m=1
M34 N_16 N_5 N_47 VDD mp5  l=0.42u w=0.62u m=1
.ends dfprb1
* SPICE INPUT		Mon Sep 24 12:19:49 2018	dfprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb2
.subckt dfprb2 GND QN Q VDD D SN CK
M1 QN N_14 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_5 CK GND GND mn5  l=0.5u w=0.6u m=1
M3 Q N_8 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_8 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_19 SN N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_11 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_20 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_12 N_5 N_20 GND mn5  l=0.5u w=0.6u m=1
M9 N_21 N_11 N_12 GND mn5  l=0.5u w=0.6u m=1
M10 GND N_12 N_19 GND mn5  l=0.5u w=0.6u m=1
M11 N_21 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_23 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M13 GND SN N_22 GND mn5  l=0.5u w=0.6u m=1
M14 N_24 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_22 N_16 N_14 GND mn5  l=0.5u w=0.6u m=1
M16 N_16 N_11 N_23 GND mn5  l=0.5u w=0.6u m=1
M17 N_24 N_5 N_16 GND mn5  l=0.5u w=0.6u m=1
M18 Q N_8 VDD VDD mp5  l=0.42u w=1.28u m=1
M19 N_8 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_5 CK VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_9 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_47 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 VDD N_5 N_11 VDD mp5  l=0.42u w=0.6u m=1
M24 N_45 D VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_46 N_5 N_12 VDD mp5  l=0.42u w=0.6u m=1
M26 N_45 N_11 N_12 VDD mp5  l=0.42u w=0.62u m=1
M27 N_9 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M28 QN N_14 VDD VDD mp5  l=0.42u w=1.28u m=1
M29 N_14 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M30 VDD N_14 N_48 VDD mp5  l=0.42u w=0.6u m=1
M31 N_46 N_9 VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_14 N_16 VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_48 N_11 N_16 VDD mp5  l=0.42u w=0.6u m=1
M34 N_16 N_5 N_47 VDD mp5  l=0.42u w=0.62u m=1
.ends dfprb2
* SPICE INPUT		Mon Sep 24 12:19:58 2018	dfprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq1
.subckt dfprq1 GND Q VDD CK D SN
M1 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M2 N_17 N_14 N_5 GND mn5  l=0.5u w=0.6u m=1
M3 Q N_14 N_16 GND mn5  l=0.5u w=0.72u m=1
M4 N_17 SN GND GND mn5  l=0.5u w=0.6u m=1
M5 GND SN N_16 GND mn5  l=0.5u w=0.72u m=1
M6 N_18 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_10 N_9 N_18 GND mn5  l=0.5u w=0.6u m=1
M8 N_10 N_3 N_19 GND mn5  l=0.5u w=0.6u m=1
M9 N_19 D GND GND mn5  l=0.5u w=0.6u m=1
M10 N_9 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_20 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_14 N_3 N_20 GND mn5  l=0.5u w=0.6u m=1
M13 N_14 N_9 N_22 GND mn5  l=0.5u w=0.6u m=1
M14 N_22 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_21 N_10 N_12 GND mn5  l=0.5u w=0.6u m=1
M16 N_21 SN GND GND mn5  l=0.5u w=0.6u m=1
M17 N_43 N_5 VDD VDD mp5  l=0.42u w=0.6u m=1
M18 N_43 N_9 N_14 VDD mp5  l=0.42u w=0.6u m=1
M19 N_14 N_3 N_42 VDD mp5  l=0.42u w=0.62u m=1
M20 N_42 N_12 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_12 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_41 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M23 N_40 N_9 N_10 VDD mp5  l=0.42u w=0.62u m=1
M24 N_41 N_3 N_10 VDD mp5  l=0.42u w=0.6u m=1
M25 N_40 D VDD VDD mp5  l=0.42u w=0.62u m=1
M26 VDD N_3 N_9 VDD mp5  l=0.42u w=0.6u m=1
M27 N_5 N_14 VDD VDD mp5  l=0.42u w=0.6u m=1
M28 VDD N_14 Q VDD mp5  l=0.42u w=0.96u m=1
M29 N_5 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M30 VDD SN Q VDD mp5  l=0.42u w=0.96u m=1
M31 N_12 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_3 CK VDD VDD mp5  l=0.42u w=0.6u m=1
.ends dfprq1
* SPICE INPUT		Mon Sep 24 12:20:07 2018	dfprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq2
.subckt dfprq2 GND Q VDD CK D SN
M1 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M2 N_17 N_14 N_5 GND mn5  l=0.5u w=0.6u m=1
M3 Q N_14 N_16 GND mn5  l=0.5u w=0.98u m=1
M4 N_17 SN GND GND mn5  l=0.5u w=0.6u m=1
M5 GND SN N_16 GND mn5  l=0.5u w=0.98u m=1
M6 N_18 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_10 N_9 N_18 GND mn5  l=0.5u w=0.6u m=1
M8 N_10 N_3 N_19 GND mn5  l=0.5u w=0.6u m=1
M9 N_19 D GND GND mn5  l=0.5u w=0.6u m=1
M10 N_9 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_20 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_14 N_3 N_20 GND mn5  l=0.5u w=0.6u m=1
M13 N_14 N_9 N_22 GND mn5  l=0.5u w=0.6u m=1
M14 N_22 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_21 N_10 N_12 GND mn5  l=0.5u w=0.6u m=1
M16 N_21 SN GND GND mn5  l=0.5u w=0.6u m=1
M17 N_43 N_5 VDD VDD mp5  l=0.42u w=0.6u m=1
M18 N_43 N_9 N_14 VDD mp5  l=0.42u w=0.6u m=1
M19 N_14 N_3 N_42 VDD mp5  l=0.42u w=0.62u m=1
M20 N_42 N_12 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_12 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_41 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M23 N_40 N_9 N_10 VDD mp5  l=0.42u w=0.62u m=1
M24 N_41 N_3 N_10 VDD mp5  l=0.42u w=0.6u m=1
M25 N_40 D VDD VDD mp5  l=0.42u w=0.62u m=1
M26 VDD N_3 N_9 VDD mp5  l=0.42u w=0.6u m=1
M27 N_5 N_14 VDD VDD mp5  l=0.42u w=0.6u m=1
M28 VDD N_14 Q VDD mp5  l=0.42u w=1.28u m=1
M29 N_5 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M30 VDD SN Q VDD mp5  l=0.42u w=1.28u m=1
M31 N_12 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M32 N_3 CK VDD VDD mp5  l=0.42u w=0.6u m=1
.ends dfprq2
* SPICE INPUT		Mon Sep 24 12:20:16 2018	dl01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d0
.subckt dl01d0 A GND Y VDD
M1 GND N_5 N_2 GND mn5  l=0.5u w=0.92u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.92u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_3 N_2 GND GND mn5  l=0.5u w=0.92u m=1
M5 N_2 N_5 VDD VDD mp5  l=0.42u w=1.17u m=1
M6 N_5 A VDD VDD mp5  l=0.42u w=1.17u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_3 N_2 VDD VDD mp5  l=0.42u w=1.17u m=1
.ends dl01d0
* SPICE INPUT		Mon Sep 24 12:20:24 2018	dl01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d1
.subckt dl01d1 A VDD Y GND
M1 N_4 A GND GND mn5  l=0.5u w=0.92u m=1
M2 N_2 N_4 GND GND mn5  l=0.5u w=0.92u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_3 N_2 GND GND mn5  l=0.5u w=0.92u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_3 N_2 VDD VDD mp5  l=0.42u w=1.17u m=1
M7 N_4 A VDD VDD mp5  l=0.42u w=1.17u m=1
M8 N_2 N_4 VDD VDD mp5  l=0.42u w=1.17u m=1
.ends dl01d1
* SPICE INPUT		Mon Sep 24 12:20:33 2018	dl01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d2
.subckt dl01d2 A VDD Y GND
M1 N_4 A GND GND mn5  l=0.5u w=0.92u m=1
M2 N_2 N_4 GND GND mn5  l=0.5u w=0.92u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_3 N_2 GND GND mn5  l=0.5u w=0.92u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M6 N_3 N_2 VDD VDD mp5  l=0.42u w=1.17u m=1
M7 N_4 A VDD VDD mp5  l=0.42u w=1.17u m=1
M8 N_2 N_4 VDD VDD mp5  l=0.42u w=1.17u m=1
.ends dl01d2
* SPICE INPUT		Mon Sep 24 12:20:41 2018	dl02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d0
.subckt dl02d0 A VDD Y GND
M1 N_4 A GND GND mn5  l=0.5u w=0.92u m=1
M2 N_2 N_4 GND GND mn5  l=1u w=0.92u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_3 N_2 GND GND mn5  l=1u w=0.92u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_3 N_2 VDD VDD mp5  l=0.84u w=1.17u m=1
M7 N_4 A VDD VDD mp5  l=0.42u w=1.17u m=1
M8 N_2 N_4 VDD VDD mp5  l=0.84u w=1.17u m=1
.ends dl02d0
* SPICE INPUT		Mon Sep 24 12:20:50 2018	dl02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d1
.subckt dl02d1 A VDD Y GND
M1 N_4 A GND GND mn5  l=0.5u w=0.92u m=1
M2 N_2 N_4 GND GND mn5  l=1u w=0.92u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_3 N_2 GND GND mn5  l=1u w=0.92u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_3 N_2 VDD VDD mp5  l=0.84u w=1.17u m=1
M7 N_4 A VDD VDD mp5  l=0.42u w=1.17u m=1
M8 N_2 N_4 VDD VDD mp5  l=0.84u w=1.17u m=1
.ends dl02d1
* SPICE INPUT		Mon Sep 24 12:20:58 2018	dl02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d2
.subckt dl02d2 A VDD Y GND
M1 N_4 A GND GND mn5  l=0.5u w=0.92u m=1
M2 N_2 N_4 GND GND mn5  l=1u w=0.92u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_3 N_2 GND GND mn5  l=1u w=0.92u m=1
M5 Y N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M6 N_3 N_2 VDD VDD mp5  l=0.84u w=1.17u m=1
M7 N_4 A VDD VDD mp5  l=0.42u w=1.17u m=1
M8 N_2 N_4 VDD VDD mp5  l=0.84u w=1.17u m=1
.ends dl02d2
* SPICE INPUT		Mon Sep 24 12:53:56 2018	fillercap16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap16
.subckt fillercap16 VDD GND
M1 GND VDD GND GND mn5  l=6.58u w=0.81u m=1
M2 VDD GND VDD VDD mp5  l=6.58u w=1.07u m=1
.ends fillercap16
* SPICE INPUT		Mon Sep 24 12:54:03 2018	fillercap32
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap32
.subckt fillercap32 VDD GND
M1 GND VDD GND GND mn5  l=14.12u w=0.81u m=1
M2 VDD GND VDD VDD mp5  l=14.12u w=1.04u m=1
.ends fillercap32
* SPICE INPUT		Mon Sep 24 12:53:41 2018	fillercap4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap4
.subckt fillercap4 VDD GND
M1 GND VDD GND GND mn5  l=0.86u w=0.81u m=1
M2 VDD GND VDD VDD mp5  l=0.86u w=1.07u m=1
.ends fillercap4
* SPICE INPUT		Mon Sep 24 12:54:10 2018	fillercap64
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap64
.subckt fillercap64 VDD GND
M1 GND VDD GND GND mn5  l=29.43u w=0.81u m=1
M2 VDD GND VDD VDD mp5  l=29.43u w=1.04u m=1
.ends fillercap64
* SPICE INPUT		Mon Sep 24 12:53:48 2018	fillercap8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap8
.subckt fillercap8 GND VDD
M1 GND VDD GND GND mn5  l=2.77u w=0.81u m=1
M2 VDD GND VDD VDD mp5  l=2.77u w=1.07u m=1
.ends fillercap8
* SPICE INPUT		Mon Sep 24 12:21:07 2018	inv0d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d0
.subckt inv0d0 GND VDD A Y
M1 Y A GND GND mn5  l=0.5u w=0.6u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends inv0d0
* SPICE INPUT		Mon Sep 24 12:21:16 2018	inv0d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d1
.subckt inv0d1 GND VDD A Y
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d1
* SPICE INPUT		Mon Sep 24 12:21:27 2018	inv0d10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d10
.subckt inv0d10 A Y GND VDD
M1 Y A GND GND mn5  l=0.5u w=0.98u m=1
M2 Y A GND GND mn5  l=0.5u w=0.98u m=1
M3 Y A GND GND mn5  l=0.5u w=0.98u m=1
M4 GND A Y GND mn5  l=0.5u w=0.98u m=1
M5 Y A GND GND mn5  l=0.5u w=0.98u m=1
M6 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
M7 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
M8 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
M9 VDD A Y VDD mp5  l=0.42u w=1.28u m=1
M10 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
.ends inv0d10
* SPICE INPUT		Mon Sep 24 12:21:36 2018	inv0d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d2
.subckt inv0d2 VDD Y GND A
M1 Y A GND GND mn5  l=0.5u w=0.98u m=1
M2 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
.ends inv0d2
* SPICE INPUT		Mon Sep 24 12:21:45 2018	inv0d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d3
.subckt inv0d3 Y GND VDD A
M1 GND A Y GND mn5  l=0.5u w=0.735u m=1
M2 GND A Y GND mn5  l=0.5u w=0.735u m=1
M3 VDD A Y VDD mp5  l=0.42u w=0.96u m=1
M4 VDD A Y VDD mp5  l=0.42u w=0.96u m=1
.ends inv0d3
* SPICE INPUT		Mon Sep 24 12:21:53 2018	inv0d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d4
.subckt inv0d4 Y GND VDD A
M1 GND A Y GND mn5  l=0.5u w=0.98u m=1
M2 GND A Y GND mn5  l=0.5u w=0.98u m=1
M3 VDD A Y VDD mp5  l=0.42u w=1.28u m=1
M4 VDD A Y VDD mp5  l=0.42u w=1.28u m=1
.ends inv0d4
* SPICE INPUT		Mon Sep 24 12:22:02 2018	inv0d5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d5
.subckt inv0d5 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.9u m=1
M2 Y A GND GND mn5  l=0.5u w=0.9u m=1
M3 Y A GND GND mn5  l=0.5u w=0.65u m=1
M4 Y A VDD VDD mp5  l=0.42u w=1.1u m=1
M5 Y A VDD VDD mp5  l=0.42u w=1.1u m=1
M6 Y A VDD VDD mp5  l=0.42u w=1u m=1
.ends inv0d5
* SPICE INPUT		Mon Sep 24 12:22:11 2018	inv0d6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d6
.subckt inv0d6 GND Y VDD A
M1 Y A GND GND mn5  l=0.5u w=0.98u m=1
M2 Y A GND GND mn5  l=0.5u w=0.98u m=1
M3 Y A GND GND mn5  l=0.5u w=0.98u m=1
M4 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
M5 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
M6 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
.ends inv0d6
* SPICE INPUT		Mon Sep 24 12:22:19 2018	inv0d8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d8
.subckt inv0d8 Y GND VDD A
M1 GND A Y GND mn5  l=0.5u w=0.98u m=1
M2 GND A Y GND mn5  l=0.5u w=0.98u m=1
M3 GND A Y GND mn5  l=0.5u w=0.98u m=1
M4 Y A GND GND mn5  l=0.5u w=0.98u m=1
M5 VDD A Y VDD mp5  l=0.42u w=1.28u m=1
M6 VDD A Y VDD mp5  l=0.42u w=1.28u m=1
M7 VDD A Y VDD mp5  l=0.42u w=1.28u m=1
M8 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
.ends inv0d8
* SPICE INPUT		Mon Sep 24 12:22:28 2018	invtd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtd0
.subckt invtd0 A OE GND VDD Y
M1 N_3 OE GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_3 N_14 GND mn5  l=0.5u w=0.6u m=1
M3 GND A N_14 GND mn5  l=0.5u w=0.6u m=1
M4 N_3 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M5 Y OE N_9 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD A N_9 VDD mp5  l=0.42u w=0.62u m=1
.ends invtd0
* SPICE INPUT		Mon Sep 24 12:22:38 2018	invtd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtd1
.subckt invtd1 A OE GND VDD Y
M1 N_2 OE GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A N_14 GND mn5  l=0.5u w=0.72u m=1
M3 Y N_2 N_14 GND mn5  l=0.5u w=0.72u m=1
M4 N_2 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M5 VDD A N_9 VDD mp5  l=0.42u w=0.96u m=1
M6 Y OE N_9 VDD mp5  l=0.42u w=0.96u m=1
.ends invtd1
* SPICE INPUT		Mon Sep 24 12:22:49 2018	invtd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtd2
.subckt invtd2 A OE GND Y VDD
M1 N_3 OE GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_3 N_14 GND mn5  l=0.5u w=0.98u m=1
M3 GND A N_14 GND mn5  l=0.5u w=0.98u m=1
M4 N_3 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M5 Y OE N_9 VDD mp5  l=0.42u w=1.28u m=1
M6 VDD A N_9 VDD mp5  l=0.42u w=1.28u m=1
.ends invtd2
* SPICE INPUT		Mon Sep 24 12:22:59 2018	invtld0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld0
.subckt invtld0 A OE GND VDD Y
M1 N_5 OE GND GND mn5  l=0.5u w=0.6u m=1
M2 Y OE N_14 GND mn5  l=0.5u w=0.6u m=1
M3 GND A N_14 GND mn5  l=0.5u w=0.6u m=1
M4 N_5 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M5 Y N_5 N_9 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD A N_9 VDD mp5  l=0.42u w=0.62u m=1
.ends invtld0
* SPICE INPUT		Mon Sep 24 12:23:10 2018	invtld1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld1
.subckt invtld1 OE A GND VDD Y
M1 N_5 OE GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A N_14 GND mn5  l=0.5u w=0.72u m=1
M3 Y OE N_14 GND mn5  l=0.5u w=0.72u m=1
M4 N_5 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M5 VDD A N_9 VDD mp5  l=0.42u w=0.96u m=1
M6 Y N_5 N_9 VDD mp5  l=0.42u w=0.96u m=1
.ends invtld1
* SPICE INPUT		Mon Sep 24 12:23:19 2018	invtld2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld2
.subckt invtld2 A OE GND Y VDD
M1 N_5 OE GND GND mn5  l=0.5u w=0.6u m=1
M2 Y OE N_14 GND mn5  l=0.5u w=0.98u m=1
M3 GND A N_14 GND mn5  l=0.5u w=0.98u m=1
M4 N_5 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M5 Y N_5 N_9 VDD mp5  l=0.42u w=1.28u m=1
M6 VDD A N_9 VDD mp5  l=0.42u w=1.28u m=1
.ends invtld2
* SPICE INPUT		Mon Sep 24 12:23:28 2018	labhb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=labhb1
.subckt labhb1 RN D SN G QN VDD GND Q
M1 Q N_2 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_4 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_6 G GND GND mn5  l=0.5u w=0.6u m=1
M4 N_7 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_3 SN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_21 D GND GND mn5  l=0.5u w=0.6u m=1
M7 N_22 RN N_21 GND mn5  l=0.5u w=0.6u m=1
M8 N_2 N_7 N_22 GND mn5  l=0.5u w=0.6u m=1
M9 N_23 N_6 N_2 GND mn5  l=0.5u w=0.6u m=1
M10 N_24 RN N_23 GND mn5  l=0.5u w=0.6u m=1
M11 N_24 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_4 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_4 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 VDD SN N_3 VDD mp5  l=0.42u w=0.62u m=1
M16 N_40 D VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_2 N_6 N_41 VDD mp5  l=0.42u w=0.62u m=1
M18 N_42 N_7 N_2 VDD mp5  l=0.42u w=0.62u m=1
M19 N_43 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 VDD RN N_39 VDD mp5  l=0.42u w=0.62u m=1
M21 N_2 N_3 N_39 VDD mp5  l=0.42u w=0.62u m=1
M22 N_41 N_3 N_40 VDD mp5  l=0.42u w=0.62u m=1
M23 N_43 N_3 N_42 VDD mp5  l=0.42u w=0.62u m=1
M24 N_6 G VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_7 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M26 Q N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M27 QN N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends labhb1
* SPICE INPUT		Mon Sep 24 12:23:37 2018	labhb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=labhb2
.subckt labhb2 GND QN Q VDD G SN D RN
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M3 N_6 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_9 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_18 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_18 RN N_17 GND mn5  l=0.5u w=0.6u m=1
M7 N_17 N_4 N_9 GND mn5  l=0.5u w=0.6u m=1
M8 N_9 N_3 N_16 GND mn5  l=0.5u w=0.6u m=1
M9 N_16 RN N_15 GND mn5  l=0.5u w=0.6u m=1
M10 N_15 D GND GND mn5  l=0.5u w=0.6u m=1
M11 N_8 SN GND GND mn5  l=0.5u w=0.6u m=1
M12 QN N_6 GND GND mn5  l=0.5u w=0.98u m=1
M13 Q N_9 GND GND mn5  l=0.5u w=0.98u m=1
M14 N_6 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_9 N_8 N_38 VDD mp5  l=0.42u w=0.62u m=1
M16 N_40 N_8 N_39 VDD mp5  l=0.42u w=0.62u m=1
M17 N_42 N_8 N_41 VDD mp5  l=0.42u w=0.62u m=1
M18 VDD RN N_38 VDD mp5  l=0.42u w=0.62u m=1
M19 N_42 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_41 N_3 N_9 VDD mp5  l=0.42u w=0.62u m=1
M21 N_9 N_4 N_40 VDD mp5  l=0.42u w=0.62u m=1
M22 N_39 D VDD VDD mp5  l=0.42u w=0.62u m=1
M23 VDD SN N_8 VDD mp5  l=0.42u w=0.62u m=1
M24 QN N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M25 Q N_9 VDD VDD mp5  l=0.42u w=1.28u m=1
M26 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M27 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
.ends labhb2
* SPICE INPUT		Mon Sep 24 12:23:46 2018	lablb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb1
.subckt lablb1 GND QN Q VDD RN D SN GN
M1 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_12 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_7 GN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_11 SN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_15 D GND GND mn5  l=0.5u w=0.6u m=1
M7 N_16 RN N_15 GND mn5  l=0.5u w=0.6u m=1
M8 N_12 N_7 N_16 GND mn5  l=0.5u w=0.6u m=1
M9 N_9 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_17 N_6 N_12 GND mn5  l=0.5u w=0.6u m=1
M11 N_18 RN N_17 GND mn5  l=0.5u w=0.6u m=1
M12 N_18 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_12 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_7 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_6 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M17 Q N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M18 N_9 N_12 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 VDD SN N_11 VDD mp5  l=0.42u w=0.62u m=1
M20 N_39 D VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_12 N_6 N_40 VDD mp5  l=0.42u w=0.62u m=1
M22 N_41 N_7 N_12 VDD mp5  l=0.42u w=0.62u m=1
M23 N_42 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M24 VDD RN N_38 VDD mp5  l=0.42u w=0.62u m=1
M25 N_12 N_11 N_38 VDD mp5  l=0.42u w=0.62u m=1
M26 N_40 N_11 N_39 VDD mp5  l=0.42u w=0.62u m=1
M27 N_42 N_11 N_41 VDD mp5  l=0.42u w=0.62u m=1
.ends lablb1
* SPICE INPUT		Mon Sep 24 12:23:55 2018	lablb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb2
.subckt lablb2 GND QN Q VDD RN D SN GN
M1 N_4 GN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_8 SN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_15 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_16 RN N_15 GND mn5  l=0.5u w=0.6u m=1
M6 N_9 N_4 N_16 GND mn5  l=0.5u w=0.6u m=1
M7 N_6 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_17 N_3 N_9 GND mn5  l=0.5u w=0.6u m=1
M9 N_18 RN N_17 GND mn5  l=0.5u w=0.6u m=1
M10 N_18 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_9 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M12 QN N_6 GND GND mn5  l=0.5u w=0.98u m=1
M13 Q N_9 GND GND mn5  l=0.5u w=0.98u m=1
M14 N_4 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 QN N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M17 Q N_9 VDD VDD mp5  l=0.42u w=1.28u m=1
M18 N_6 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 VDD SN N_8 VDD mp5  l=0.42u w=0.62u m=1
M20 N_39 D VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_9 N_3 N_40 VDD mp5  l=0.42u w=0.62u m=1
M22 N_41 N_4 N_9 VDD mp5  l=0.42u w=0.62u m=1
M23 N_42 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M24 VDD RN N_38 VDD mp5  l=0.42u w=0.62u m=1
M25 N_9 N_8 N_38 VDD mp5  l=0.42u w=0.62u m=1
M26 N_40 N_8 N_39 VDD mp5  l=0.42u w=0.62u m=1
M27 N_42 N_8 N_41 VDD mp5  l=0.42u w=0.62u m=1
.ends lablb2
* SPICE INPUT		Mon Sep 24 12:24:03 2018	lachb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb1
.subckt lachb1 GND QN Q VDD RN D G
M1 Q N_11 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_7 G GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_13 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_14 RN N_13 GND mn5  l=0.5u w=0.6u m=1
M7 N_11 N_6 N_14 GND mn5  l=0.5u w=0.6u m=1
M8 N_15 N_7 N_11 GND mn5  l=0.5u w=0.6u m=1
M9 N_16 RN N_15 GND mn5  l=0.5u w=0.6u m=1
M10 N_16 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_9 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_7 G VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_6 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_9 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 Q N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 QN N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M17 N_34 D VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_11 N_7 N_34 VDD mp5  l=0.42u w=0.62u m=1
M19 N_35 N_6 N_11 VDD mp5  l=0.42u w=0.62u m=1
M20 N_11 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_35 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lachb1
* SPICE INPUT		Mon Sep 24 12:24:12 2018	lachb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb2
.subckt lachb2 GND QN Q VDD D RN G
M1 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_13 D GND GND mn5  l=0.5u w=0.6u m=1
M4 N_14 RN N_13 GND mn5  l=0.5u w=0.6u m=1
M5 N_8 N_3 N_14 GND mn5  l=0.5u w=0.6u m=1
M6 N_15 N_4 N_8 GND mn5  l=0.5u w=0.6u m=1
M7 N_16 RN N_15 GND mn5  l=0.5u w=0.6u m=1
M8 N_16 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_6 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M10 Q N_8 GND GND mn5  l=0.5u w=0.98u m=1
M11 QN N_6 GND GND mn5  l=0.5u w=0.98u m=1
M12 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_6 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 Q N_8 VDD VDD mp5  l=0.42u w=1.28u m=1
M16 QN N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M17 N_34 D VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_8 N_4 N_34 VDD mp5  l=0.42u w=0.62u m=1
M19 N_35 N_3 N_8 VDD mp5  l=0.42u w=0.62u m=1
M20 N_8 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_35 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lachb2
* SPICE INPUT		Mon Sep 24 12:24:20 2018	lachq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachq1
.subckt lachq1 GND Q VDD D RN G
M1 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 D GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 RN N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_8 N_3 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_4 N_8 GND mn5  l=0.5u w=0.6u m=1
M7 N_15 RN N_14 GND mn5  l=0.5u w=0.6u m=1
M8 N_15 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_6 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M10 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_6 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M15 N_32 D VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_8 N_4 N_32 VDD mp5  l=0.42u w=0.62u m=1
M17 N_33 N_3 N_8 VDD mp5  l=0.42u w=0.62u m=1
M18 N_8 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_33 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lachq1
* SPICE INPUT		Mon Sep 24 12:24:30 2018	lachq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachq2
.subckt lachq2 GND Q VDD D RN G
M1 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 D GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 RN N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_8 N_3 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_4 N_8 GND mn5  l=0.5u w=0.6u m=1
M7 N_15 RN N_14 GND mn5  l=0.5u w=0.6u m=1
M8 N_15 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_6 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M10 Q N_8 GND GND mn5  l=0.5u w=0.98u m=1
M11 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_6 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 Q N_8 VDD VDD mp5  l=0.42u w=1.28u m=1
M15 N_32 D VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_8 N_4 N_32 VDD mp5  l=0.42u w=0.62u m=1
M17 N_33 N_3 N_8 VDD mp5  l=0.42u w=0.62u m=1
M18 N_8 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_33 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lachq2
* SPICE INPUT		Mon Sep 24 12:24:38 2018	laclb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb1
.subckt laclb1 RN D GN Q QN VDD GND
M1 Q N_8 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_2 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_4 GN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_31 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_32 RN N_31 GND mn5  l=0.5u w=0.6u m=1
M7 N_8 N_4 N_32 GND mn5  l=0.5u w=0.6u m=1
M8 N_33 N_5 N_8 GND mn5  l=0.5u w=0.6u m=1
M9 N_34 RN N_33 GND mn5  l=0.5u w=0.6u m=1
M10 N_34 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_2 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_4 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_2 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 Q N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 QN N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M17 N_18 D VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_8 N_5 N_18 VDD mp5  l=0.42u w=0.62u m=1
M19 N_19 N_4 N_8 VDD mp5  l=0.42u w=0.62u m=1
M20 N_8 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_19 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends laclb1
* SPICE INPUT		Mon Sep 24 12:24:47 2018	laclb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb2
.subckt laclb2 RN D GN QN Q VDD GND
M1 N_4 GN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_18 D GND GND mn5  l=0.5u w=0.6u m=1
M4 N_19 RN N_18 GND mn5  l=0.5u w=0.6u m=1
M5 N_8 N_4 N_19 GND mn5  l=0.5u w=0.6u m=1
M6 N_20 N_5 N_8 GND mn5  l=0.5u w=0.6u m=1
M7 N_21 RN N_20 GND mn5  l=0.5u w=0.6u m=1
M8 N_21 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_2 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M10 Q N_8 GND GND mn5  l=0.5u w=0.98u m=1
M11 QN N_2 GND GND mn5  l=0.5u w=0.98u m=1
M12 N_4 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_2 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 Q N_8 VDD VDD mp5  l=0.42u w=1.28u m=1
M16 QN N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
M17 N_35 D VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_8 N_5 N_35 VDD mp5  l=0.42u w=0.62u m=1
M19 N_36 N_4 N_8 VDD mp5  l=0.42u w=0.62u m=1
M20 N_8 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_36 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends laclb2
* SPICE INPUT		Mon Sep 24 12:24:56 2018	laclq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclq1
.subckt laclq1 VDD Q GND RN D GN
M1 Q N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 GN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_30 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_31 RN N_30 GND mn5  l=0.5u w=0.6u m=1
M6 N_6 N_4 N_31 GND mn5  l=0.5u w=0.6u m=1
M7 N_32 N_3 N_6 GND mn5  l=0.5u w=0.6u m=1
M8 N_33 RN N_32 GND mn5  l=0.5u w=0.6u m=1
M9 N_33 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_10 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_4 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_14 D VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_6 N_3 N_14 VDD mp5  l=0.42u w=0.62u m=1
M15 N_15 N_4 N_6 VDD mp5  l=0.42u w=0.62u m=1
M16 N_6 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_15 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_10 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 Q N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends laclq1
* SPICE INPUT		Mon Sep 24 12:25:07 2018	laclq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclq2
.subckt laclq2 RN D GN GND VDD Q
M1 Q N_7 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_4 GN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_28 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_29 RN N_28 GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_4 N_29 GND mn5  l=0.5u w=0.6u m=1
M7 N_30 N_5 N_7 GND mn5  l=0.5u w=0.6u m=1
M8 N_31 RN N_30 GND mn5  l=0.5u w=0.6u m=1
M9 N_31 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_2 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_4 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 Q N_7 VDD VDD mp5  l=0.42u w=1.28u m=1
M15 N_16 D VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_7 N_5 N_16 VDD mp5  l=0.42u w=0.62u m=1
M17 N_17 N_4 N_7 VDD mp5  l=0.42u w=0.62u m=1
M18 N_7 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_17 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends laclq2
* SPICE INPUT		Mon Sep 24 12:25:17 2018	lanhb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb1
.subckt lanhb1 D G VDD QN Q GND
M1 Q N_2 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_15 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_2 N_5 N_15 GND mn5  l=0.5u w=0.6u m=1
M7 N_16 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M8 N_16 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M10 Q N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 QN N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_28 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_4 N_28 VDD mp5  l=0.42u w=0.62u m=1
M14 N_29 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M15 N_29 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanhb1
* SPICE INPUT		Mon Sep 24 12:25:27 2018	lanhb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb2
.subckt lanhb2 GND QN Q VDD D G
M1 Q N_11 GND GND mn5  l=0.5u w=0.98u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_6 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_7 G GND GND mn5  l=0.5u w=0.6u m=1
M5 N_13 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_11 N_6 N_13 GND mn5  l=0.5u w=0.6u m=1
M7 N_14 N_7 N_11 GND mn5  l=0.5u w=0.6u m=1
M8 N_14 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_9 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M10 Q N_11 VDD VDD mp5  l=0.42u w=1.28u m=1
M11 QN N_9 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 N_29 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_11 N_7 N_29 VDD mp5  l=0.42u w=0.62u m=1
M14 N_30 N_6 N_11 VDD mp5  l=0.42u w=0.62u m=1
M15 N_30 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_9 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_6 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_7 G VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanhb2
* SPICE INPUT		Mon Sep 24 12:25:35 2018	lanhn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhn1
.subckt lanhn1 D G GND VDD QN
M1 QN N_3 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_14 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_5 N_14 GND mn5  l=0.5u w=0.6u m=1
M6 N_15 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_15 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 QN N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_26 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_4 N_26 VDD mp5  l=0.42u w=0.62u m=1
M14 N_27 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M15 N_27 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanhn1
* SPICE INPUT		Mon Sep 24 12:25:44 2018	lanhn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhn2
.subckt lanhn2 D G GND QN VDD
M1 QN N_3 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_14 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_5 N_14 GND mn5  l=0.5u w=0.6u m=1
M6 N_15 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_15 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 QN N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 N_26 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_4 N_26 VDD mp5  l=0.42u w=0.62u m=1
M14 N_27 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M15 N_27 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanhn2
* SPICE INPUT		Mon Sep 24 12:25:52 2018	lanhq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhq1
.subckt lanhq1 D G GND VDD Q
M1 Q N_2 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_5 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_14 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 Q N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_4 N_25 VDD mp5  l=0.42u w=0.62u m=1
M14 N_26 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M15 N_26 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanhq1
* SPICE INPUT		Mon Sep 24 12:26:01 2018	lanhq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhq2
.subckt lanhq2 D G GND VDD Q
M1 Q N_2 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_5 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_14 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_5 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 Q N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_4 N_25 VDD mp5  l=0.42u w=0.62u m=1
M14 N_26 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M15 N_26 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanhq2
* SPICE INPUT		Mon Sep 24 12:26:10 2018	lanht1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanht1
.subckt lanht1 GND VDD D G OE Q
M1 GND N_12 N_14 GND mn5  l=0.5u w=0.72u m=1
M2 Q OE N_14 GND mn5  l=0.5u w=0.72u m=1
M3 N_10 OE GND GND mn5  l=0.5u w=0.6u m=1
M4 N_9 G GND GND mn5  l=0.5u w=0.6u m=1
M5 N_8 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M6 GND N_12 N_13 GND mn5  l=0.5u w=0.6u m=1
M7 N_31 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_31 N_9 N_12 GND mn5  l=0.5u w=0.6u m=1
M9 N_12 N_8 N_30 GND mn5  l=0.5u w=0.6u m=1
M10 N_30 D GND GND mn5  l=0.5u w=0.6u m=1
M11 N_13 N_12 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_29 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_29 N_8 N_12 VDD mp5  l=0.42u w=0.62u m=1
M14 N_28 D VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_12 N_9 N_28 VDD mp5  l=0.42u w=0.62u m=1
M16 N_10 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M17 VDD N_12 N_14 VDD mp5  l=0.42u w=0.96u m=1
M18 Q N_10 N_14 VDD mp5  l=0.42u w=0.96u m=1
M19 N_9 G VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_8 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanht1
* SPICE INPUT		Mon Sep 24 12:26:18 2018	lanht2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanht2
.subckt lanht2 GND VDD D G OE Q
M1 GND N_12 N_14 GND mn5  l=0.5u w=0.98u m=1
M2 Q OE N_14 GND mn5  l=0.5u w=0.98u m=1
M3 N_10 OE GND GND mn5  l=0.5u w=0.6u m=1
M4 N_9 G GND GND mn5  l=0.5u w=0.6u m=1
M5 N_8 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M6 GND N_12 N_13 GND mn5  l=0.5u w=0.6u m=1
M7 N_31 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_31 N_9 N_12 GND mn5  l=0.5u w=0.6u m=1
M9 N_12 N_8 N_30 GND mn5  l=0.5u w=0.6u m=1
M10 N_30 D GND GND mn5  l=0.5u w=0.6u m=1
M11 N_13 N_12 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_29 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_29 N_8 N_12 VDD mp5  l=0.42u w=0.62u m=1
M14 N_28 D VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_12 N_9 N_28 VDD mp5  l=0.42u w=0.62u m=1
M16 N_10 OE VDD VDD mp5  l=0.42u w=0.62u m=1
M17 VDD N_12 N_14 VDD mp5  l=0.42u w=1.28u m=1
M18 Q N_10 N_14 VDD mp5  l=0.42u w=1.28u m=1
M19 N_9 G VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_8 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanht2
* SPICE INPUT		Mon Sep 24 12:26:27 2018	lanlb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb1
.subckt lanlb1 D GN GND QN Q VDD
M1 Q N_2 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_5 GN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_4 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_15 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_2 N_5 N_15 GND mn5  l=0.5u w=0.6u m=1
M7 N_16 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M8 N_16 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_5 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_4 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Q N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 QN N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_28 D VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_2 N_4 N_28 VDD mp5  l=0.42u w=0.62u m=1
M16 N_29 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M17 N_29 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanlb1
* SPICE INPUT		Mon Sep 24 12:26:35 2018	lanlb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb2
.subckt lanlb2 GND QN Q VDD D GN
M1 Q N_11 GND GND mn5  l=0.5u w=0.98u m=1
M2 QN N_9 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_7 GN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_13 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_11 N_7 N_13 GND mn5  l=0.5u w=0.6u m=1
M7 N_14 N_6 N_11 GND mn5  l=0.5u w=0.6u m=1
M8 N_14 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_9 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_7 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_6 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Q N_11 VDD VDD mp5  l=0.42u w=1.28u m=1
M13 QN N_9 VDD VDD mp5  l=0.42u w=1.28u m=1
M14 N_29 D VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_11 N_6 N_29 VDD mp5  l=0.42u w=0.62u m=1
M16 N_30 N_7 N_11 VDD mp5  l=0.42u w=0.62u m=1
M17 N_30 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_9 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanlb2
* SPICE INPUT		Mon Sep 24 12:26:43 2018	lanln1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanln1
.subckt lanln1 D GN GND VDD QN
M1 QN N_3 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_5 GN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_4 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_14 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_5 N_14 GND mn5  l=0.5u w=0.6u m=1
M6 N_15 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_15 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_5 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_4 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 QN N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_26 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_4 N_26 VDD mp5  l=0.42u w=0.62u m=1
M14 N_27 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M15 N_27 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanln1
* SPICE INPUT		Mon Sep 24 12:26:51 2018	lanln2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanln2
.subckt lanln2 D GN GND VDD QN
M1 QN N_3 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_5 GN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_4 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_14 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_5 N_14 GND mn5  l=0.5u w=0.6u m=1
M6 N_15 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_15 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_5 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_4 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 QN N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 N_26 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_4 N_26 VDD mp5  l=0.42u w=0.62u m=1
M14 N_27 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M15 N_27 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanln2
* SPICE INPUT		Mon Sep 24 12:26:59 2018	lanlq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlq1
.subckt lanlq1 D GN GND Q VDD
M1 Q N_2 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_5 GN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_4 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_5 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_14 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_5 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_4 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 Q N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_4 N_25 VDD mp5  l=0.42u w=0.62u m=1
M14 N_26 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M15 N_26 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanlq1
* SPICE INPUT		Mon Sep 24 12:27:07 2018	lanlq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlq2
.subckt lanlq2 D GN VDD Q GND
M1 Q N_2 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_5 GN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_4 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_5 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_14 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_3 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_5 GN VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_4 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 Q N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_2 N_4 N_25 VDD mp5  l=0.42u w=0.62u m=1
M14 N_26 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M15 N_26 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_3 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends lanlq2
* SPICE INPUT		Mon Sep 24 12:27:16 2018	laphb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb1
.subckt laphb1 GND QN Q VDD D SN G
M1 N_4 G GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_8 SN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_16 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_6 N_3 N_16 GND mn5  l=0.5u w=0.6u m=1
M6 N_17 N_4 N_6 GND mn5  l=0.5u w=0.6u m=1
M7 N_6 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_17 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M9 Q N_6 GND GND mn5  l=0.5u w=0.72u m=1
M10 QN N_14 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_14 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_4 G VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_14 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 VDD SN N_8 VDD mp5  l=0.42u w=0.62u m=1
M16 N_35 D VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_6 N_4 N_36 VDD mp5  l=0.42u w=0.62u m=1
M18 N_37 N_3 N_6 VDD mp5  l=0.42u w=0.62u m=1
M19 N_36 N_8 N_35 VDD mp5  l=0.42u w=0.62u m=1
M20 N_38 N_8 N_37 VDD mp5  l=0.42u w=0.62u m=1
M21 N_38 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 Q N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M23 QN N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends laphb1
* SPICE INPUT		Mon Sep 24 12:27:24 2018	laphb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb2
.subckt laphb2 GND QN Q VDD D G SN
M1 Q N_11 GND GND mn5  l=0.5u w=0.98u m=1
M2 QN N_6 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_6 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_8 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_9 G GND GND mn5  l=0.5u w=0.6u m=1
M6 N_13 SN GND GND mn5  l=0.5u w=0.6u m=1
M7 N_16 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_17 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_11 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_17 N_9 N_11 GND mn5  l=0.5u w=0.6u m=1
M11 N_11 N_8 N_16 GND mn5  l=0.5u w=0.6u m=1
M12 Q N_11 VDD VDD mp5  l=0.42u w=1.28u m=1
M13 QN N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M14 VDD SN N_13 VDD mp5  l=0.42u w=0.62u m=1
M15 N_6 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_35 D VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_38 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_36 N_13 N_35 VDD mp5  l=0.42u w=0.62u m=1
M19 N_38 N_13 N_37 VDD mp5  l=0.42u w=0.62u m=1
M20 N_37 N_8 N_11 VDD mp5  l=0.42u w=0.62u m=1
M21 N_11 N_9 N_36 VDD mp5  l=0.42u w=0.62u m=1
M22 N_8 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_9 G VDD VDD mp5  l=0.42u w=0.62u m=1
.ends laphb2
* SPICE INPUT		Mon Sep 24 12:27:32 2018	laplb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb1
.subckt laplb1 GND QN Q VDD GN SN D
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_4 GN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_17 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_17 N_3 N_6 GND mn5  l=0.5u w=0.6u m=1
M6 N_6 N_4 N_16 GND mn5  l=0.5u w=0.6u m=1
M7 N_16 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_8 SN GND GND mn5  l=0.5u w=0.6u m=1
M9 QN N_14 GND GND mn5  l=0.5u w=0.72u m=1
M10 Q N_6 GND GND mn5  l=0.5u w=0.72u m=1
M11 N_14 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_14 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_38 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_36 N_8 N_35 VDD mp5  l=0.42u w=0.62u m=1
M15 N_38 N_8 N_37 VDD mp5  l=0.42u w=0.62u m=1
M16 N_37 N_4 N_6 VDD mp5  l=0.42u w=0.62u m=1
M17 N_6 N_3 N_36 VDD mp5  l=0.42u w=0.62u m=1
M18 N_35 D VDD VDD mp5  l=0.42u w=0.62u m=1
M19 VDD SN N_8 VDD mp5  l=0.42u w=0.62u m=1
M20 QN N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M21 Q N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M22 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_4 GN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends laplb1
* SPICE INPUT		Mon Sep 24 12:27:43 2018	laplb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb2
.subckt laplb2 GND QN Q VDD GN SN D
M1 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_4 GN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_17 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_17 N_3 N_6 GND mn5  l=0.5u w=0.6u m=1
M6 N_6 N_4 N_16 GND mn5  l=0.5u w=0.6u m=1
M7 N_16 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_8 SN GND GND mn5  l=0.5u w=0.6u m=1
M9 QN N_14 GND GND mn5  l=0.5u w=0.98u m=1
M10 Q N_6 GND GND mn5  l=0.5u w=0.98u m=1
M11 N_14 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_14 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_38 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_36 N_8 N_35 VDD mp5  l=0.42u w=0.62u m=1
M15 N_38 N_8 N_37 VDD mp5  l=0.42u w=0.62u m=1
M16 N_37 N_4 N_6 VDD mp5  l=0.42u w=0.62u m=1
M17 N_6 N_3 N_36 VDD mp5  l=0.42u w=0.62u m=1
M18 N_35 D VDD VDD mp5  l=0.42u w=0.62u m=1
M19 VDD SN N_8 VDD mp5  l=0.42u w=0.62u m=1
M20 QN N_14 VDD VDD mp5  l=0.42u w=1.28u m=1
M21 Q N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M22 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_4 GN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends laplb2
* SPICE INPUT		Mon Sep 24 12:27:52 2018	mi02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d0
.subckt mi02d0 S0 B A GND VDD Y
M1 N_12 A GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 S0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_10 B GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 S0 Y GND mn5  l=0.5u w=0.6u m=1
M6 N_12 A VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_10 B VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y S0 N_12 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_3 N_10 VDD mp5  l=0.42u w=0.62u m=1
.ends mi02d0
* SPICE INPUT		Mon Sep 24 12:28:01 2018	mi02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d1
.subckt mi02d1 S0 B A VDD Y GND
M1 N_11 A GND GND mn5  l=0.5u w=0.6u m=1
M2 Y S0 N_9 GND mn5  l=0.5u w=0.72u m=1
M3 N_9 B GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 N_11 GND mn5  l=0.5u w=0.72u m=1
M5 N_3 S0 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_11 A VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y S0 N_11 VDD mp5  l=0.42u w=0.96u m=1
M8 N_9 B VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_3 N_9 VDD mp5  l=0.42u w=0.96u m=1
M10 N_3 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends mi02d1
* SPICE INPUT		Mon Sep 24 12:28:10 2018	mi02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d2
.subckt mi02d2 S0 B A VDD Y GND
M1 N_11 A GND GND mn5  l=0.5u w=0.6u m=1
M2 Y S0 N_9 GND mn5  l=0.5u w=0.98u m=1
M3 N_9 B GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 N_11 GND mn5  l=0.5u w=0.98u m=1
M5 N_3 S0 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_11 A VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y S0 N_11 VDD mp5  l=0.42u w=1.28u m=1
M8 N_9 B VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_3 N_9 VDD mp5  l=0.42u w=1.28u m=1
M10 N_3 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends mi02d2
* SPICE INPUT		Mon Sep 24 12:28:19 2018	mi04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi04d0
.subckt mi04d0 VDD Y GND D B A S0 S1 C
M1 N_10 N_8 N_11 GND mn5  l=0.5u w=0.6u m=1
M2 GND D N_12 GND mn5  l=0.5u w=0.6u m=1
M3 N_8 S0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 B GND GND mn5  l=0.5u w=0.6u m=1
M5 N_17 S1 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_20 N_13 GND mn5  l=0.5u w=0.6u m=1
M7 N_17 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_3 A GND GND mn5  l=0.5u w=0.6u m=1
M9 N_3 N_8 N_6 GND mn5  l=0.5u w=0.6u m=1
M10 N_6 S0 N_5 GND mn5  l=0.5u w=0.6u m=1
M11 N_11 C GND GND mn5  l=0.5u w=0.6u m=1
M12 N_14 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_10 S0 N_12 GND mn5  l=0.5u w=0.6u m=1
M14 N_20 S1 GND GND mn5  l=0.5u w=0.6u m=1
M15 Y N_13 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_5 B VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_3 A VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_6 N_8 N_5 VDD mp5  l=0.42u w=0.62u m=1
M19 N_6 S0 N_3 VDD mp5  l=0.42u w=0.62u m=1
M20 N_12 D VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_8 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_11 C VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_12 N_8 N_10 VDD mp5  l=0.42u w=0.62u m=1
M24 N_11 S0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M25 N_14 S1 N_13 VDD mp5  l=0.42u w=0.62u m=1
M26 N_17 N_20 N_13 VDD mp5  l=0.42u w=0.62u m=1
M27 N_17 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_14 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_20 S1 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 Y N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends mi04d0
* SPICE INPUT		Mon Sep 24 12:28:26 2018	mi04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi04d1
.subckt mi04d1 S1 S0 C A B D GND Y VDD
M1 N_10 N_8 N_25 GND mn5  l=0.5u w=0.6u m=1
M2 GND D N_21 GND mn5  l=0.5u w=0.6u m=1
M3 N_8 S0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_22 B GND GND mn5  l=0.5u w=0.6u m=1
M5 N_26 S1 N_2 GND mn5  l=0.5u w=0.6u m=1
M6 N_23 N_11 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_26 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_19 A GND GND mn5  l=0.5u w=0.6u m=1
M9 N_19 N_8 N_5 GND mn5  l=0.5u w=0.6u m=1
M10 N_5 S0 N_22 GND mn5  l=0.5u w=0.6u m=1
M11 N_25 C GND GND mn5  l=0.5u w=0.6u m=1
M12 N_23 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_10 S0 N_21 GND mn5  l=0.5u w=0.6u m=1
M14 N_11 S1 GND GND mn5  l=0.5u w=0.6u m=1
M15 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M16 N_22 B VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_19 A VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_5 N_8 N_22 VDD mp5  l=0.42u w=0.62u m=1
M19 N_5 S0 N_19 VDD mp5  l=0.42u w=0.62u m=1
M20 N_21 D VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_8 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_25 C VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_21 N_8 N_10 VDD mp5  l=0.42u w=0.62u m=1
M24 N_25 S0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M25 N_23 S1 N_2 VDD mp5  l=0.42u w=0.62u m=1
M26 N_26 N_11 N_2 VDD mp5  l=0.42u w=0.62u m=1
M27 N_26 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_23 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_11 S1 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends mi04d1
* SPICE INPUT		Mon Sep 24 12:28:34 2018	mi04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi04d2
.subckt mi04d2 S1 S0 C A B D GND Y VDD
M1 N_10 N_8 N_25 GND mn5  l=0.5u w=0.6u m=1
M2 GND D N_21 GND mn5  l=0.5u w=0.6u m=1
M3 N_8 S0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_22 B GND GND mn5  l=0.5u w=0.6u m=1
M5 N_26 S1 N_2 GND mn5  l=0.5u w=0.6u m=1
M6 N_23 N_11 N_2 GND mn5  l=0.5u w=0.6u m=1
M7 N_26 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_19 A GND GND mn5  l=0.5u w=0.6u m=1
M9 N_19 N_8 N_5 GND mn5  l=0.5u w=0.6u m=1
M10 N_5 S0 N_22 GND mn5  l=0.5u w=0.6u m=1
M11 N_25 C GND GND mn5  l=0.5u w=0.6u m=1
M12 N_23 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_10 S0 N_21 GND mn5  l=0.5u w=0.6u m=1
M14 N_11 S1 GND GND mn5  l=0.5u w=0.6u m=1
M15 Y N_2 GND GND mn5  l=0.5u w=0.98u m=1
M16 N_22 B VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_19 A VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_5 N_8 N_22 VDD mp5  l=0.42u w=0.62u m=1
M19 N_5 S0 N_19 VDD mp5  l=0.42u w=0.62u m=1
M20 N_21 D VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_8 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_25 C VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_21 N_8 N_10 VDD mp5  l=0.42u w=0.62u m=1
M24 N_25 S0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M25 N_23 S1 N_2 VDD mp5  l=0.42u w=0.62u m=1
M26 N_26 N_11 N_2 VDD mp5  l=0.42u w=0.62u m=1
M27 N_26 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_23 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_11 S1 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 Y N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends mi04d2
* SPICE INPUT		Mon Sep 24 12:28:42 2018	mx02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d0
.subckt mx02d0 S0 A B GND VDD Y
M1 N_11 S0 N_5 GND mn5  l=0.5u w=0.6u m=1
M2 N_11 B GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_12 A GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 S0 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_5 N_2 N_12 GND mn5  l=0.5u w=0.6u m=1
M7 N_11 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_12 A VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_2 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_5 S0 N_12 VDD mp5  l=0.42u w=0.62u m=1
M12 N_11 N_2 N_5 VDD mp5  l=0.42u w=0.62u m=1
.ends mx02d0
* SPICE INPUT		Mon Sep 24 12:28:50 2018	mx02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d1
.subckt mx02d1 B S0 A GND Y VDD
M1 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_11 A GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 S0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_10 S0 N_7 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 B GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_2 N_11 GND mn5  l=0.5u w=0.6u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_11 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_2 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_7 S0 N_11 VDD mp5  l=0.42u w=0.62u m=1
M11 N_10 B VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_10 N_2 N_7 VDD mp5  l=0.42u w=0.62u m=1
.ends mx02d1
* SPICE INPUT		Mon Sep 24 12:28:58 2018	mx02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d2
.subckt mx02d2 B S0 A GND Y VDD
M1 Y N_7 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_10 A GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 S0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 S0 N_7 GND mn5  l=0.5u w=0.6u m=1
M5 N_13 B GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_2 N_10 GND mn5  l=0.5u w=0.6u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 N_10 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_2 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_7 S0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M11 N_13 B VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_13 N_2 N_7 VDD mp5  l=0.42u w=0.62u m=1
.ends mx02d2
* SPICE INPUT		Mon Sep 24 12:29:06 2018	mx04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d0
.subckt mx04d0 S0 A B D C S1 GND VDD Y
M1 N_20 N_13 N_12 GND mn5  l=0.5u w=0.6u m=1
M2 N_23 S1 N_12 GND mn5  l=0.5u w=0.6u m=1
M3 Y N_12 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 S1 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_25 C GND GND mn5  l=0.5u w=0.6u m=1
M6 N_23 N_5 N_25 GND mn5  l=0.5u w=0.6u m=1
M7 GND D N_24 GND mn5  l=0.5u w=0.6u m=1
M8 N_22 B GND GND mn5  l=0.5u w=0.6u m=1
M9 N_20 S0 N_22 GND mn5  l=0.5u w=0.6u m=1
M10 N_20 N_5 N_21 GND mn5  l=0.5u w=0.6u m=1
M11 N_21 A GND GND mn5  l=0.5u w=0.6u m=1
M12 N_23 S0 N_24 GND mn5  l=0.5u w=0.6u m=1
M13 N_5 S0 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_25 C VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_24 N_5 N_23 VDD mp5  l=0.42u w=0.6u m=1
M16 N_24 D VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_23 S0 N_25 VDD mp5  l=0.42u w=0.6u m=1
M18 N_5 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_22 B VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_20 N_5 N_22 VDD mp5  l=0.42u w=0.6u m=1
M21 N_20 S0 N_21 VDD mp5  l=0.42u w=0.6u m=1
M22 N_21 A VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.6u m=1
M24 N_20 S1 N_12 VDD mp5  l=0.42u w=0.6u m=1
M25 Y N_12 VDD VDD mp5  l=0.42u w=0.62u m=1
M26 N_13 S1 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends mx04d0
* SPICE INPUT		Mon Sep 24 12:29:14 2018	mx04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d1
.subckt mx04d1 S0 A B D C S1 GND VDD Y
M1 N_20 N_13 N_12 GND mn5  l=0.5u w=0.6u m=1
M2 N_23 S1 N_12 GND mn5  l=0.5u w=0.6u m=1
M3 Y N_12 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_13 S1 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_25 C GND GND mn5  l=0.5u w=0.6u m=1
M6 N_23 N_5 N_25 GND mn5  l=0.5u w=0.6u m=1
M7 GND D N_24 GND mn5  l=0.5u w=0.6u m=1
M8 N_22 B GND GND mn5  l=0.5u w=0.6u m=1
M9 N_20 S0 N_22 GND mn5  l=0.5u w=0.6u m=1
M10 N_20 N_5 N_21 GND mn5  l=0.5u w=0.6u m=1
M11 N_21 A GND GND mn5  l=0.5u w=0.6u m=1
M12 N_23 S0 N_24 GND mn5  l=0.5u w=0.6u m=1
M13 N_5 S0 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_25 C VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_24 N_5 N_23 VDD mp5  l=0.42u w=0.6u m=1
M16 N_24 D VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_23 S0 N_25 VDD mp5  l=0.42u w=0.6u m=1
M18 N_5 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_22 B VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_20 N_5 N_22 VDD mp5  l=0.42u w=0.6u m=1
M21 N_20 S0 N_21 VDD mp5  l=0.42u w=0.6u m=1
M22 N_21 A VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.6u m=1
M24 N_20 S1 N_12 VDD mp5  l=0.42u w=0.6u m=1
M25 Y N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 N_13 S1 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends mx04d1
* SPICE INPUT		Mon Sep 24 12:29:22 2018	mx04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d2
.subckt mx04d2 S0 A B D C S1 GND VDD Y
M1 N_20 N_13 N_12 GND mn5  l=0.5u w=0.6u m=1
M2 N_23 S1 N_12 GND mn5  l=0.5u w=0.6u m=1
M3 Y N_12 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_13 S1 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_25 C GND GND mn5  l=0.5u w=0.6u m=1
M6 N_23 N_5 N_25 GND mn5  l=0.5u w=0.6u m=1
M7 GND D N_24 GND mn5  l=0.5u w=0.6u m=1
M8 N_22 B GND GND mn5  l=0.5u w=0.6u m=1
M9 N_20 S0 N_22 GND mn5  l=0.5u w=0.6u m=1
M10 N_20 N_5 N_21 GND mn5  l=0.5u w=0.6u m=1
M11 N_21 A GND GND mn5  l=0.5u w=0.6u m=1
M12 N_23 S0 N_24 GND mn5  l=0.5u w=0.6u m=1
M13 N_5 S0 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_25 C VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_24 N_5 N_23 VDD mp5  l=0.42u w=0.6u m=1
M16 N_24 D VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_23 S0 N_25 VDD mp5  l=0.42u w=0.6u m=1
M18 N_5 S0 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_22 B VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_20 N_5 N_22 VDD mp5  l=0.42u w=0.6u m=1
M21 N_20 S0 N_21 VDD mp5  l=0.42u w=0.6u m=1
M22 N_21 A VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_23 N_13 N_12 VDD mp5  l=0.42u w=0.6u m=1
M24 N_20 S1 N_12 VDD mp5  l=0.42u w=0.6u m=1
M25 Y N_12 VDD VDD mp5  l=0.42u w=1.28u m=1
M26 N_13 S1 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends mx04d2
* SPICE INPUT		Mon Sep 24 12:29:30 2018	nd02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d0
.subckt nd02d0 Y GND VDD B A
M1 Y A N_5 GND mn5  l=0.5u w=0.6u m=1
M2 GND B N_5 GND mn5  l=0.5u w=0.6u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.62u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.62u m=1
.ends nd02d0
* SPICE INPUT		Mon Sep 24 12:29:38 2018	nd02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d1
.subckt nd02d1 Y GND VDD B A
M1 Y A N_5 GND mn5  l=0.5u w=0.72u m=1
M2 GND B N_5 GND mn5  l=0.5u w=0.72u m=1
M3 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd02d1
* SPICE INPUT		Mon Sep 24 12:29:46 2018	nd02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d2
.subckt nd02d2 Y GND VDD A B
M1 GND B N_5 GND mn5  l=0.5u w=0.98u m=1
M2 Y A N_5 GND mn5  l=0.5u w=0.98u m=1
M3 Y B VDD VDD mp5  l=0.42u w=1.28u m=1
M4 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
.ends nd02d2
* SPICE INPUT		Mon Sep 24 12:29:54 2018	nd03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d0
.subckt nd03d0 A C B GND Y VDD
M1 N_9 B N_8 GND mn5  l=0.5u w=0.6u m=1
M2 N_9 C GND GND mn5  l=0.5u w=0.6u m=1
M3 Y A N_8 GND mn5  l=0.5u w=0.6u m=1
M4 Y B VDD VDD mp5  l=0.42u w=0.62u m=1
M5 Y C VDD VDD mp5  l=0.42u w=0.62u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends nd03d0
* SPICE INPUT		Mon Sep 24 12:30:02 2018	nd03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d1
.subckt nd03d1 C B A GND Y VDD
M1 Y A N_8 GND mn5  l=0.5u w=0.72u m=1
M2 N_9 B N_8 GND mn5  l=0.5u w=0.72u m=1
M3 N_9 C GND GND mn5  l=0.5u w=0.72u m=1
M4 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M5 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd03d1
* SPICE INPUT		Mon Sep 24 12:30:10 2018	nd03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d2
.subckt nd03d2 C B A GND Y VDD
M1 Y A N_8 GND mn5  l=0.5u w=0.98u m=1
M2 N_9 B N_8 GND mn5  l=0.5u w=0.98u m=1
M3 N_9 C GND GND mn5  l=0.5u w=0.98u m=1
M4 Y A VDD VDD mp5  l=0.42u w=1.28u m=1
M5 Y B VDD VDD mp5  l=0.42u w=1.28u m=1
M6 Y C VDD VDD mp5  l=0.42u w=1.28u m=1
.ends nd03d2
* SPICE INPUT		Mon Sep 24 12:30:17 2018	nd04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d0
.subckt nd04d0 C B A D VDD Y GND
M1 N_10 D GND GND mn5  l=0.5u w=0.6u m=1
M2 Y A N_9 GND mn5  l=0.5u w=0.6u m=1
M3 N_11 B N_9 GND mn5  l=0.5u w=0.6u m=1
M4 N_11 C N_10 GND mn5  l=0.5u w=0.6u m=1
M5 Y D VDD VDD mp5  l=0.42u w=0.62u m=1
M6 Y A VDD VDD mp5  l=0.42u w=0.62u m=1
M7 VDD B Y VDD mp5  l=0.42u w=0.62u m=1
M8 VDD C Y VDD mp5  l=0.42u w=0.62u m=1
.ends nd04d0
* SPICE INPUT		Mon Sep 24 12:30:25 2018	nd04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d1
.subckt nd04d1 B C D A Y GND VDD
M1 Y A N_9 GND mn5  l=0.5u w=0.72u m=1
M2 N_10 D GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 C N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_11 B N_9 GND mn5  l=0.5u w=0.72u m=1
M5 Y A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y D VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M8 VDD B Y VDD mp5  l=0.42u w=0.96u m=1
.ends nd04d1
* SPICE INPUT		Mon Sep 24 12:30:33 2018	nd04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d2
.subckt nd04d2 A B C D GND Y VDD
M1 N_10 D GND GND mn5  l=0.5u w=0.98u m=1
M2 N_11 C N_10 GND mn5  l=0.5u w=0.98u m=1
M3 N_11 B N_9 GND mn5  l=0.5u w=0.98u m=1
M4 Y A N_9 GND mn5  l=0.5u w=0.98u m=1
M5 Y D VDD VDD mp5  l=0.42u w=1.28u m=1
M6 VDD C Y VDD mp5  l=0.42u w=1.28u m=1
M7 VDD B Y VDD mp5  l=0.42u w=1.28u m=1
M8 VDD A Y VDD mp5  l=0.42u w=1.28u m=1
.ends nd04d2
* SPICE INPUT		Mon Sep 24 12:30:41 2018	nd12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d0
.subckt nd12d0 AN B Y VDD GND
M1 GND B N_12 GND mn5  l=0.5u w=0.6u m=1
M2 Y N_3 N_12 GND mn5  l=0.5u w=0.6u m=1
M3 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M4 VDD B Y VDD mp5  l=0.42u w=0.62u m=1
M5 VDD N_3 Y VDD mp5  l=0.42u w=0.62u m=1
M6 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends nd12d0
* SPICE INPUT		Mon Sep 24 12:30:50 2018	nd12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d1
.subckt nd12d1 AN B VDD GND Y
M1 GND B N_8 GND mn5  l=0.5u w=0.72u m=1
M2 Y N_3 N_8 GND mn5  l=0.5u w=0.72u m=1
M3 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M4 VDD B Y VDD mp5  l=0.42u w=0.96u m=1
M5 VDD N_3 Y VDD mp5  l=0.42u w=0.96u m=1
M6 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends nd12d1
* SPICE INPUT		Mon Sep 24 12:30:58 2018	nd12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d2
.subckt nd12d2 AN B GND Y VDD
M1 GND B N_8 GND mn5  l=0.5u w=0.98u m=1
M2 Y N_3 N_8 GND mn5  l=0.5u w=0.98u m=1
M3 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M4 VDD B Y VDD mp5  l=0.42u w=1.28u m=1
M5 VDD N_3 Y VDD mp5  l=0.42u w=1.28u m=1
M6 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends nd12d2
* SPICE INPUT		Mon Sep 24 12:31:07 2018	nd13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d0
.subckt nd13d0 AN B C GND VDD Y
M1 N_14 C GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_4 N_13 GND mn5  l=0.5u w=0.6u m=1
M3 N_14 B N_13 GND mn5  l=0.5u w=0.6u m=1
M4 N_4 AN GND GND mn5  l=0.5u w=0.6u m=1
M5 Y C VDD VDD mp5  l=0.42u w=0.62u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 VDD AN N_4 VDD mp5  l=0.42u w=0.62u m=1
.ends nd13d0
* SPICE INPUT		Mon Sep 24 12:31:16 2018	nd13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d1
.subckt nd13d1 AN B C GND VDD Y
M1 N_10 C GND GND mn5  l=0.5u w=0.72u m=1
M2 Y N_4 N_9 GND mn5  l=0.5u w=0.72u m=1
M3 N_10 B N_9 GND mn5  l=0.5u w=0.72u m=1
M4 N_4 AN GND GND mn5  l=0.5u w=0.6u m=1
M5 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y B VDD VDD mp5  l=0.42u w=0.96u m=1
M8 VDD AN N_4 VDD mp5  l=0.42u w=0.62u m=1
.ends nd13d1
* SPICE INPUT		Mon Sep 24 12:31:25 2018	nd13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d2
.subckt nd13d2 B C AN VDD Y GND
M1 N_4 AN GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_4 N_9 GND mn5  l=0.5u w=0.98u m=1
M3 N_10 C GND GND mn5  l=0.5u w=0.98u m=1
M4 N_10 B N_9 GND mn5  l=0.5u w=0.98u m=1
M5 VDD AN N_4 VDD mp5  l=0.42u w=0.62u m=1
M6 Y N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 Y C VDD VDD mp5  l=0.42u w=1.28u m=1
M8 Y B VDD VDD mp5  l=0.42u w=1.28u m=1
.ends nd13d2
* SPICE INPUT		Mon Sep 24 12:31:33 2018	nd14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d0
.subckt nd14d0 D AN C B GND Y VDD
M1 Y N_6 N_10 GND mn5  l=0.5u w=0.6u m=1
M2 N_12 B N_10 GND mn5  l=0.5u w=0.6u m=1
M3 N_12 C N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_6 AN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_11 D GND GND mn5  l=0.5u w=0.6u m=1
M6 VDD N_6 Y VDD mp5  l=0.42u w=0.62u m=1
M7 VDD B Y VDD mp5  l=0.42u w=0.62u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.62u m=1
M9 VDD AN N_6 VDD mp5  l=0.42u w=0.62u m=1
M10 Y D VDD VDD mp5  l=0.42u w=0.62u m=1
.ends nd14d0
* SPICE INPUT		Mon Sep 24 12:31:41 2018	nd14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d1
.subckt nd14d1 D AN C B GND Y VDD
M1 Y N_6 N_10 GND mn5  l=0.5u w=0.72u m=1
M2 N_12 B N_10 GND mn5  l=0.5u w=0.72u m=1
M3 N_12 C N_11 GND mn5  l=0.5u w=0.72u m=1
M4 N_6 AN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_11 D GND GND mn5  l=0.5u w=0.72u m=1
M6 VDD N_6 Y VDD mp5  l=0.42u w=0.96u m=1
M7 VDD B Y VDD mp5  l=0.42u w=0.96u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M9 VDD AN N_6 VDD mp5  l=0.42u w=0.62u m=1
M10 Y D VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd14d1
* SPICE INPUT		Mon Sep 24 12:31:50 2018	nd14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d2
.subckt nd14d2 Y GND VDD C D B AN
M1 Y N_4 N_6 GND mn5  l=0.5u w=0.98u m=1
M2 N_8 B N_6 GND mn5  l=0.5u w=0.98u m=1
M3 N_8 C N_7 GND mn5  l=0.5u w=0.98u m=1
M4 N_4 AN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_7 D GND GND mn5  l=0.5u w=0.98u m=1
M6 VDD N_4 Y VDD mp5  l=0.42u w=1.28u m=1
M7 VDD B Y VDD mp5  l=0.42u w=1.28u m=1
M8 VDD C Y VDD mp5  l=0.42u w=1.28u m=1
M9 VDD AN N_4 VDD mp5  l=0.42u w=0.62u m=1
M10 Y D VDD VDD mp5  l=0.42u w=1.28u m=1
.ends nd14d2
* SPICE INPUT		Mon Sep 24 12:31:58 2018	nd23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd23d0
.subckt nd23d0 C BN AN Y GND VDD
M1 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_2 BN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_16 C GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 N_15 GND mn5  l=0.5u w=0.6u m=1
M5 N_16 N_2 N_15 GND mn5  l=0.5u w=0.6u m=1
M6 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_2 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends nd23d0
* SPICE INPUT		Mon Sep 24 12:32:07 2018	nd23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd23d1
.subckt nd23d1 C BN AN GND VDD Y
M1 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 BN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_11 C GND GND mn5  l=0.5u w=0.72u m=1
M4 N_11 N_3 N_10 GND mn5  l=0.5u w=0.72u m=1
M5 Y N_2 N_10 GND mn5  l=0.5u w=0.72u m=1
M6 N_2 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends nd23d1
* SPICE INPUT		Mon Sep 24 12:32:15 2018	nd23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd23d2
.subckt nd23d2 C BN AN GND VDD Y
M1 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 BN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_11 C GND GND mn5  l=0.5u w=0.98u m=1
M4 N_11 N_3 N_10 GND mn5  l=0.5u w=0.98u m=1
M5 Y N_2 N_10 GND mn5  l=0.5u w=0.98u m=1
M6 N_2 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y C VDD VDD mp5  l=0.42u w=1.28u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M10 Y N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends nd23d2
* SPICE INPUT		Mon Sep 24 12:32:24 2018	nd24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d0
.subckt nd24d0 BN C D AN GND Y VDD
M1 Y N_7 N_11 GND mn5  l=0.5u w=0.6u m=1
M2 N_7 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 D GND GND mn5  l=0.5u w=0.6u m=1
M4 N_13 C N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_13 N_3 N_11 GND mn5  l=0.5u w=0.6u m=1
M6 N_3 BN GND GND mn5  l=0.5u w=0.6u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_7 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y D VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y C VDD VDD mp5  l=0.42u w=0.62u m=1
M11 VDD N_3 Y VDD mp5  l=0.42u w=0.62u m=1
M12 N_3 BN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends nd24d0
* SPICE INPUT		Mon Sep 24 12:32:33 2018	nd24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d1
.subckt nd24d1 BN C D AN GND Y VDD
M1 Y N_7 N_11 GND mn5  l=0.5u w=0.72u m=1
M2 N_7 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 D GND GND mn5  l=0.5u w=0.72u m=1
M4 N_13 C N_12 GND mn5  l=0.5u w=0.72u m=1
M5 N_13 N_3 N_11 GND mn5  l=0.5u w=0.72u m=1
M6 N_3 BN GND GND mn5  l=0.5u w=0.6u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_7 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y D VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y C VDD VDD mp5  l=0.42u w=0.96u m=1
M11 VDD N_3 Y VDD mp5  l=0.42u w=0.96u m=1
M12 N_3 BN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends nd24d1
* SPICE INPUT		Mon Sep 24 12:32:42 2018	nd24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d2
.subckt nd24d2 D C AN BN GND VDD Y
M1 N_5 BN GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_6 N_11 GND mn5  l=0.5u w=0.98u m=1
M3 N_13 N_5 N_11 GND mn5  l=0.5u w=0.98u m=1
M4 N_6 AN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_13 C N_12 GND mn5  l=0.5u w=0.98u m=1
M6 N_12 D GND GND mn5  l=0.5u w=0.98u m=1
M7 N_5 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M9 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M10 N_6 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M11 VDD C Y VDD mp5  l=0.42u w=1.28u m=1
M12 Y D VDD VDD mp5  l=0.42u w=1.28u m=1
.ends nd24d2
* SPICE INPUT		Mon Sep 24 12:32:50 2018	nr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d0
.subckt nr02d0 GND VDD Y B A
M1 GND B Y GND mn5  l=0.5u w=0.6u m=1
M2 GND A Y GND mn5  l=0.5u w=0.6u m=1
M3 Y B N_7 VDD mp5  l=0.42u w=0.62u m=1
M4 VDD A N_7 VDD mp5  l=0.42u w=0.62u m=1
.ends nr02d0
* SPICE INPUT		Mon Sep 24 12:32:58 2018	nr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d1
.subckt nr02d1 Y VDD GND A B
M1 GND B Y GND mn5  l=0.5u w=0.72u m=1
M2 GND A Y GND mn5  l=0.5u w=0.72u m=1
M3 Y B N_5 VDD mp5  l=0.42u w=0.96u m=1
M4 VDD A N_5 VDD mp5  l=0.42u w=0.96u m=1
.ends nr02d1
* SPICE INPUT		Mon Sep 24 12:33:06 2018	nr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d2
.subckt nr02d2 Y VDD GND A B
M1 GND B Y GND mn5  l=0.5u w=0.98u m=1
M2 GND A Y GND mn5  l=0.5u w=0.98u m=1
M3 Y B N_5 VDD mp5  l=0.42u w=1.28u m=1
M4 VDD A N_5 VDD mp5  l=0.42u w=1.28u m=1
.ends nr02d2
* SPICE INPUT		Mon Sep 24 12:33:15 2018	nr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d0
.subckt nr03d0 B A C Y VDD GND
M1 Y C GND GND mn5  l=0.5u w=0.6u m=1
M2 Y A GND GND mn5  l=0.5u w=0.6u m=1
M3 Y B GND GND mn5  l=0.5u w=0.6u m=1
M4 Y C N_8 VDD mp5  l=0.42u w=0.62u m=1
M5 N_9 A VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_9 B N_8 VDD mp5  l=0.42u w=0.62u m=1
.ends nr03d0
* SPICE INPUT		Mon Sep 24 12:33:23 2018	nr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d1
.subckt nr03d1 B A C Y VDD GND
M1 Y C GND GND mn5  l=0.5u w=0.72u m=1
M2 Y A GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C N_8 VDD mp5  l=0.42u w=0.96u m=1
M5 N_9 A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_9 B N_8 VDD mp5  l=0.42u w=0.96u m=1
.ends nr03d1
* SPICE INPUT		Mon Sep 24 12:33:32 2018	nr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d2
.subckt nr03d2 B C A VDD Y GND
M1 Y A GND GND mn5  l=0.5u w=0.98u m=1
M2 Y C GND GND mn5  l=0.5u w=0.98u m=1
M3 Y B GND GND mn5  l=0.5u w=0.98u m=1
M4 N_9 A VDD VDD mp5  l=0.42u w=1.28u m=1
M5 Y C N_8 VDD mp5  l=0.42u w=1.28u m=1
M6 N_9 B N_8 VDD mp5  l=0.42u w=1.28u m=1
.ends nr03d2
* SPICE INPUT		Mon Sep 24 12:33:40 2018	nr04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d0
.subckt nr04d0 C D B A VDD Y GND
M1 Y A GND GND mn5  l=0.5u w=0.6u m=1
M2 Y B GND GND mn5  l=0.5u w=0.6u m=1
M3 Y D GND GND mn5  l=0.5u w=0.6u m=1
M4 GND C Y GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_11 B N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 Y D N_9 VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 C N_9 VDD mp5  l=0.42u w=0.62u m=1
.ends nr04d0
* SPICE INPUT		Mon Sep 24 12:33:49 2018	nr04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d1
.subckt nr04d1 C D B A VDD Y GND
M1 Y A GND GND mn5  l=0.5u w=0.72u m=1
M2 Y B GND GND mn5  l=0.5u w=0.72u m=1
M3 Y D GND GND mn5  l=0.5u w=0.72u m=1
M4 GND C Y GND mn5  l=0.5u w=0.72u m=1
M5 N_10 A VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_11 B N_10 VDD mp5  l=0.42u w=0.96u m=1
M7 Y D N_9 VDD mp5  l=0.42u w=0.96u m=1
M8 N_11 C N_9 VDD mp5  l=0.42u w=0.96u m=1
.ends nr04d1
* SPICE INPUT		Mon Sep 24 12:33:58 2018	nr04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d2
.subckt nr04d2 D B A C Y VDD GND
M1 GND C Y GND mn5  l=0.5u w=0.98u m=1
M2 Y A GND GND mn5  l=0.5u w=0.98u m=1
M3 GND B Y GND mn5  l=0.5u w=0.98u m=1
M4 GND D Y GND mn5  l=0.5u w=0.98u m=1
M5 N_11 C N_9 VDD mp5  l=0.42u w=1.28u m=1
M6 N_10 A VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_11 B N_10 VDD mp5  l=0.42u w=1.28u m=1
M8 Y D N_9 VDD mp5  l=0.42u w=1.28u m=1
.ends nr04d2
* SPICE INPUT		Mon Sep 24 12:34:12 2018	nr12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d0
.subckt nr12d0 AN B VDD Y GND
M1 Y B GND GND mn5  l=0.5u w=0.6u m=1
M2 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 GND N_2 Y GND mn5  l=0.5u w=0.6u m=1
M4 Y B N_8 VDD mp5  l=0.42u w=0.62u m=1
M5 VDD AN N_2 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD N_2 N_8 VDD mp5  l=0.42u w=0.62u m=1
.ends nr12d0
* SPICE INPUT		Mon Sep 24 12:34:21 2018	nr12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d1
.subckt nr12d1 AN B VDD Y GND
M1 Y B GND GND mn5  l=0.5u w=0.72u m=1
M2 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 GND N_2 Y GND mn5  l=0.5u w=0.72u m=1
M4 Y B N_8 VDD mp5  l=0.42u w=0.96u m=1
M5 VDD AN N_2 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD N_2 N_8 VDD mp5  l=0.42u w=0.96u m=1
.ends nr12d1
* SPICE INPUT		Mon Sep 24 12:34:30 2018	nr12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d2
.subckt nr12d2 AN B VDD Y GND
M1 GND B Y GND mn5  l=0.5u w=0.98u m=1
M2 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 GND N_2 Y GND mn5  l=0.5u w=0.98u m=1
M4 Y B N_8 VDD mp5  l=0.42u w=1.28u m=1
M5 VDD AN N_2 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD N_2 N_8 VDD mp5  l=0.42u w=1.28u m=1
.ends nr12d2
* SPICE INPUT		Mon Sep 24 12:34:38 2018	nr13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d0
.subckt nr13d0 C AN B VDD Y GND
M1 Y B GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.6u m=1
M4 Y C GND GND mn5  l=0.5u w=0.6u m=1
M5 N_10 B N_9 VDD mp5  l=0.42u w=0.62u m=1
M6 VDD AN N_3 VDD mp5  l=0.42u w=0.62u m=1
M7 N_10 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y C N_9 VDD mp5  l=0.42u w=0.62u m=1
.ends nr13d0
* SPICE INPUT		Mon Sep 24 12:34:46 2018	nr13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d1
.subckt nr13d1 C AN B VDD Y GND
M1 Y B GND GND mn5  l=0.5u w=0.72u m=1
M2 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y C GND GND mn5  l=0.5u w=0.72u m=1
M5 N_10 B N_9 VDD mp5  l=0.42u w=0.96u m=1
M6 VDD AN N_3 VDD mp5  l=0.42u w=0.62u m=1
M7 N_10 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y C N_9 VDD mp5  l=0.42u w=0.96u m=1
.ends nr13d1
* SPICE INPUT		Mon Sep 24 12:34:55 2018	nr13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d2
.subckt nr13d2 B AN C Y GND VDD
M1 Y C GND GND mn5  l=0.5u w=0.98u m=1
M2 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 Y B GND GND mn5  l=0.5u w=0.98u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.98u m=1
M5 Y C N_9 VDD mp5  l=0.42u w=1.28u m=1
M6 VDD AN N_2 VDD mp5  l=0.42u w=0.62u m=1
M7 N_10 B N_9 VDD mp5  l=0.42u w=1.28u m=1
M8 N_10 N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends nr13d2
* SPICE INPUT		Mon Sep 24 12:35:04 2018	nr14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d0
.subckt nr14d0 D C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.6u m=1
M3 Y B GND GND mn5  l=0.5u w=0.6u m=1
M4 GND C Y GND mn5  l=0.5u w=0.6u m=1
M5 Y D GND GND mn5  l=0.5u w=0.6u m=1
M6 VDD AN N_5 VDD mp5  l=0.42u w=0.62u m=1
M7 N_11 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_12 B N_11 VDD mp5  l=0.42u w=0.62u m=1
M9 N_12 C N_10 VDD mp5  l=0.42u w=0.62u m=1
M10 Y D N_10 VDD mp5  l=0.42u w=0.62u m=1
.ends nr14d0
* SPICE INPUT		Mon Sep 24 12:35:13 2018	nr14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d1
.subckt nr14d1 D C B AN GND VDD Y
M1 N_5 AN GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B GND GND mn5  l=0.5u w=0.72u m=1
M4 GND C Y GND mn5  l=0.5u w=0.72u m=1
M5 Y D GND GND mn5  l=0.5u w=0.72u m=1
M6 VDD AN N_5 VDD mp5  l=0.42u w=0.62u m=1
M7 N_11 N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_12 B N_11 VDD mp5  l=0.42u w=0.96u m=1
M9 N_12 C N_10 VDD mp5  l=0.42u w=0.96u m=1
M10 Y D N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends nr14d1
* SPICE INPUT		Mon Sep 24 12:35:21 2018	nr14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d2
.subckt nr14d2 Y VDD GND D C B AN
M1 GND C Y GND mn5  l=0.5u w=0.98u m=1
M2 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 GND B Y GND mn5  l=0.5u w=0.98u m=1
M4 GND D Y GND mn5  l=0.5u w=0.98u m=1
M5 Y N_3 GND GND mn5  l=0.5u w=0.98u m=1
M6 N_8 C N_6 VDD mp5  l=0.42u w=1.28u m=1
M7 VDD AN N_3 VDD mp5  l=0.42u w=0.62u m=1
M8 N_8 B N_7 VDD mp5  l=0.42u w=1.28u m=1
M9 Y D N_6 VDD mp5  l=0.42u w=1.28u m=1
M10 N_7 N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends nr14d2
* SPICE INPUT		Mon Sep 24 12:35:30 2018	nr23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr23d0
.subckt nr23d0 AN BN C VDD GND Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.6u m=1
M3 Y C GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 BN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_6 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_5 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_6 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_11 N_5 N_10 VDD mp5  l=0.42u w=0.62u m=1
M10 Y C N_10 VDD mp5  l=0.42u w=0.62u m=1
.ends nr23d0
* SPICE INPUT		Mon Sep 24 12:35:39 2018	nr23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr23d1
.subckt nr23d1 AN BN C VDD GND Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y C GND GND mn5  l=0.5u w=0.72u m=1
M4 N_5 BN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_6 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_5 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_6 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_11 N_5 N_10 VDD mp5  l=0.42u w=0.96u m=1
M10 Y C N_10 VDD mp5  l=0.42u w=0.96u m=1
.ends nr23d1
* SPICE INPUT		Mon Sep 24 12:35:47 2018	nr23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr23d2
.subckt nr23d2 AN BN C VDD Y GND
M1 Y C GND GND mn5  l=0.5u w=0.98u m=1
M2 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M3 Y N_4 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_5 BN GND GND mn5  l=0.5u w=0.6u m=1
M5 N_4 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_5 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_4 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y C N_10 VDD mp5  l=0.42u w=1.28u m=1
M9 N_11 N_5 N_10 VDD mp5  l=0.42u w=1.28u m=1
M10 N_11 N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends nr23d2
* SPICE INPUT		Mon Sep 24 12:36:00 2018	nr24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d0
.subckt nr24d0 AN BN D C VDD Y GND
M1 Y N_7 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_6 GND GND mn5  l=0.5u w=0.6u m=1
M3 GND C Y GND mn5  l=0.5u w=0.6u m=1
M4 Y D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_6 BN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 AN GND GND mn5  l=0.5u w=0.6u m=1
M7 N_6 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_7 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_12 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.62u m=1
M11 N_13 C N_11 VDD mp5  l=0.42u w=0.62u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=0.62u m=1
.ends nr24d0
* SPICE INPUT		Mon Sep 24 12:36:09 2018	nr24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d1
.subckt nr24d1 AN BN D C VDD Y GND
M1 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M3 GND C Y GND mn5  l=0.5u w=0.72u m=1
M4 Y D GND GND mn5  l=0.5u w=0.72u m=1
M5 N_6 BN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 AN GND GND mn5  l=0.5u w=0.6u m=1
M7 N_6 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_7 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_12 N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_13 N_6 N_12 VDD mp5  l=0.42u w=0.96u m=1
M11 N_13 C N_11 VDD mp5  l=0.42u w=0.96u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=0.96u m=1
.ends nr24d1
* SPICE INPUT		Mon Sep 24 12:36:17 2018	nr24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d2
.subckt nr24d2 BN AN D C GND VDD Y
M1 GND C Y GND mn5  l=0.5u w=0.98u m=1
M2 GND N_6 Y GND mn5  l=0.5u w=0.98u m=1
M3 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M4 GND D Y GND mn5  l=0.5u w=0.98u m=1
M5 N_5 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_6 BN GND GND mn5  l=0.5u w=0.6u m=1
M7 N_5 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 BN VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_13 C N_11 VDD mp5  l=0.42u w=1.28u m=1
M10 N_13 N_6 N_12 VDD mp5  l=0.42u w=1.28u m=1
M11 N_12 N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 Y D N_11 VDD mp5  l=0.42u w=1.28u m=1
.ends nr24d2
* SPICE INPUT		Mon Sep 24 12:36:26 2018	oai211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d0
.subckt oai211d0 C0 B0 A1 A0 VDD GND Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_9 B0 N_16 GND mn5  l=0.5u w=0.6u m=1
M4 Y C0 N_16 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M6 Y A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends oai211d0
* SPICE INPUT		Mon Sep 24 12:36:34 2018	oai211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d1
.subckt oai211d1 C0 B0 A1 A0 GND VDD Y
M1 N_9 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 B0 N_16 GND mn5  l=0.5u w=0.72u m=1
M4 Y C0 N_16 GND mn5  l=0.5u w=0.72u m=1
M5 N_10 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 Y A1 N_10 VDD mp5  l=0.42u w=0.96u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oai211d1
* SPICE INPUT		Mon Sep 24 12:36:43 2018	oai211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d2
.subckt oai211d2 VDD Y GND C0 B0 A1 A0
M1 GND A0 N_10 GND mn5  l=0.5u w=0.98u m=1
M2 N_10 A1 GND GND mn5  l=0.5u w=0.98u m=1
M3 Y C0 N_18 GND mn5  l=0.5u w=0.98u m=1
M4 N_10 B0 N_18 GND mn5  l=0.5u w=0.98u m=1
M5 N_7 A0 VDD VDD mp5  l=0.42u w=1.28u m=1
M6 Y A1 N_7 VDD mp5  l=0.42u w=1.28u m=1
M7 Y C0 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 Y B0 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends oai211d2
* SPICE INPUT		Mon Sep 24 12:36:51 2018	oai21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d0
.subckt oai21d0 B0 A1 A0 Y VDD GND
M1 N_8 A0 GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A1 N_8 GND mn5  l=0.5u w=0.6u m=1
M3 N_8 B0 Y GND mn5  l=0.5u w=0.6u m=1
M4 N_9 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M5 N_9 A1 Y VDD mp5  l=0.42u w=0.62u m=1
M6 VDD B0 Y VDD mp5  l=0.42u w=0.62u m=1
.ends oai21d0
* SPICE INPUT		Mon Sep 24 12:36:58 2018	oai21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d1
.subckt oai21d1 B0 A1 A0 Y VDD GND
M1 N_8 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 GND A1 N_8 GND mn5  l=0.5u w=0.72u m=1
M3 N_8 B0 Y GND mn5  l=0.5u w=0.72u m=1
M4 N_9 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M5 N_9 A1 Y VDD mp5  l=0.42u w=0.96u m=1
M6 VDD B0 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai21d1
* SPICE INPUT		Mon Sep 24 12:37:06 2018	oai21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d2
.subckt oai21d2 A0 A1 B0 Y VDD GND
M1 N_5 B0 Y GND mn5  l=0.5u w=0.98u m=1
M2 GND A1 N_5 GND mn5  l=0.5u w=0.98u m=1
M3 GND A0 N_5 GND mn5  l=0.5u w=0.98u m=1
M4 VDD B0 Y VDD mp5  l=0.42u w=1.28u m=1
M5 N_9 A1 Y VDD mp5  l=0.42u w=1.28u m=1
M6 N_9 A0 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends oai21d2
* SPICE INPUT		Mon Sep 24 12:37:14 2018	oai221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d0
.subckt oai221d0 B0 B1 A1 A0 C0 Y VDD GND
M1 Y C0 N_8 GND mn5  l=0.5u w=0.6u m=1
M2 N_9 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_9 A1 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_9 B1 N_8 GND mn5  l=0.5u w=0.6u m=1
M5 N_8 B0 N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_12 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y A1 N_12 VDD mp5  l=0.42u w=0.62u m=1
M8 N_13 B1 Y VDD mp5  l=0.42u w=0.62u m=1
M9 N_13 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends oai221d0
* SPICE INPUT		Mon Sep 24 12:37:22 2018	oai221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d1
.subckt oai221d1 C0 B0 B1 A1 A0 GND VDD Y
M1 GND A0 N_11 GND mn5  l=0.5u w=0.72u m=1
M2 N_11 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_11 B1 N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_11 B0 N_10 GND mn5  l=0.5u w=0.72u m=1
M5 Y C0 N_10 GND mn5  l=0.5u w=0.72u m=1
M6 N_12 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y A1 N_12 VDD mp5  l=0.42u w=0.96u m=1
M8 N_13 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M9 N_13 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oai221d1
* SPICE INPUT		Mon Sep 24 12:37:30 2018	oai221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d2
.subckt oai221d2 C0 A0 A1 B1 B0 GND VDD Y
M1 N_11 B0 N_10 GND mn5  l=0.5u w=0.98u m=1
M2 N_11 B1 N_10 GND mn5  l=0.5u w=0.98u m=1
M3 N_11 A1 GND GND mn5  l=0.5u w=0.98u m=1
M4 GND A0 N_11 GND mn5  l=0.5u w=0.98u m=1
M5 Y C0 N_10 GND mn5  l=0.5u w=0.98u m=1
M6 Y C0 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_13 B0 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 N_13 B1 Y VDD mp5  l=0.42u w=1.28u m=1
M9 Y A1 N_12 VDD mp5  l=0.42u w=1.28u m=1
M10 N_12 A0 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends oai221d2
* SPICE INPUT		Mon Sep 24 12:37:38 2018	oai222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d0
.subckt oai222d0 C0 B1 A0 B0 A1 C1 GND Y VDD
M1 N_9 C1 Y GND mn5  l=0.5u w=0.6u m=1
M2 N_13 A1 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_13 B0 N_9 GND mn5  l=0.5u w=0.6u m=1
M4 N_13 A0 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_9 B1 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 N_9 C0 Y GND mn5  l=0.5u w=0.6u m=1
M7 Y A1 N_14 VDD mp5  l=0.42u w=0.62u m=1
M8 N_12 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 VDD A0 N_14 VDD mp5  l=0.42u w=0.62u m=1
M10 VDD C1 N_15 VDD mp5  l=0.42u w=0.62u m=1
M11 Y B1 N_12 VDD mp5  l=0.42u w=0.62u m=1
M12 Y C0 N_15 VDD mp5  l=0.42u w=0.62u m=1
.ends oai222d0
* SPICE INPUT		Mon Sep 24 12:37:46 2018	oai222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d1
.subckt oai222d1 C0 B1 A1 A0 B0 C1 VDD GND Y
M1 N_11 C1 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_13 B0 N_11 GND mn5  l=0.5u w=0.72u m=1
M3 N_13 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_13 A1 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_11 B1 N_13 GND mn5  l=0.5u w=0.72u m=1
M6 N_11 C0 Y GND mn5  l=0.5u w=0.72u m=1
M7 VDD B0 N_12 VDD mp5  l=0.42u w=0.96u m=1
M8 VDD A0 N_14 VDD mp5  l=0.42u w=0.96u m=1
M9 Y A1 N_14 VDD mp5  l=0.42u w=0.96u m=1
M10 VDD C1 N_15 VDD mp5  l=0.42u w=0.96u m=1
M11 Y B1 N_12 VDD mp5  l=0.42u w=0.96u m=1
M12 Y C0 N_15 VDD mp5  l=0.42u w=0.96u m=1
.ends oai222d1
* SPICE INPUT		Mon Sep 24 12:37:54 2018	oai222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d2
.subckt oai222d2 Y VDD GND C1 C0 B1 A1 A0 B0
M1 N_15 B0 N_11 GND mn5  l=0.5u w=0.98u m=1
M2 N_15 A0 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_15 A1 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_11 B1 N_15 GND mn5  l=0.5u w=0.98u m=1
M5 N_11 C0 Y GND mn5  l=0.5u w=0.98u m=1
M6 N_11 C1 Y GND mn5  l=0.5u w=0.98u m=1
M7 VDD B0 N_3 VDD mp5  l=0.42u w=1.28u m=1
M8 VDD A0 N_9 VDD mp5  l=0.42u w=1.28u m=1
M9 Y A1 N_9 VDD mp5  l=0.42u w=1.28u m=1
M10 Y B1 N_3 VDD mp5  l=0.42u w=1.28u m=1
M11 Y C0 N_10 VDD mp5  l=0.42u w=1.28u m=1
M12 VDD C1 N_10 VDD mp5  l=0.42u w=1.28u m=1
.ends oai222d2
* SPICE INPUT		Mon Sep 24 12:38:02 2018	oai22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d0
.subckt oai22d0 A0 A1 B0 B1 VDD GND Y
M1 Y B1 N_9 GND mn5  l=0.5u w=0.6u m=1
M2 Y B0 N_9 GND mn5  l=0.5u w=0.6u m=1
M3 N_9 A1 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_9 A0 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_11 B1 Y VDD mp5  l=0.42u w=0.62u m=1
M6 N_11 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 VDD A0 N_10 VDD mp5  l=0.42u w=0.62u m=1
.ends oai22d0
* SPICE INPUT		Mon Sep 24 12:38:10 2018	oai22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d1
.subckt oai22d1 B0 A0 A1 B1 VDD GND Y
M1 Y B1 N_9 GND mn5  l=0.5u w=0.72u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_9 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 N_9 GND mn5  l=0.5u w=0.72u m=1
M5 N_11 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M6 Y A1 N_10 VDD mp5  l=0.42u w=0.96u m=1
M7 VDD A0 N_10 VDD mp5  l=0.42u w=0.96u m=1
M8 N_11 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oai22d1
* SPICE INPUT		Mon Sep 24 12:38:19 2018	oai22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d2
.subckt oai22d2 A0 B1 B0 A1 Y GND VDD
M1 N_8 A1 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_8 B0 Y GND mn5  l=0.5u w=0.98u m=1
M3 Y B1 N_8 GND mn5  l=0.5u w=0.98u m=1
M4 N_8 A0 GND GND mn5  l=0.5u w=0.98u m=1
M5 Y A1 N_10 VDD mp5  l=0.42u w=1.28u m=1
M6 N_11 B0 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_11 B1 Y VDD mp5  l=0.42u w=1.28u m=1
M8 VDD A0 N_10 VDD mp5  l=0.42u w=1.28u m=1
.ends oai22d2
* SPICE INPUT		Mon Sep 24 12:38:27 2018	oai311d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai311d0
.subckt oai311d0 B0 C0 A0 A1 A2 Y VDD GND
M1 N_9 A2 GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A1 N_9 GND mn5  l=0.5u w=0.6u m=1
M3 N_9 A0 GND GND mn5  l=0.5u w=0.6u m=1
M4 Y C0 N_13 GND mn5  l=0.5u w=0.6u m=1
M5 N_9 B0 N_13 GND mn5  l=0.5u w=0.6u m=1
M6 N_11 A2 Y VDD mp5  l=0.42u w=0.62u m=1
M7 N_12 A1 N_11 VDD mp5  l=0.42u w=0.62u m=1
M8 N_12 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 VDD C0 Y VDD mp5  l=0.42u w=0.62u m=1
M10 VDD B0 Y VDD mp5  l=0.42u w=0.62u m=1
.ends oai311d0
* SPICE INPUT		Mon Sep 24 12:38:36 2018	oai311d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai311d1
.subckt oai311d1 B0 A1 A2 C0 A0 Y GND VDD
M1 N_8 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 Y C0 N_11 GND mn5  l=0.5u w=0.72u m=1
M3 N_8 A2 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_8 A1 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_8 B0 N_11 GND mn5  l=0.5u w=0.72u m=1
M6 N_18 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 VDD C0 Y VDD mp5  l=0.42u w=0.96u m=1
M8 N_17 A2 Y VDD mp5  l=0.42u w=0.96u m=1
M9 N_18 A1 N_17 VDD mp5  l=0.42u w=0.96u m=1
M10 VDD B0 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai311d1
* SPICE INPUT		Mon Sep 24 12:38:45 2018	oai311d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai311d2
.subckt oai311d2 B0 A1 A2 C0 A0 Y GND VDD
M1 N_7 A0 GND GND mn5  l=0.5u w=0.98u m=1
M2 Y C0 N_19 GND mn5  l=0.5u w=0.98u m=1
M3 N_7 A2 GND GND mn5  l=0.5u w=0.98u m=1
M4 GND A1 N_7 GND mn5  l=0.5u w=0.98u m=1
M5 N_7 B0 N_19 GND mn5  l=0.5u w=0.98u m=1
M6 VDD A0 N_12 VDD mp5  l=0.42u w=1.28u m=1
M7 VDD C0 Y VDD mp5  l=0.42u w=1.28u m=1
M8 N_11 A2 Y VDD mp5  l=0.42u w=1.28u m=1
M9 N_12 A1 N_11 VDD mp5  l=0.42u w=1.28u m=1
M10 VDD B0 Y VDD mp5  l=0.42u w=1.28u m=1
.ends oai311d2
* SPICE INPUT		Mon Sep 24 12:38:53 2018	oai31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d0
.subckt oai31d0 A2 B0 A1 A0 GND VDD Y
M1 GND A0 N_9 GND mn5  l=0.5u w=0.6u m=1
M2 GND A1 N_9 GND mn5  l=0.5u w=0.6u m=1
M3 Y B0 N_9 GND mn5  l=0.5u w=0.6u m=1
M4 N_9 A2 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_11 A0 N_10 VDD mp5  l=0.42u w=0.62u m=1
M6 N_11 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_10 A2 Y VDD mp5  l=0.42u w=0.62u m=1
.ends oai31d0
* SPICE INPUT		Mon Sep 24 12:39:02 2018	oai31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d1
.subckt oai31d1 A2 B0 A1 A0 Y GND VDD
M1 N_9 A0 GND GND mn5  l=0.5u w=0.72u m=1
M2 GND A1 N_9 GND mn5  l=0.5u w=0.72u m=1
M3 Y B0 N_9 GND mn5  l=0.5u w=0.72u m=1
M4 N_9 A2 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_11 A0 N_10 VDD mp5  l=0.42u w=0.96u m=1
M6 N_11 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=0.6u m=1
M8 N_10 A2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai31d1
* SPICE INPUT		Mon Sep 24 12:39:11 2018	oai31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d2
.subckt oai31d2 A2 A0 A1 B0 Y VDD GND
M1 Y B0 N_8 GND mn5  l=0.5u w=0.98u m=1
M2 GND A1 N_8 GND mn5  l=0.5u w=0.98u m=1
M3 GND A0 N_8 GND mn5  l=0.5u w=0.98u m=1
M4 N_8 A2 GND GND mn5  l=0.5u w=0.98u m=1
M5 Y B0 VDD VDD mp5  l=0.42u w=1.28u m=1
M6 N_11 A1 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_11 A0 N_10 VDD mp5  l=0.42u w=1.28u m=1
M8 N_10 A2 Y VDD mp5  l=0.42u w=1.28u m=1
.ends oai31d2
* SPICE INPUT		Mon Sep 24 12:39:21 2018	oai321d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai321d0
.subckt oai321d0 B1 B0 A0 A1 A2 C0 GND VDD Y
M1 Y C0 N_11 GND mn5  l=0.5u w=0.6u m=1
M2 N_12 A2 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 A1 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_12 A0 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_12 B0 N_11 GND mn5  l=0.5u w=0.6u m=1
M6 N_11 B1 N_12 GND mn5  l=0.5u w=0.6u m=1
M7 N_13 A2 Y VDD mp5  l=0.42u w=0.62u m=1
M8 N_14 A1 N_13 VDD mp5  l=0.42u w=0.62u m=1
M9 N_14 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_15 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_15 B1 Y VDD mp5  l=0.42u w=0.62u m=1
M12 Y C0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends oai321d0
* SPICE INPUT		Mon Sep 24 12:39:30 2018	oai321d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai321d1
.subckt oai321d1 C0 A1 A2 A0 B0 B1 GND VDD Y
M1 N_11 B1 N_12 GND mn5  l=0.5u w=0.72u m=1
M2 N_11 B0 N_12 GND mn5  l=0.5u w=0.72u m=1
M3 N_11 A0 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_11 A2 GND GND mn5  l=0.5u w=0.72u m=1
M5 GND A1 N_11 GND mn5  l=0.5u w=0.72u m=1
M6 Y C0 N_12 GND mn5  l=0.5u w=0.72u m=1
M7 VDD C0 Y VDD mp5  l=0.42u w=0.96u m=1
M8 N_15 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M9 N_15 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 VDD A0 N_14 VDD mp5  l=0.42u w=0.96u m=1
M11 N_13 A2 Y VDD mp5  l=0.42u w=0.96u m=1
M12 N_14 A1 N_13 VDD mp5  l=0.42u w=0.96u m=1
.ends oai321d1
* SPICE INPUT		Mon Sep 24 12:39:39 2018	oai321d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai321d2
.subckt oai321d2 Y VDD GND A0 B1 A1 C0 B0 A2
M1 N_13 B1 N_14 GND mn5  l=0.5u w=0.98u m=1
M2 N_13 B0 N_14 GND mn5  l=0.5u w=0.98u m=1
M3 N_13 A0 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_13 A2 GND GND mn5  l=0.5u w=0.98u m=1
M5 GND A1 N_13 GND mn5  l=0.5u w=0.98u m=1
M6 Y C0 N_14 GND mn5  l=0.5u w=0.98u m=1
M7 VDD C0 Y VDD mp5  l=0.42u w=1.28u m=1
M8 N_9 B1 Y VDD mp5  l=0.42u w=1.28u m=1
M9 N_9 B0 VDD VDD mp5  l=0.42u w=1.28u m=1
M10 VDD A0 N_8 VDD mp5  l=0.42u w=1.28u m=1
M11 N_7 A2 Y VDD mp5  l=0.42u w=1.28u m=1
M12 N_8 A1 N_7 VDD mp5  l=0.42u w=1.28u m=1
.ends oai321d2
* SPICE INPUT		Mon Sep 24 12:39:48 2018	oai322d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai322d0
.subckt oai322d0 B0 C1 A2 A1 C0 A0 B1 VDD GND Y
M1 N_10 B1 N_12 GND mn5  l=0.5u w=0.6u m=1
M2 N_10 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 C0 Y GND mn5  l=0.5u w=0.6u m=1
M4 GND A1 N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A2 GND GND mn5  l=0.5u w=0.6u m=1
M6 Y C1 N_12 GND mn5  l=0.5u w=0.6u m=1
M7 N_12 B0 N_10 GND mn5  l=0.5u w=0.6u m=1
M8 Y B1 N_9 VDD mp5  l=0.42u w=0.62u m=1
M9 N_15 C0 Y VDD mp5  l=0.42u w=0.62u m=1
M10 N_15 C1 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_17 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_9 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_17 A1 N_16 VDD mp5  l=0.42u w=0.62u m=1
M14 N_16 A2 Y VDD mp5  l=0.42u w=0.62u m=1
.ends oai322d0
* SPICE INPUT		Mon Sep 24 12:39:56 2018	oai322d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai322d1
.subckt oai322d1 B0 C1 A2 A0 C0 A1 B1 VDD Y GND
M1 N_14 B1 N_9 GND mn5  l=0.5u w=0.72u m=1
M2 GND A1 N_14 GND mn5  l=0.5u w=0.72u m=1
M3 N_9 C0 Y GND mn5  l=0.5u w=0.72u m=1
M4 N_14 A0 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_14 A2 GND GND mn5  l=0.5u w=0.72u m=1
M6 Y C1 N_9 GND mn5  l=0.5u w=0.72u m=1
M7 N_9 B0 N_14 GND mn5  l=0.5u w=0.72u m=1
M8 N_10 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M9 N_15 C0 Y VDD mp5  l=0.42u w=0.96u m=1
M10 N_15 C1 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 N_17 A1 N_16 VDD mp5  l=0.42u w=0.96u m=1
M12 N_10 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M13 N_17 A0 VDD VDD mp5  l=0.42u w=0.96u m=1
M14 N_16 A2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai322d1
* SPICE INPUT		Mon Sep 24 12:40:04 2018	oai322d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai322d2
.subckt oai322d2 Y VDD GND C0 B1 A2 C1 A1 A0 B0
M1 N_18 B1 N_16 GND mn5  l=0.5u w=0.98u m=1
M2 Y C1 N_16 GND mn5  l=0.5u w=0.98u m=1
M3 GND A0 N_18 GND mn5  l=0.5u w=0.98u m=1
M4 GND A1 N_18 GND mn5  l=0.5u w=0.98u m=1
M5 GND A2 N_18 GND mn5  l=0.5u w=0.98u m=1
M6 N_16 C0 Y GND mn5  l=0.5u w=0.98u m=1
M7 N_16 B0 N_18 GND mn5  l=0.5u w=0.98u m=1
M8 N_3 B1 Y VDD mp5  l=0.42u w=1.28u m=1
M9 N_9 C1 VDD VDD mp5  l=0.42u w=1.28u m=1
M10 N_9 C0 Y VDD mp5  l=0.42u w=1.28u m=1
M11 N_11 A0 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 N_3 B0 VDD VDD mp5  l=0.42u w=1.28u m=1
M13 N_11 A1 N_10 VDD mp5  l=0.42u w=1.28u m=1
M14 N_10 A2 Y VDD mp5  l=0.42u w=1.28u m=1
.ends oai322d2
* SPICE INPUT		Mon Sep 24 12:40:13 2018	oai32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d0
.subckt oai32d0 A2 B1 B0 A1 A0 GND VDD Y
M1 GND A0 N_10 GND mn5  l=0.5u w=0.6u m=1
M2 N_10 A1 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_10 B0 Y GND mn5  l=0.5u w=0.6u m=1
M4 N_10 B1 Y GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A2 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_13 A0 N_12 VDD mp5  l=0.42u w=0.62u m=1
M7 N_13 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 VDD B0 N_11 VDD mp5  l=0.42u w=0.62u m=1
M9 Y B1 N_11 VDD mp5  l=0.42u w=0.62u m=1
M10 N_12 A2 Y VDD mp5  l=0.42u w=0.62u m=1
.ends oai32d0
* SPICE INPUT		Mon Sep 24 12:40:21 2018	oai32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d1
.subckt oai32d1 B1 A2 A0 A1 B0 Y VDD GND
M1 N_9 B0 Y GND mn5  l=0.5u w=0.72u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 GND A0 N_9 GND mn5  l=0.5u w=0.72u m=1
M4 GND A2 N_9 GND mn5  l=0.5u w=0.72u m=1
M5 N_9 B1 Y GND mn5  l=0.5u w=0.72u m=1
M6 VDD B0 N_11 VDD mp5  l=0.42u w=0.96u m=1
M7 N_13 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_13 A0 N_12 VDD mp5  l=0.42u w=0.96u m=1
M9 N_12 A2 Y VDD mp5  l=0.42u w=0.96u m=1
M10 Y B1 N_11 VDD mp5  l=0.42u w=0.96u m=1
.ends oai32d1
* SPICE INPUT		Mon Sep 24 12:40:30 2018	oai32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d2
.subckt oai32d2 B1 A2 A0 A1 B0 Y VDD GND
M1 N_9 B0 Y GND mn5  l=0.5u w=0.98u m=1
M2 N_9 A1 GND GND mn5  l=0.5u w=0.98u m=1
M3 GND A0 N_9 GND mn5  l=0.5u w=0.98u m=1
M4 N_9 A2 GND GND mn5  l=0.5u w=0.98u m=1
M5 N_9 B1 Y GND mn5  l=0.5u w=0.98u m=1
M6 VDD B0 N_11 VDD mp5  l=0.42u w=1.28u m=1
M7 N_13 A1 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 N_13 A0 N_12 VDD mp5  l=0.42u w=1.28u m=1
M9 N_12 A2 Y VDD mp5  l=0.42u w=1.28u m=1
M10 Y B1 N_11 VDD mp5  l=0.42u w=1.28u m=1
.ends oai32d2
* SPICE INPUT		Mon Sep 24 12:40:38 2018	oai33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d0
.subckt oai33d0 A2 A0 B0 B2 A1 B1 Y VDD GND
M1 Y B1 N_8 GND mn5  l=0.5u w=0.6u m=1
M2 N_8 A1 GND GND mn5  l=0.5u w=0.6u m=1
M3 Y B2 N_8 GND mn5  l=0.5u w=0.6u m=1
M4 Y B0 N_8 GND mn5  l=0.5u w=0.6u m=1
M5 N_8 A0 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_8 A2 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_15 B1 N_12 VDD mp5  l=0.42u w=0.62u m=1
M8 N_14 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y B2 N_12 VDD mp5  l=0.42u w=0.62u m=1
M10 N_15 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_14 A0 N_13 VDD mp5  l=0.42u w=0.62u m=1
M12 N_13 A2 Y VDD mp5  l=0.42u w=0.62u m=1
.ends oai33d0
* SPICE INPUT		Mon Sep 24 12:40:47 2018	oai33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d1
.subckt oai33d1 A2 A0 B0 B2 A1 B1 Y VDD GND
M1 Y B1 N_8 GND mn5  l=0.5u w=0.72u m=1
M2 N_8 A1 GND GND mn5  l=0.5u w=0.72u m=1
M3 Y B2 N_8 GND mn5  l=0.5u w=0.72u m=1
M4 Y B0 N_8 GND mn5  l=0.5u w=0.72u m=1
M5 GND A0 N_8 GND mn5  l=0.5u w=0.72u m=1
M6 N_8 A2 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_15 B1 N_12 VDD mp5  l=0.42u w=0.96u m=1
M8 N_14 A1 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 Y B2 N_12 VDD mp5  l=0.42u w=0.96u m=1
M10 N_15 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M11 N_14 A0 N_13 VDD mp5  l=0.42u w=0.96u m=1
M12 N_13 A2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oai33d1
* SPICE INPUT		Mon Sep 24 12:40:55 2018	oai33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d2
.subckt oai33d2 Y VDD GND A1 A2 B2 B0 B1 A0
M1 Y B1 N_13 GND mn5  l=0.5u w=0.98u m=1
M2 N_13 A1 GND GND mn5  l=0.5u w=0.98u m=1
M3 Y B2 N_13 GND mn5  l=0.5u w=0.98u m=1
M4 Y B0 N_13 GND mn5  l=0.5u w=0.98u m=1
M5 GND A0 N_13 GND mn5  l=0.5u w=0.98u m=1
M6 N_13 A2 GND GND mn5  l=0.5u w=0.98u m=1
M7 N_9 B1 N_6 VDD mp5  l=0.42u w=1.28u m=1
M8 N_8 A1 VDD VDD mp5  l=0.42u w=1.28u m=1
M9 Y B2 N_6 VDD mp5  l=0.42u w=1.28u m=1
M10 N_9 B0 VDD VDD mp5  l=0.42u w=1.28u m=1
M11 N_8 A0 N_7 VDD mp5  l=0.42u w=1.28u m=1
M12 N_7 A2 Y VDD mp5  l=0.42u w=1.28u m=1
.ends oai33d2
* SPICE INPUT		Mon Sep 24 12:41:03 2018	oaim211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim211d0
.subckt oaim211d0 C0 B0 A0N A1N GND VDD Y
M1 N_11 A1N N_4 GND mn5  l=0.5u w=0.6u m=1
M2 N_11 A0N GND GND mn5  l=0.5u w=0.6u m=1
M3 N_12 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_12 B0 N_10 GND mn5  l=0.5u w=0.6u m=1
M5 Y C0 N_10 GND mn5  l=0.5u w=0.6u m=1
M6 N_4 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_4 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends oaim211d0
* SPICE INPUT		Mon Sep 24 12:41:11 2018	oaim211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim211d1
.subckt oaim211d1 B0 A0N C0 A1N Y GND VDD
M1 N_15 A1N N_3 GND mn5  l=0.5u w=0.6u m=1
M2 Y C0 N_14 GND mn5  l=0.5u w=0.72u m=1
M3 N_15 A0N GND GND mn5  l=0.5u w=0.6u m=1
M4 N_16 N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_16 B0 N_14 GND mn5  l=0.5u w=0.72u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_3 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y B0 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oaim211d1
* SPICE INPUT		Mon Sep 24 12:41:20 2018	oaim211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim211d2
.subckt oaim211d2 C0 A0N B0 A1N Y GND VDD
M1 N_11 A1N N_3 GND mn5  l=0.5u w=0.6u m=1
M2 N_12 B0 N_10 GND mn5  l=0.5u w=0.98u m=1
M3 N_11 A0N GND GND mn5  l=0.5u w=0.6u m=1
M4 N_12 N_3 GND GND mn5  l=0.5u w=0.98u m=1
M5 Y C0 N_10 GND mn5  l=0.5u w=0.98u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y B0 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 N_3 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends oaim211d2
* SPICE INPUT		Mon Sep 24 12:41:28 2018	oaim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d0
.subckt oaim21d0 B0 A1N A0N GND VDD Y
M1 N_10 A0N N_3 GND mn5  l=0.5u w=0.6u m=1
M2 N_10 A1N GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_3 N_9 GND mn5  l=0.5u w=0.6u m=1
M4 GND B0 N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_3 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_3 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
M7 Y N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 VDD B0 Y VDD mp5  l=0.42u w=0.62u m=1
.ends oaim21d0
* SPICE INPUT		Mon Sep 24 12:41:36 2018	oaim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d1
.subckt oaim21d1 A1N B0 A0N VDD Y GND
M1 N_10 A0N N_2 GND mn5  l=0.5u w=0.6u m=1
M2 GND B0 N_9 GND mn5  l=0.5u w=0.72u m=1
M3 N_10 A1N GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_2 N_9 GND mn5  l=0.5u w=0.72u m=1
M5 N_2 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M6 VDD B0 Y VDD mp5  l=0.42u w=0.96u m=1
M7 N_2 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
M8 VDD N_2 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oaim21d1
* SPICE INPUT		Mon Sep 24 12:41:45 2018	oaim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d2
.subckt oaim21d2 B0 A1N A0N VDD Y GND
M1 N_10 A0N N_2 GND mn5  l=0.5u w=0.6u m=1
M2 N_10 A1N GND GND mn5  l=0.5u w=0.6u m=1
M3 GND B0 N_9 GND mn5  l=0.5u w=0.98u m=1
M4 Y N_2 N_9 GND mn5  l=0.5u w=0.98u m=1
M5 N_2 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_2 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
M7 VDD B0 Y VDD mp5  l=0.42u w=1.28u m=1
M8 VDD N_2 Y VDD mp5  l=0.42u w=1.28u m=1
.ends oaim21d2
* SPICE INPUT		Mon Sep 24 12:41:53 2018	oaim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d0
.subckt oaim22d0 A1N A0N B0 B1 GND VDD Y
M1 Y N_6 N_10 GND mn5  l=0.5u w=0.6u m=1
M2 N_10 B1 GND GND mn5  l=0.5u w=0.6u m=1
M3 GND B0 N_10 GND mn5  l=0.5u w=0.6u m=1
M4 N_6 A0N N_19 GND mn5  l=0.5u w=0.6u m=1
M5 GND A1N N_19 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_11 B1 Y VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
.ends oaim22d0
* SPICE INPUT		Mon Sep 24 12:42:01 2018	oaim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d1
.subckt oaim22d1 A1N A0N B0 B1 GND VDD Y
M1 Y N_6 N_10 GND mn5  l=0.5u w=0.72u m=1
M2 N_10 B1 GND GND mn5  l=0.5u w=0.72u m=1
M3 GND B0 N_10 GND mn5  l=0.5u w=0.72u m=1
M4 N_6 A0N N_11 GND mn5  l=0.5u w=0.6u m=1
M5 GND A1N N_11 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_19 B1 Y VDD mp5  l=0.42u w=0.96u m=1
M8 N_19 B0 VDD VDD mp5  l=0.42u w=0.96u m=1
M9 N_6 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
.ends oaim22d1
* SPICE INPUT		Mon Sep 24 12:42:10 2018	oaim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d2
.subckt oaim22d2 A1N A0N B0 B1 GND VDD Y
M1 GND B1 N_10 GND mn5  l=0.5u w=0.98u m=1
M2 GND B0 N_10 GND mn5  l=0.5u w=0.98u m=1
M3 Y N_4 N_10 GND mn5  l=0.5u w=0.98u m=1
M4 N_4 A0N N_11 GND mn5  l=0.5u w=0.6u m=1
M5 N_11 A1N GND GND mn5  l=0.5u w=0.6u m=1
M6 N_19 B1 Y VDD mp5  l=0.42u w=1.28u m=1
M7 N_19 B0 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 Y N_4 VDD VDD mp5  l=0.42u w=1.28u m=1
M9 N_4 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_4 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
.ends oaim22d2
* SPICE INPUT		Mon Sep 24 12:42:18 2018	oaim2m11d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim2m11d0
.subckt oaim2m11d0 B0N A1N A0N C0 Y VDD GND
M1 GND N_6 N_11 GND mn5  l=0.5u w=0.6u m=1
M2 Y C0 N_11 GND mn5  l=0.5u w=0.6u m=1
M3 N_12 A0N N_6 GND mn5  l=0.5u w=0.6u m=1
M4 N_12 A1N GND GND mn5  l=0.5u w=0.6u m=1
M5 N_6 B0N GND GND mn5  l=0.5u w=0.6u m=1
M6 VDD A0N N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 VDD A1N N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 B0N N_10 VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y C0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends oaim2m11d0
* SPICE INPUT		Mon Sep 24 12:42:27 2018	oaim2m11d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim2m11d1
.subckt oaim2m11d1 B0N A1N A0N C0 GND VDD Y
M1 Y C0 N_11 GND mn5  l=0.5u w=0.72u m=1
M2 GND N_5 N_11 GND mn5  l=0.5u w=0.72u m=1
M3 N_12 A0N N_5 GND mn5  l=0.5u w=0.6u m=1
M4 N_12 A1N GND GND mn5  l=0.5u w=0.6u m=1
M5 N_5 B0N GND GND mn5  l=0.5u w=0.6u m=1
M6 VDD A0N N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 VDD A1N N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 B0N N_10 VDD mp5  l=0.42u w=0.62u m=1
M9 Y C0 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends oaim2m11d1
* SPICE INPUT		Mon Sep 24 12:42:34 2018	oaim2m11d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim2m11d2
.subckt oaim2m11d2 B0N A1N A0N C0 GND VDD Y
M1 Y C0 N_17 GND mn5  l=0.5u w=0.98u m=1
M2 GND N_5 N_17 GND mn5  l=0.5u w=0.98u m=1
M3 N_18 A0N N_5 GND mn5  l=0.5u w=0.6u m=1
M4 N_18 A1N GND GND mn5  l=0.5u w=0.6u m=1
M5 N_5 B0N GND GND mn5  l=0.5u w=0.6u m=1
M6 VDD A0N N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 VDD A1N N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 B0N N_10 VDD mp5  l=0.42u w=0.62u m=1
M9 Y C0 VDD VDD mp5  l=0.42u w=1.28u m=1
M10 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends oaim2m11d2
* SPICE INPUT		Mon Sep 24 12:42:42 2018	oaim31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim31d0
.subckt oaim31d0 B0 A2N A1N A0N Y GND VDD
M1 Y N_6 N_10 GND mn5  l=0.5u w=0.6u m=1
M2 N_11 A0N N_6 GND mn5  l=0.5u w=0.6u m=1
M3 N_12 A1N N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_12 A2N GND GND mn5  l=0.5u w=0.6u m=1
M5 GND B0 N_10 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_6 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 A2N VDD VDD mp5  l=0.42u w=0.62u m=1
M10 VDD B0 Y VDD mp5  l=0.42u w=0.62u m=1
.ends oaim31d0
* SPICE INPUT		Mon Sep 24 12:42:50 2018	oaim31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim31d1
.subckt oaim31d1 B0 A2N A1N A0N Y GND VDD
M1 Y N_6 N_10 GND mn5  l=0.5u w=0.72u m=1
M2 N_11 A0N N_6 GND mn5  l=0.5u w=0.6u m=1
M3 N_12 A1N N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_12 A2N GND GND mn5  l=0.5u w=0.6u m=1
M5 GND B0 N_10 GND mn5  l=0.5u w=0.72u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_6 A0N VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 A2N VDD VDD mp5  l=0.42u w=0.62u m=1
M10 VDD B0 Y VDD mp5  l=0.42u w=0.96u m=1
.ends oaim31d1
* SPICE INPUT		Mon Sep 24 12:42:58 2018	oaim31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim31d2
.subckt oaim31d2 Y GND VDD B0 A2N A1N A0N
M1 Y N_3 N_6 GND mn5  l=0.5u w=0.98u m=1
M2 N_7 A0N N_3 GND mn5  l=0.5u w=0.6u m=1
M3 N_8 A1N N_7 GND mn5  l=0.5u w=0.6u m=1
M4 N_8 A2N GND GND mn5  l=0.5u w=0.6u m=1
M5 GND B0 N_6 GND mn5  l=0.5u w=0.98u m=1
M6 Y N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 VDD A0N N_3 VDD mp5  l=0.42u w=0.62u m=1
M8 N_3 A1N VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_3 A2N VDD VDD mp5  l=0.42u w=0.62u m=1
M10 VDD B0 Y VDD mp5  l=0.42u w=1.28u m=1
.ends oaim31d2
* SPICE INPUT		Mon Sep 24 12:43:07 2018	or02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d0
.subckt or02d0 B A Y GND VDD
M1 Y N_4 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_4 A GND GND mn5  l=0.5u w=0.6u m=1
M3 N_4 B GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M5 N_8 A VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_8 B N_4 VDD mp5  l=0.42u w=0.62u m=1
.ends or02d0
* SPICE INPUT		Mon Sep 24 12:43:15 2018	or02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d1
.subckt or02d1 A B GND VDD Y
M1 N_2 B GND GND mn5  l=0.5u w=0.6u m=1
M2 N_2 A GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_8 B N_2 VDD mp5  l=0.42u w=0.62u m=1
M5 N_8 A VDD VDD mp5  l=0.42u w=0.62u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends or02d1
* SPICE INPUT		Mon Sep 24 12:43:24 2018	or02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d2
.subckt or02d2 A B GND VDD Y
M1 N_2 B GND GND mn5  l=0.5u w=0.6u m=1
M2 N_2 A GND GND mn5  l=0.5u w=0.6u m=1
M3 Y N_2 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_8 B N_2 VDD mp5  l=0.42u w=0.62u m=1
M5 N_8 A VDD VDD mp5  l=0.42u w=0.62u m=1
M6 Y N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends or02d2
* SPICE INPUT		Mon Sep 24 12:43:33 2018	or03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d0
.subckt or03d0 C B A GND Y VDD
M1 Y N_5 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 B GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 C GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_10 A VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_10 B N_9 VDD mp5  l=0.42u w=0.62u m=1
M8 N_9 C N_5 VDD mp5  l=0.42u w=0.62u m=1
.ends or03d0
* SPICE INPUT		Mon Sep 24 12:43:42 2018	or03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d1
.subckt or03d1 C B A GND VDD Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 B GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 C GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_10 A VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_10 B N_9 VDD mp5  l=0.42u w=0.62u m=1
M8 N_9 C N_5 VDD mp5  l=0.42u w=0.62u m=1
.ends or03d1
* SPICE INPUT		Mon Sep 24 12:43:50 2018	or03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d2
.subckt or03d2 C B A GND VDD Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_5 A GND GND mn5  l=0.5u w=0.6u m=1
M3 N_5 B GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 C GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M6 N_10 A VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_10 B N_9 VDD mp5  l=0.42u w=0.62u m=1
M8 N_9 C N_5 VDD mp5  l=0.42u w=0.62u m=1
.ends or03d2
* SPICE INPUT		Mon Sep 24 12:43:59 2018	or04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d0
.subckt or04d0 D A B C GND VDD Y
M1 N_3 C GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 B GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 A GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_3 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_11 C N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 N_12 B N_11 VDD mp5  l=0.42u w=0.62u m=1
M8 N_12 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_10 D N_3 VDD mp5  l=0.42u w=0.62u m=1
.ends or04d0
* SPICE INPUT		Mon Sep 24 12:44:08 2018	or04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d1
.subckt or04d1 D A B C GND VDD Y
M1 N_3 C GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 B GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 A GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M5 N_3 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_11 C N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 N_12 B N_11 VDD mp5  l=0.42u w=0.62u m=1
M8 N_12 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M10 N_10 D N_3 VDD mp5  l=0.42u w=0.62u m=1
.ends or04d1
* SPICE INPUT		Mon Sep 24 12:44:16 2018	or04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d2
.subckt or04d2 A B C D GND VDD Y
M1 N_3 D GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 C GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 B GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_3 GND GND mn5  l=0.5u w=0.98u m=1
M5 N_3 A GND GND mn5  l=0.5u w=0.6u m=1
M6 N_10 D N_3 VDD mp5  l=0.42u w=0.62u m=1
M7 N_11 C N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_12 B N_11 VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M10 N_12 A VDD VDD mp5  l=0.42u w=0.62u m=1
.ends or04d2
* SPICE INPUT		Mon Sep 24 12:44:25 2018	or12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or12d0
.subckt or12d0 AN B GND Y VDD
M1 N_2 B GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_2 B N_9 VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 VDD N_3 N_9 VDD mp5  l=0.42u w=0.62u m=1
.ends or12d0
* SPICE INPUT		Mon Sep 24 12:44:33 2018	or12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or12d1
.subckt or12d1 AN B GND Y VDD
M1 N_2 B GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M5 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M6 N_2 B N_9 VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 VDD N_3 N_9 VDD mp5  l=0.42u w=0.62u m=1
.ends or12d1
* SPICE INPUT		Mon Sep 24 12:44:42 2018	or12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or12d2
.subckt or12d2 AN B GND Y VDD
M1 N_2 B GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M4 Y N_2 GND GND mn5  l=0.5u w=0.98u m=1
M5 Y N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
M6 N_2 B N_9 VDD mp5  l=0.42u w=0.62u m=1
M7 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M8 VDD N_3 N_9 VDD mp5  l=0.42u w=0.62u m=1
.ends or12d2
* SPICE INPUT		Mon Sep 24 12:44:51 2018	or13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or13d0
.subckt or13d0 AN B C Y GND VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_6 C GND GND mn5  l=0.5u w=0.6u m=1
M3 N_6 B GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_6 C N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 N_11 B N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends or13d0
* SPICE INPUT		Mon Sep 24 12:44:59 2018	or13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or13d1
.subckt or13d1 B AN C GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_6 C GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_6 B GND GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_6 C N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_11 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_11 B N_10 VDD mp5  l=0.42u w=0.62u m=1
.ends or13d1
* SPICE INPUT		Mon Sep 24 12:45:07 2018	or13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or13d2
.subckt or13d2 B AN C GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_6 C GND GND mn5  l=0.5u w=0.6u m=1
M3 N_3 AN GND GND mn5  l=0.5u w=0.6u m=1
M4 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_6 B GND GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_6 C N_10 VDD mp5  l=0.42u w=0.62u m=1
M8 N_3 AN VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_11 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_11 B N_10 VDD mp5  l=0.42u w=0.62u m=1
.ends or13d2
* SPICE INPUT		Mon Sep 24 12:45:16 2018	or23d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or23d0
.subckt or23d0 AN C BN GND Y VDD
M1 Y N_7 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_4 BN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_7 C GND GND mn5  l=0.5u w=0.6u m=1
M4 N_7 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 C N_11 VDD mp5  l=0.42u w=0.62u m=1
M8 N_12 N_4 N_11 VDD mp5  l=0.42u w=0.62u m=1
M9 VDD AN N_2 VDD mp5  l=0.42u w=0.62u m=1
M10 VDD N_2 N_12 VDD mp5  l=0.42u w=0.62u m=1
M11 Y N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 N_4 BN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends or23d0
* SPICE INPUT		Mon Sep 24 12:45:25 2018	or23d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or23d1
.subckt or23d1 AN C BN GND Y VDD
M1 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_4 BN GND GND mn5  l=0.5u w=0.6u m=1
M3 GND C N_7 GND mn5  l=0.5u w=0.6u m=1
M4 N_7 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 C N_11 VDD mp5  l=0.42u w=0.62u m=1
M8 N_12 N_4 N_11 VDD mp5  l=0.42u w=0.62u m=1
M9 VDD AN N_2 VDD mp5  l=0.42u w=0.62u m=1
M10 VDD N_2 N_12 VDD mp5  l=0.42u w=0.62u m=1
M11 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_4 BN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends or23d1
* SPICE INPUT		Mon Sep 24 12:45:34 2018	or23d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or23d2
.subckt or23d2 AN C BN GND Y VDD
M1 Y N_7 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_4 BN GND GND mn5  l=0.5u w=0.6u m=1
M3 GND C N_7 GND mn5  l=0.5u w=0.6u m=1
M4 N_7 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 AN GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 C N_11 VDD mp5  l=0.42u w=0.62u m=1
M8 N_12 N_4 N_11 VDD mp5  l=0.42u w=0.62u m=1
M9 VDD AN N_2 VDD mp5  l=0.42u w=0.62u m=1
M10 VDD N_2 N_12 VDD mp5  l=0.42u w=0.62u m=1
M11 Y N_7 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 N_4 BN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends or23d2
* SPICE INPUT		Mon Sep 24 12:45:42 2018	ora211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d0
.subckt ora211d0 A1 A0 C0 B0 GND Y VDD
M1 Y N_6 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_8 B0 N_19 GND mn5  l=0.5u w=0.6u m=1
M3 N_19 C0 N_6 GND mn5  l=0.5u w=0.6u m=1
M4 N_8 A0 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_8 A1 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_6 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 VDD C0 N_6 VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 A1 N_11 VDD mp5  l=0.42u w=0.62u m=1
M10 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends ora211d0
* SPICE INPUT		Mon Sep 24 12:45:51 2018	ora211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d1
.subckt ora211d1 C0 B0 A1 A0 GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_10 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_10 A1 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_10 B0 N_19 GND mn5  l=0.5u w=0.6u m=1
M5 N_6 C0 N_19 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_11 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 A1 N_11 VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 C0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends ora211d1
* SPICE INPUT		Mon Sep 24 12:45:59 2018	ora211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d2
.subckt ora211d2 C0 B0 A1 A0 GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_10 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_10 A1 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_10 B0 N_19 GND mn5  l=0.5u w=0.6u m=1
M5 N_6 C0 N_19 GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_11 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 A1 N_11 VDD mp5  l=0.42u w=0.62u m=1
M9 N_6 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 C0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends ora211d2
* SPICE INPUT		Mon Sep 24 12:46:08 2018	ora21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d0
.subckt ora21d0 B0 A0 A1 VDD GND Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A1 N_8 GND mn5  l=0.5u w=0.6u m=1
M3 N_8 A0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 B0 N_8 GND mn5  l=0.5u w=0.6u m=1
M5 N_5 A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M6 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_5 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends ora21d0
* SPICE INPUT		Mon Sep 24 12:46:16 2018	ora21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d1
.subckt ora21d1 B0 A0 A1 VDD GND Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.72u m=1
M2 GND A1 N_8 GND mn5  l=0.5u w=0.6u m=1
M3 N_8 A0 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_5 B0 N_8 GND mn5  l=0.5u w=0.6u m=1
M5 N_5 A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M6 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_5 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends ora21d1
* SPICE INPUT		Mon Sep 24 12:46:25 2018	ora21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d2
.subckt ora21d2 B0 A1 A0 GND VDD Y
M1 Y N_5 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_9 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 GND A1 N_9 GND mn5  l=0.5u w=0.6u m=1
M4 N_5 B0 N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M6 N_5 A1 N_10 VDD mp5  l=0.42u w=0.62u m=1
M7 N_5 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 Y N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends ora21d2
* SPICE INPUT		Mon Sep 24 12:46:33 2018	ora311d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora311d1
.subckt ora311d1 C0 A1 B0 A2 A0 Y GND VDD
M1 Y N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_8 A2 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_8 B0 N_21 GND mn5  l=0.5u w=0.6u m=1
M5 N_8 A1 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 C0 N_21 GND mn5  l=0.5u w=0.6u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M8 N_12 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_7 A2 N_13 VDD mp5  l=0.42u w=0.62u m=1
M10 N_7 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_13 A1 N_12 VDD mp5  l=0.42u w=0.62u m=1
M12 N_7 C0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends ora311d1
* SPICE INPUT		Mon Sep 24 12:46:42 2018	ora311d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora311d2
.subckt ora311d2 C0 A1 B0 A2 A0 Y GND VDD
M1 Y N_7 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_8 A0 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_8 A2 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_8 B0 N_21 GND mn5  l=0.5u w=0.6u m=1
M5 N_8 A1 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 C0 N_21 GND mn5  l=0.5u w=0.6u m=1
M7 Y N_7 VDD VDD mp5  l=0.42u w=1.28u m=1
M8 N_12 A0 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_7 A2 N_13 VDD mp5  l=0.42u w=0.62u m=1
M10 N_7 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M11 N_13 A1 N_12 VDD mp5  l=0.42u w=0.62u m=1
M12 N_7 C0 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends ora311d2
* SPICE INPUT		Mon Sep 24 12:46:51 2018	ora31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d0
.subckt ora31d0 A2 A1 A0 B0 VDD Y GND
M1 Y N_6 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_6 B0 N_10 GND mn5  l=0.5u w=0.6u m=1
M3 GND A0 N_10 GND mn5  l=0.5u w=0.6u m=1
M4 N_10 A1 GND GND mn5  l=0.5u w=0.6u m=1
M5 GND A2 N_10 GND mn5  l=0.5u w=0.6u m=1
M6 N_6 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M7 N_12 A0 N_11 VDD mp5  l=0.42u w=0.62u m=1
M8 N_11 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M9 Y N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_6 A2 N_12 VDD mp5  l=0.42u w=0.62u m=1
.ends ora31d0
* SPICE INPUT		Mon Sep 24 12:46:59 2018	ora31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d1
.subckt ora31d1 A0 A1 A2 B0 GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_6 B0 N_10 GND mn5  l=0.5u w=0.6u m=1
M3 GND A2 N_10 GND mn5  l=0.5u w=0.6u m=1
M4 N_10 A1 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A0 GND GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M7 N_6 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 A2 N_12 VDD mp5  l=0.42u w=0.62u m=1
M9 N_11 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_12 A0 N_11 VDD mp5  l=0.42u w=0.62u m=1
.ends ora31d1
* SPICE INPUT		Mon Sep 24 12:47:08 2018	ora31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d2
.subckt ora31d2 A0 A1 A2 B0 GND VDD Y
M1 Y N_6 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_6 B0 N_10 GND mn5  l=0.5u w=0.6u m=1
M3 GND A2 N_10 GND mn5  l=0.5u w=0.6u m=1
M4 N_10 A1 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_10 A0 GND GND mn5  l=0.5u w=0.6u m=1
M6 Y N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M7 N_6 B0 VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_6 A2 N_12 VDD mp5  l=0.42u w=0.62u m=1
M9 N_11 A1 VDD VDD mp5  l=0.42u w=0.62u m=1
M10 N_12 A0 N_11 VDD mp5  l=0.42u w=0.62u m=1
.ends ora31d2
* SPICE INPUT		Mon Sep 24 12:47:17 2018	sdbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb1
.subckt sdbfb1 VDD Q QN GND RN SN SI SE D CKN
M1 Q N_19 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_10 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_20 RN GND GND mn5  l=0.5u w=0.6u m=1
M4 GND N_10 N_19 GND mn5  l=0.5u w=0.6u m=1
M5 N_4 N_12 N_36 GND mn5  l=0.5u w=0.6u m=1
M6 N_4 N_13 N_68 GND mn5  l=0.5u w=0.6u m=1
M7 N_68 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_16 SE GND GND mn5  l=0.5u w=0.6u m=1
M9 N_70 D GND GND mn5  l=0.5u w=0.6u m=1
M10 N_36 N_16 N_70 GND mn5  l=0.5u w=0.6u m=1
M11 N_36 SI N_69 GND mn5  l=0.5u w=0.6u m=1
M12 N_69 SE GND GND mn5  l=0.5u w=0.6u m=1
M13 N_13 CKN GND GND mn5  l=0.5u w=0.6u m=1
M14 GND N_13 N_12 GND mn5  l=0.5u w=0.6u m=1
M15 N_6 N_4 N_35 GND mn5  l=0.5u w=0.6u m=1
M16 N_6 N_20 N_35 GND mn5  l=0.5u w=0.6u m=1
M17 GND SN N_35 GND mn5  l=0.5u w=0.6u m=1
M18 N_71 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M19 N_8 N_13 N_71 GND mn5  l=0.5u w=0.6u m=1
M20 N_72 N_12 N_8 GND mn5  l=0.5u w=0.6u m=1
M21 GND N_10 N_72 GND mn5  l=0.5u w=0.6u m=1
M22 N_33 SN GND GND mn5  l=0.5u w=0.6u m=1
M23 N_33 N_20 N_10 GND mn5  l=0.5u w=0.6u m=1
M24 N_33 N_8 N_10 GND mn5  l=0.5u w=0.6u m=1
M25 N_4 N_13 N_3 VDD mp5  l=0.42u w=0.62u m=1
M26 N_26 N_12 N_4 VDD mp5  l=0.42u w=0.62u m=1
M27 VDD N_6 N_26 VDD mp5  l=0.42u w=0.62u m=1
M28 N_27 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_27 N_20 N_6 VDD mp5  l=0.42u w=0.62u m=1
M30 VDD SN N_6 VDD mp5  l=0.42u w=0.62u m=1
M31 N_28 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_28 N_12 N_8 VDD mp5  l=0.42u w=0.62u m=1
M33 N_29 N_13 N_8 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD N_10 N_29 VDD mp5  l=0.42u w=0.6u m=1
M35 N_10 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_10 N_20 N_25 VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_8 N_25 VDD mp5  l=0.42u w=0.62u m=1
M38 N_13 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M39 N_12 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M40 N_16 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M41 N_31 D VDD VDD mp5  l=0.42u w=0.62u m=1
M42 N_3 SE N_31 VDD mp5  l=0.42u w=0.62u m=1
M43 N_3 N_16 N_30 VDD mp5  l=0.42u w=0.62u m=1
M44 N_30 SI VDD VDD mp5  l=0.42u w=0.62u m=1
M45 N_20 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M46 N_19 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M47 Q N_19 VDD VDD mp5  l=0.42u w=0.96u m=1
M48 QN N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdbfb1
* SPICE INPUT		Mon Sep 24 12:47:25 2018	sdbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb2
.subckt sdbfb2 VDD Q QN GND RN SN SI SE D CKN
M1 N_13 RN GND GND mn5  l=0.5u w=0.6u m=1
M2 GND N_10 N_12 GND mn5  l=0.5u w=0.6u m=1
M3 N_4 N_18 N_36 GND mn5  l=0.5u w=0.6u m=1
M4 N_4 N_19 N_68 GND mn5  l=0.5u w=0.6u m=1
M5 N_68 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_22 SE GND GND mn5  l=0.5u w=0.6u m=1
M7 N_70 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_36 N_22 N_70 GND mn5  l=0.5u w=0.6u m=1
M9 N_36 SI N_69 GND mn5  l=0.5u w=0.6u m=1
M10 N_69 SE GND GND mn5  l=0.5u w=0.6u m=1
M11 N_19 CKN GND GND mn5  l=0.5u w=0.6u m=1
M12 GND N_19 N_18 GND mn5  l=0.5u w=0.6u m=1
M13 N_6 N_4 N_35 GND mn5  l=0.5u w=0.6u m=1
M14 N_6 N_13 N_35 GND mn5  l=0.5u w=0.6u m=1
M15 GND SN N_35 GND mn5  l=0.5u w=0.6u m=1
M16 N_71 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M17 N_8 N_19 N_71 GND mn5  l=0.5u w=0.6u m=1
M18 N_72 N_18 N_8 GND mn5  l=0.5u w=0.6u m=1
M19 GND N_10 N_72 GND mn5  l=0.5u w=0.6u m=1
M20 N_33 SN GND GND mn5  l=0.5u w=0.6u m=1
M21 N_33 N_13 N_10 GND mn5  l=0.5u w=0.6u m=1
M22 N_33 N_8 N_10 GND mn5  l=0.5u w=0.6u m=1
M23 Q N_12 GND GND mn5  l=0.5u w=0.98u m=1
M24 QN N_10 GND GND mn5  l=0.5u w=0.98u m=1
M25 N_4 N_19 N_3 VDD mp5  l=0.42u w=0.62u m=1
M26 N_26 N_18 N_4 VDD mp5  l=0.42u w=0.62u m=1
M27 VDD N_6 N_26 VDD mp5  l=0.42u w=0.62u m=1
M28 N_27 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_27 N_13 N_6 VDD mp5  l=0.42u w=0.62u m=1
M30 VDD SN N_6 VDD mp5  l=0.42u w=0.62u m=1
M31 N_28 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_28 N_18 N_8 VDD mp5  l=0.42u w=0.62u m=1
M33 N_29 N_19 N_8 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD N_10 N_29 VDD mp5  l=0.42u w=0.6u m=1
M35 N_10 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_10 N_13 N_25 VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_8 N_25 VDD mp5  l=0.42u w=0.62u m=1
M38 N_13 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M39 N_12 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M40 Q N_12 VDD VDD mp5  l=0.42u w=1.28u m=1
M41 QN N_10 VDD VDD mp5  l=0.42u w=1.28u m=1
M42 N_19 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M43 N_18 N_19 VDD VDD mp5  l=0.42u w=0.62u m=1
M44 N_22 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M45 N_31 D VDD VDD mp5  l=0.42u w=0.62u m=1
M46 N_3 SE N_31 VDD mp5  l=0.42u w=0.62u m=1
M47 N_3 N_22 N_30 VDD mp5  l=0.42u w=0.62u m=1
M48 N_30 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdbfb2
* SPICE INPUT		Mon Sep 24 12:47:34 2018	sdbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb1
.subckt sdbrb1 VDD Q QN GND RN SN SI SE D CK
M1 N_13 RN GND GND mn5  l=0.5u w=0.6u m=1
M2 GND N_10 N_12 GND mn5  l=0.5u w=0.6u m=1
M3 N_3 N_18 N_36 GND mn5  l=0.5u w=0.6u m=1
M4 N_3 N_19 N_68 GND mn5  l=0.5u w=0.6u m=1
M5 N_68 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_22 SE GND GND mn5  l=0.5u w=0.6u m=1
M7 N_70 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_36 N_22 N_70 GND mn5  l=0.5u w=0.6u m=1
M9 N_36 SI N_69 GND mn5  l=0.5u w=0.6u m=1
M10 N_69 SE GND GND mn5  l=0.5u w=0.6u m=1
M11 N_19 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M12 GND CK N_18 GND mn5  l=0.5u w=0.6u m=1
M13 N_6 N_3 N_35 GND mn5  l=0.5u w=0.6u m=1
M14 N_6 N_13 N_35 GND mn5  l=0.5u w=0.6u m=1
M15 GND SN N_35 GND mn5  l=0.5u w=0.6u m=1
M16 N_71 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M17 N_8 N_19 N_71 GND mn5  l=0.5u w=0.6u m=1
M18 N_72 N_18 N_8 GND mn5  l=0.5u w=0.6u m=1
M19 GND N_10 N_72 GND mn5  l=0.5u w=0.6u m=1
M20 N_33 SN GND GND mn5  l=0.5u w=0.6u m=1
M21 N_33 N_13 N_10 GND mn5  l=0.5u w=0.6u m=1
M22 N_33 N_8 N_10 GND mn5  l=0.5u w=0.6u m=1
M23 Q N_12 GND GND mn5  l=0.5u w=0.72u m=1
M24 QN N_10 GND GND mn5  l=0.5u w=0.72u m=1
M25 N_4 N_19 N_3 VDD mp5  l=0.42u w=0.62u m=1
M26 N_26 N_18 N_3 VDD mp5  l=0.42u w=0.6u m=1
M27 VDD N_6 N_26 VDD mp5  l=0.42u w=0.6u m=1
M28 N_27 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_27 N_13 N_6 VDD mp5  l=0.42u w=0.62u m=1
M30 VDD SN N_6 VDD mp5  l=0.42u w=0.62u m=1
M31 N_28 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_28 N_18 N_8 VDD mp5  l=0.42u w=0.62u m=1
M33 N_29 N_19 N_8 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD N_10 N_29 VDD mp5  l=0.42u w=0.6u m=1
M35 N_10 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_10 N_13 N_25 VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_8 N_25 VDD mp5  l=0.42u w=0.62u m=1
M38 N_13 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M39 N_12 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M40 Q N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M41 QN N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
M42 N_19 N_18 VDD VDD mp5  l=0.42u w=0.62u m=1
M43 N_18 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M44 N_22 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M45 N_31 D VDD VDD mp5  l=0.42u w=0.62u m=1
M46 N_4 SE N_31 VDD mp5  l=0.42u w=0.62u m=1
M47 N_4 N_22 N_30 VDD mp5  l=0.42u w=0.62u m=1
M48 N_30 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdbrb1
* SPICE INPUT		Mon Sep 24 12:47:42 2018	sdbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb2
.subckt sdbrb2 VDD Q QN GND RN SN SI SE D CK
M1 N_13 RN GND GND mn5  l=0.5u w=0.6u m=1
M2 GND N_10 N_12 GND mn5  l=0.5u w=0.6u m=1
M3 N_3 N_18 N_36 GND mn5  l=0.5u w=0.6u m=1
M4 N_3 N_19 N_68 GND mn5  l=0.5u w=0.6u m=1
M5 N_68 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_22 SE GND GND mn5  l=0.5u w=0.6u m=1
M7 N_70 D GND GND mn5  l=0.5u w=0.6u m=1
M8 N_36 N_22 N_70 GND mn5  l=0.5u w=0.6u m=1
M9 N_36 SI N_69 GND mn5  l=0.5u w=0.6u m=1
M10 N_69 SE GND GND mn5  l=0.5u w=0.6u m=1
M11 N_19 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M12 GND CK N_18 GND mn5  l=0.5u w=0.6u m=1
M13 N_6 N_3 N_35 GND mn5  l=0.5u w=0.6u m=1
M14 N_6 N_13 N_35 GND mn5  l=0.5u w=0.6u m=1
M15 GND SN N_35 GND mn5  l=0.5u w=0.6u m=1
M16 N_71 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M17 N_8 N_19 N_71 GND mn5  l=0.5u w=0.6u m=1
M18 N_72 N_18 N_8 GND mn5  l=0.5u w=0.6u m=1
M19 GND N_10 N_72 GND mn5  l=0.5u w=0.6u m=1
M20 N_33 SN GND GND mn5  l=0.5u w=0.6u m=1
M21 N_33 N_13 N_10 GND mn5  l=0.5u w=0.6u m=1
M22 N_33 N_8 N_10 GND mn5  l=0.5u w=0.6u m=1
M23 Q N_12 GND GND mn5  l=0.5u w=0.98u m=1
M24 QN N_10 GND GND mn5  l=0.5u w=0.98u m=1
M25 N_4 N_19 N_3 VDD mp5  l=0.42u w=0.62u m=1
M26 N_26 N_18 N_3 VDD mp5  l=0.42u w=0.6u m=1
M27 VDD N_6 N_26 VDD mp5  l=0.42u w=0.6u m=1
M28 N_27 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_27 N_13 N_6 VDD mp5  l=0.42u w=0.62u m=1
M30 VDD SN N_6 VDD mp5  l=0.42u w=0.62u m=1
M31 N_28 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_28 N_18 N_8 VDD mp5  l=0.42u w=0.62u m=1
M33 N_29 N_19 N_8 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD N_10 N_29 VDD mp5  l=0.42u w=0.6u m=1
M35 N_10 SN VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_10 N_13 N_25 VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_8 N_25 VDD mp5  l=0.42u w=0.62u m=1
M38 N_13 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M39 N_12 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M40 Q N_12 VDD VDD mp5  l=0.42u w=1.28u m=1
M41 QN N_10 VDD VDD mp5  l=0.42u w=1.28u m=1
M42 N_19 N_18 VDD VDD mp5  l=0.42u w=0.62u m=1
M43 N_18 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M44 N_22 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M45 N_31 D VDD VDD mp5  l=0.42u w=0.62u m=1
M46 N_4 SE N_31 VDD mp5  l=0.42u w=0.62u m=1
M47 N_4 N_22 N_30 VDD mp5  l=0.42u w=0.62u m=1
M48 N_30 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdbrb2
* SPICE INPUT		Mon Sep 24 12:47:51 2018	sdbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq1
.subckt sdbrq1 VDD Q GND D CK SE SI SN RN
M1 N_43 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_7 N_17 N_43 GND mn5  l=0.5u w=0.6u m=1
M3 N_7 N_16 N_37 GND mn5  l=0.5u w=0.6u m=1
M4 N_20 SE GND GND mn5  l=0.5u w=0.6u m=1
M5 N_45 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_37 N_20 N_45 GND mn5  l=0.5u w=0.6u m=1
M7 N_44 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_37 SI N_44 GND mn5  l=0.5u w=0.6u m=1
M9 GND CK N_16 GND mn5  l=0.5u w=0.6u m=1
M10 N_17 N_16 GND GND mn5  l=0.5u w=0.6u m=1
M11 GND SN N_41 GND mn5  l=0.5u w=0.6u m=1
M12 GND N_14 N_47 GND mn5  l=0.5u w=0.6u m=1
M13 N_41 N_3 N_14 GND mn5  l=0.5u w=0.6u m=1
M14 N_41 N_12 N_14 GND mn5  l=0.5u w=0.6u m=1
M15 N_12 N_17 N_46 GND mn5  l=0.5u w=0.6u m=1
M16 N_47 N_16 N_12 GND mn5  l=0.5u w=0.6u m=1
M17 GND SN N_40 GND mn5  l=0.5u w=0.6u m=1
M18 N_10 N_3 N_40 GND mn5  l=0.5u w=0.6u m=1
M19 N_10 N_7 N_40 GND mn5  l=0.5u w=0.6u m=1
M20 N_46 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M21 N_33 SN GND GND mn5  l=0.5u w=0.72u m=1
M22 N_33 N_3 Q GND mn5  l=0.5u w=0.72u m=1
M23 Q N_12 N_33 GND mn5  l=0.5u w=0.72u m=1
M24 N_3 RN GND GND mn5  l=0.5u w=0.6u m=1
M25 Q SN VDD VDD mp5  l=0.42u w=0.96u m=1
M26 Q N_3 N_23 VDD mp5  l=0.42u w=0.96u m=1
M27 N_23 N_12 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_3 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_27 N_16 N_12 VDD mp5  l=0.42u w=0.62u m=1
M30 N_14 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M31 VDD N_14 N_28 VDD mp5  l=0.42u w=0.6u m=1
M32 N_14 N_3 N_24 VDD mp5  l=0.42u w=0.6u m=1
M33 VDD N_12 N_24 VDD mp5  l=0.42u w=0.6u m=1
M34 N_28 N_17 N_12 VDD mp5  l=0.42u w=0.6u m=1
M35 VDD SN N_10 VDD mp5  l=0.42u w=0.62u m=1
M36 N_26 N_3 N_10 VDD mp5  l=0.42u w=0.62u m=1
M37 N_26 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M38 VDD N_10 N_25 VDD mp5  l=0.42u w=0.6u m=1
M39 N_25 N_16 N_7 VDD mp5  l=0.42u w=0.6u m=1
M40 N_27 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M41 N_8 N_17 N_7 VDD mp5  l=0.42u w=0.62u m=1
M42 N_16 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M43 N_17 N_16 VDD VDD mp5  l=0.42u w=0.62u m=1
M44 N_20 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M45 N_30 D VDD VDD mp5  l=0.42u w=0.62u m=1
M46 N_8 SE N_30 VDD mp5  l=0.42u w=0.62u m=1
M47 N_8 N_20 N_29 VDD mp5  l=0.42u w=0.62u m=1
M48 N_29 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdbrq1
* SPICE INPUT		Mon Sep 24 12:47:59 2018	sdbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq2
.subckt sdbrq2 VDD Q GND D CK SE SI SN RN
M1 N_43 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_7 N_17 N_43 GND mn5  l=0.5u w=0.6u m=1
M3 N_7 N_16 N_37 GND mn5  l=0.5u w=0.6u m=1
M4 N_20 SE GND GND mn5  l=0.5u w=0.6u m=1
M5 N_45 D GND GND mn5  l=0.5u w=0.6u m=1
M6 N_37 N_20 N_45 GND mn5  l=0.5u w=0.6u m=1
M7 N_44 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_37 SI N_44 GND mn5  l=0.5u w=0.6u m=1
M9 GND CK N_16 GND mn5  l=0.5u w=0.6u m=1
M10 N_17 N_16 GND GND mn5  l=0.5u w=0.6u m=1
M11 GND SN N_41 GND mn5  l=0.5u w=0.6u m=1
M12 GND N_14 N_47 GND mn5  l=0.5u w=0.6u m=1
M13 N_41 N_3 N_14 GND mn5  l=0.5u w=0.6u m=1
M14 N_41 N_12 N_14 GND mn5  l=0.5u w=0.6u m=1
M15 N_12 N_17 N_46 GND mn5  l=0.5u w=0.6u m=1
M16 N_47 N_16 N_12 GND mn5  l=0.5u w=0.6u m=1
M17 GND SN N_40 GND mn5  l=0.5u w=0.6u m=1
M18 N_10 N_3 N_40 GND mn5  l=0.5u w=0.6u m=1
M19 N_10 N_7 N_40 GND mn5  l=0.5u w=0.6u m=1
M20 N_46 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M21 N_33 SN GND GND mn5  l=0.5u w=0.98u m=1
M22 N_33 N_3 Q GND mn5  l=0.5u w=0.98u m=1
M23 Q N_12 N_33 GND mn5  l=0.5u w=0.98u m=1
M24 N_3 RN GND GND mn5  l=0.5u w=0.6u m=1
M25 Q SN VDD VDD mp5  l=0.42u w=1.28u m=1
M26 Q N_3 N_23 VDD mp5  l=0.42u w=1.28u m=1
M27 N_23 N_12 VDD VDD mp5  l=0.42u w=1.28u m=1
M28 N_3 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_27 N_16 N_12 VDD mp5  l=0.42u w=0.62u m=1
M30 N_14 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M31 VDD N_14 N_28 VDD mp5  l=0.42u w=0.6u m=1
M32 N_14 N_3 N_24 VDD mp5  l=0.42u w=0.6u m=1
M33 VDD N_12 N_24 VDD mp5  l=0.42u w=0.6u m=1
M34 N_28 N_17 N_12 VDD mp5  l=0.42u w=0.6u m=1
M35 VDD SN N_10 VDD mp5  l=0.42u w=0.62u m=1
M36 N_26 N_3 N_10 VDD mp5  l=0.42u w=0.62u m=1
M37 N_26 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M38 VDD N_10 N_25 VDD mp5  l=0.42u w=0.6u m=1
M39 N_25 N_16 N_7 VDD mp5  l=0.42u w=0.6u m=1
M40 N_27 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M41 N_8 N_17 N_7 VDD mp5  l=0.42u w=0.62u m=1
M42 N_16 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M43 N_17 N_16 VDD VDD mp5  l=0.42u w=0.62u m=1
M44 N_20 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M45 N_30 D VDD VDD mp5  l=0.42u w=0.62u m=1
M46 N_8 SE N_30 VDD mp5  l=0.42u w=0.62u m=1
M47 N_8 N_20 N_29 VDD mp5  l=0.42u w=0.62u m=1
M48 N_29 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdbrq2
* SPICE INPUT		Mon Sep 24 12:48:08 2018	sdcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb1
.subckt sdcfb1 VDD Q QN GND RN CKN SI SE D
M1 GND N_16 N_21 GND mn5  l=0.5u w=0.6u m=1
M2 N_22 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_7 SE GND GND mn5  l=0.5u w=0.6u m=1
M4 N_62 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_31 N_7 N_62 GND mn5  l=0.5u w=0.6u m=1
M6 N_61 SE GND GND mn5  l=0.5u w=0.6u m=1
M7 N_31 SI N_61 GND mn5  l=0.5u w=0.6u m=1
M8 GND N_4 N_3 GND mn5  l=0.5u w=0.6u m=1
M9 N_4 CKN GND GND mn5  l=0.5u w=0.6u m=1
M10 N_63 N_4 N_10 GND mn5  l=0.5u w=0.6u m=1
M11 N_63 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M12 GND N_22 N_16 GND mn5  l=0.5u w=0.6u m=1
M13 GND N_18 N_16 GND mn5  l=0.5u w=0.6u m=1
M14 GND N_16 N_65 GND mn5  l=0.5u w=0.6u m=1
M15 N_64 N_4 N_18 GND mn5  l=0.5u w=0.6u m=1
M16 N_65 N_3 N_18 GND mn5  l=0.5u w=0.6u m=1
M17 N_64 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M18 N_9 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M19 N_10 N_3 N_31 GND mn5  l=0.5u w=0.6u m=1
M20 N_9 N_22 GND GND mn5  l=0.5u w=0.6u m=1
M21 QN N_16 GND GND mn5  l=0.5u w=0.72u m=1
M22 Q N_21 GND GND mn5  l=0.5u w=0.72u m=1
M23 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_4 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_7 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M26 N_8 SE N_25 VDD mp5  l=0.42u w=0.62u m=1
M27 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_8 N_7 N_24 VDD mp5  l=0.42u w=0.62u m=1
M29 N_24 SI VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_8 N_4 N_10 VDD mp5  l=0.42u w=0.62u m=1
M31 VDD N_9 N_27 VDD mp5  l=0.42u w=0.6u m=1
M32 VDD N_10 N_26 VDD mp5  l=0.42u w=0.62u m=1
M33 N_27 N_3 N_10 VDD mp5  l=0.42u w=0.6u m=1
M34 N_9 N_22 N_26 VDD mp5  l=0.42u w=0.62u m=1
M35 QN N_16 VDD VDD mp5  l=0.42u w=0.96u m=1
M36 Q N_21 VDD VDD mp5  l=0.42u w=0.96u m=1
M37 N_16 N_22 N_28 VDD mp5  l=0.42u w=0.62u m=1
M38 VDD N_18 N_28 VDD mp5  l=0.42u w=0.62u m=1
M39 VDD N_16 N_30 VDD mp5  l=0.42u w=0.6u m=1
M40 N_30 N_4 N_18 VDD mp5  l=0.42u w=0.6u m=1
M41 N_29 N_3 N_18 VDD mp5  l=0.42u w=0.62u m=1
M42 N_29 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M43 N_21 N_16 VDD VDD mp5  l=0.42u w=0.6u m=1
M44 N_22 RN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdcfb1
* SPICE INPUT		Mon Sep 24 12:48:17 2018	sdcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb2
.subckt sdcfb2 VDD Q QN GND RN CKN SI SE D
M1 GND N_16 N_21 GND mn5  l=0.5u w=0.6u m=1
M2 N_22 RN GND GND mn5  l=0.5u w=0.6u m=1
M3 N_7 SE GND GND mn5  l=0.5u w=0.6u m=1
M4 N_62 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_31 N_7 N_62 GND mn5  l=0.5u w=0.6u m=1
M6 N_61 SE GND GND mn5  l=0.5u w=0.6u m=1
M7 N_31 SI N_61 GND mn5  l=0.5u w=0.6u m=1
M8 GND N_4 N_3 GND mn5  l=0.5u w=0.6u m=1
M9 N_4 CKN GND GND mn5  l=0.5u w=0.6u m=1
M10 N_63 N_4 N_10 GND mn5  l=0.5u w=0.6u m=1
M11 N_63 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M12 GND N_22 N_16 GND mn5  l=0.5u w=0.6u m=1
M13 GND N_18 N_16 GND mn5  l=0.5u w=0.6u m=1
M14 GND N_16 N_65 GND mn5  l=0.5u w=0.6u m=1
M15 N_64 N_4 N_18 GND mn5  l=0.5u w=0.6u m=1
M16 N_65 N_3 N_18 GND mn5  l=0.5u w=0.6u m=1
M17 N_64 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M18 N_9 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M19 N_10 N_3 N_31 GND mn5  l=0.5u w=0.6u m=1
M20 N_9 N_22 GND GND mn5  l=0.5u w=0.6u m=1
M21 QN N_16 GND GND mn5  l=0.5u w=0.98u m=1
M22 Q N_21 GND GND mn5  l=0.5u w=0.98u m=1
M23 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_4 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_7 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M26 N_8 SE N_25 VDD mp5  l=0.42u w=0.62u m=1
M27 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_8 N_7 N_24 VDD mp5  l=0.42u w=0.62u m=1
M29 N_24 SI VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_8 N_4 N_10 VDD mp5  l=0.42u w=0.62u m=1
M31 VDD N_9 N_27 VDD mp5  l=0.42u w=0.6u m=1
M32 VDD N_10 N_26 VDD mp5  l=0.42u w=0.62u m=1
M33 N_27 N_3 N_10 VDD mp5  l=0.42u w=0.6u m=1
M34 N_9 N_22 N_26 VDD mp5  l=0.42u w=0.62u m=1
M35 QN N_16 VDD VDD mp5  l=0.42u w=1.28u m=1
M36 Q N_21 VDD VDD mp5  l=0.42u w=1.28u m=1
M37 N_16 N_22 N_28 VDD mp5  l=0.42u w=0.62u m=1
M38 VDD N_18 N_28 VDD mp5  l=0.42u w=0.62u m=1
M39 VDD N_16 N_30 VDD mp5  l=0.42u w=0.6u m=1
M40 N_30 N_4 N_18 VDD mp5  l=0.42u w=0.6u m=1
M41 N_29 N_3 N_18 VDD mp5  l=0.42u w=0.62u m=1
M42 N_29 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M43 N_21 N_16 VDD VDD mp5  l=0.42u w=0.6u m=1
M44 N_22 RN VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdcfb2
* SPICE INPUT		Mon Sep 24 12:48:26 2018	sdcfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfq1
.subckt sdcfq1 VDD Q GND RN SI SE D CKN
M1 N_14 RN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_15 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_11 SE GND GND mn5  l=0.5u w=0.6u m=1
M4 N_38 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_31 N_11 N_38 GND mn5  l=0.5u w=0.6u m=1
M6 N_31 SI N_37 GND mn5  l=0.5u w=0.6u m=1
M7 N_37 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_8 CKN GND GND mn5  l=0.5u w=0.6u m=1
M9 GND N_8 N_7 GND mn5  l=0.5u w=0.6u m=1
M10 N_3 N_7 N_31 GND mn5  l=0.5u w=0.6u m=1
M11 N_39 N_8 N_3 GND mn5  l=0.5u w=0.6u m=1
M12 N_39 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_2 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_40 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_41 N_7 N_20 GND mn5  l=0.5u w=0.6u m=1
M17 N_20 N_8 N_40 GND mn5  l=0.5u w=0.6u m=1
M18 N_41 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M19 N_18 N_20 GND GND mn5  l=0.5u w=0.6u m=1
M20 N_18 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M21 Q N_15 GND GND mn5  l=0.5u w=0.72u m=1
M22 N_4 N_8 N_3 VDD mp5  l=0.42u w=0.62u m=1
M23 N_24 N_7 N_3 VDD mp5  l=0.42u w=0.6u m=1
M24 VDD N_2 N_24 VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_3 N_23 VDD mp5  l=0.42u w=0.62u m=1
M26 N_2 N_14 N_23 VDD mp5  l=0.42u w=0.62u m=1
M27 N_8 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_7 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_11 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_26 D VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_4 SE N_26 VDD mp5  l=0.42u w=0.62u m=1
M32 N_4 N_11 N_25 VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 SI VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_14 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M35 N_15 N_18 VDD VDD mp5  l=0.42u w=0.62u m=1
M36 Q N_15 VDD VDD mp5  l=0.42u w=0.96u m=1
M37 N_28 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M38 N_28 N_7 N_20 VDD mp5  l=0.42u w=0.62u m=1
M39 N_29 N_8 N_20 VDD mp5  l=0.42u w=0.6u m=1
M40 N_29 N_18 VDD VDD mp5  l=0.42u w=0.6u m=1
M41 VDD N_20 N_27 VDD mp5  l=0.42u w=0.62u m=1
M42 N_18 N_14 N_27 VDD mp5  l=0.42u w=0.62u m=1
.ends sdcfq1
* SPICE INPUT		Mon Sep 24 12:48:34 2018	sdcfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfq2
.subckt sdcfq2 VDD Q GND RN SI SE D CKN
M1 N_14 RN GND GND mn5  l=0.5u w=0.6u m=1
M2 N_15 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_11 SE GND GND mn5  l=0.5u w=0.6u m=1
M4 N_38 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_31 N_11 N_38 GND mn5  l=0.5u w=0.6u m=1
M6 N_31 SI N_37 GND mn5  l=0.5u w=0.6u m=1
M7 N_37 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_8 CKN GND GND mn5  l=0.5u w=0.6u m=1
M9 GND N_8 N_7 GND mn5  l=0.5u w=0.6u m=1
M10 N_3 N_7 N_31 GND mn5  l=0.5u w=0.6u m=1
M11 N_39 N_8 N_3 GND mn5  l=0.5u w=0.6u m=1
M12 N_39 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_2 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_40 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_41 N_7 N_20 GND mn5  l=0.5u w=0.6u m=1
M17 N_20 N_8 N_40 GND mn5  l=0.5u w=0.6u m=1
M18 N_41 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M19 N_18 N_20 GND GND mn5  l=0.5u w=0.6u m=1
M20 N_18 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M21 Q N_15 GND GND mn5  l=0.5u w=0.98u m=1
M22 N_4 N_8 N_3 VDD mp5  l=0.42u w=0.62u m=1
M23 N_24 N_7 N_3 VDD mp5  l=0.42u w=0.6u m=1
M24 VDD N_2 N_24 VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_3 N_23 VDD mp5  l=0.42u w=0.62u m=1
M26 N_2 N_14 N_23 VDD mp5  l=0.42u w=0.62u m=1
M27 N_8 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_7 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_11 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_26 D VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_4 SE N_26 VDD mp5  l=0.42u w=0.62u m=1
M32 N_4 N_11 N_25 VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 SI VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_14 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M35 N_15 N_18 VDD VDD mp5  l=0.42u w=0.62u m=1
M36 Q N_15 VDD VDD mp5  l=0.42u w=1.28u m=1
M37 N_28 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M38 N_28 N_7 N_20 VDD mp5  l=0.42u w=0.62u m=1
M39 N_29 N_8 N_20 VDD mp5  l=0.42u w=0.6u m=1
M40 N_29 N_18 VDD VDD mp5  l=0.42u w=0.6u m=1
M41 VDD N_20 N_27 VDD mp5  l=0.42u w=0.62u m=1
M42 N_18 N_14 N_27 VDD mp5  l=0.42u w=0.62u m=1
.ends sdcfq2
* SPICE INPUT		Mon Sep 24 12:48:43 2018	sdcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb1
.subckt sdcrb1 VDD Q QN GND RN SI SE D CK
M1 N_3 N_7 N_32 GND mn5  l=0.5u w=0.6u m=1
M2 N_61 N_8 N_3 GND mn5  l=0.5u w=0.6u m=1
M3 N_61 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_19 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_62 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_63 N_7 N_15 GND mn5  l=0.5u w=0.6u m=1
M8 GND N_13 N_63 GND mn5  l=0.5u w=0.6u m=1
M9 GND N_15 N_13 GND mn5  l=0.5u w=0.6u m=1
M10 GND N_19 N_13 GND mn5  l=0.5u w=0.6u m=1
M11 N_15 N_8 N_62 GND mn5  l=0.5u w=0.6u m=1
M12 N_11 SE GND GND mn5  l=0.5u w=0.6u m=1
M13 N_65 D GND GND mn5  l=0.5u w=0.6u m=1
M14 N_32 N_11 N_65 GND mn5  l=0.5u w=0.6u m=1
M15 N_32 SI N_64 GND mn5  l=0.5u w=0.6u m=1
M16 N_64 SE GND GND mn5  l=0.5u w=0.6u m=1
M17 N_8 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M18 GND CK N_7 GND mn5  l=0.5u w=0.6u m=1
M19 N_19 RN GND GND mn5  l=0.5u w=0.6u m=1
M20 GND N_13 N_18 GND mn5  l=0.5u w=0.6u m=1
M21 QN N_13 GND GND mn5  l=0.5u w=0.72u m=1
M22 Q N_18 GND GND mn5  l=0.5u w=0.72u m=1
M23 N_4 N_8 N_3 VDD mp5  l=0.42u w=0.62u m=1
M24 N_25 N_7 N_3 VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_2 N_25 VDD mp5  l=0.42u w=0.6u m=1
M26 VDD N_3 N_24 VDD mp5  l=0.42u w=0.62u m=1
M27 N_2 N_19 N_24 VDD mp5  l=0.42u w=0.62u m=1
M28 N_8 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_7 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_11 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_27 D VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_4 SE N_27 VDD mp5  l=0.42u w=0.62u m=1
M33 N_4 N_11 N_26 VDD mp5  l=0.42u w=0.62u m=1
M34 N_26 SI VDD VDD mp5  l=0.42u w=0.62u m=1
M35 N_29 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_29 N_7 N_15 VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_13 N_30 VDD mp5  l=0.42u w=0.6u m=1
M38 VDD N_15 N_28 VDD mp5  l=0.42u w=0.62u m=1
M39 N_13 N_19 N_28 VDD mp5  l=0.42u w=0.62u m=1
M40 N_30 N_8 N_15 VDD mp5  l=0.42u w=0.6u m=1
M41 N_19 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M42 N_18 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M43 QN N_13 VDD VDD mp5  l=0.42u w=0.96u m=1
M44 Q N_18 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdcrb1
* SPICE INPUT		Mon Sep 24 12:48:52 2018	sdcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb2
.subckt sdcrb2 VDD Q QN GND RN SI SE D CK
M1 N_3 N_7 N_32 GND mn5  l=0.5u w=0.6u m=1
M2 N_61 N_8 N_3 GND mn5  l=0.5u w=0.6u m=1
M3 N_61 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_19 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_62 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_63 N_7 N_15 GND mn5  l=0.5u w=0.6u m=1
M8 GND N_13 N_63 GND mn5  l=0.5u w=0.6u m=1
M9 GND N_15 N_13 GND mn5  l=0.5u w=0.6u m=1
M10 GND N_19 N_13 GND mn5  l=0.5u w=0.6u m=1
M11 N_15 N_8 N_62 GND mn5  l=0.5u w=0.6u m=1
M12 N_11 SE GND GND mn5  l=0.5u w=0.6u m=1
M13 N_65 D GND GND mn5  l=0.5u w=0.6u m=1
M14 N_32 N_11 N_65 GND mn5  l=0.5u w=0.6u m=1
M15 N_32 SI N_64 GND mn5  l=0.5u w=0.6u m=1
M16 N_64 SE GND GND mn5  l=0.5u w=0.6u m=1
M17 N_8 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M18 GND CK N_7 GND mn5  l=0.5u w=0.6u m=1
M19 N_19 RN GND GND mn5  l=0.5u w=0.6u m=1
M20 GND N_13 N_18 GND mn5  l=0.5u w=0.6u m=1
M21 QN N_13 GND GND mn5  l=0.5u w=0.98u m=1
M22 Q N_18 GND GND mn5  l=0.5u w=0.98u m=1
M23 N_4 N_8 N_3 VDD mp5  l=0.42u w=0.62u m=1
M24 N_25 N_7 N_3 VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_2 N_25 VDD mp5  l=0.42u w=0.6u m=1
M26 VDD N_3 N_24 VDD mp5  l=0.42u w=0.62u m=1
M27 N_2 N_19 N_24 VDD mp5  l=0.42u w=0.62u m=1
M28 N_8 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_7 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_11 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_27 D VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_4 SE N_27 VDD mp5  l=0.42u w=0.62u m=1
M33 N_4 N_11 N_26 VDD mp5  l=0.42u w=0.62u m=1
M34 N_26 SI VDD VDD mp5  l=0.42u w=0.62u m=1
M35 N_29 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_29 N_7 N_15 VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_13 N_30 VDD mp5  l=0.42u w=0.6u m=1
M38 VDD N_15 N_28 VDD mp5  l=0.42u w=0.62u m=1
M39 N_13 N_19 N_28 VDD mp5  l=0.42u w=0.62u m=1
M40 N_30 N_8 N_15 VDD mp5  l=0.42u w=0.6u m=1
M41 N_19 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M42 N_18 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M43 QN N_13 VDD VDD mp5  l=0.42u w=1.28u m=1
M44 Q N_18 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends sdcrb2
* SPICE INPUT		Mon Sep 24 12:49:00 2018	sdcrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrn1
.subckt sdcrn1 VDD QN GND RN SI SE D CK
M1 N_12 RN GND GND mn5  l=0.5u w=0.6u m=1
M2 QN N_6 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_18 SE GND GND mn5  l=0.5u w=0.6u m=1
M4 N_56 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_28 N_18 N_56 GND mn5  l=0.5u w=0.6u m=1
M6 N_28 SI N_55 GND mn5  l=0.5u w=0.6u m=1
M7 N_55 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M9 GND CK N_14 GND mn5  l=0.5u w=0.6u m=1
M10 N_3 N_14 N_28 GND mn5  l=0.5u w=0.6u m=1
M11 N_57 N_15 N_3 GND mn5  l=0.5u w=0.6u m=1
M12 N_57 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_2 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_8 N_15 N_58 GND mn5  l=0.5u w=0.6u m=1
M16 N_59 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M17 GND N_8 N_6 GND mn5  l=0.5u w=0.6u m=1
M18 N_6 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M19 N_58 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M20 N_59 N_14 N_8 GND mn5  l=0.5u w=0.6u m=1
M21 N_4 N_15 N_3 VDD mp5  l=0.42u w=0.62u m=1
M22 N_22 N_14 N_3 VDD mp5  l=0.42u w=0.6u m=1
M23 VDD N_2 N_22 VDD mp5  l=0.42u w=0.6u m=1
M24 VDD N_3 N_21 VDD mp5  l=0.42u w=0.62u m=1
M25 N_2 N_12 N_21 VDD mp5  l=0.42u w=0.62u m=1
M26 N_25 N_15 N_8 VDD mp5  l=0.42u w=0.6u m=1
M27 VDD N_6 N_25 VDD mp5  l=0.42u w=0.6u m=1
M28 VDD N_8 N_23 VDD mp5  l=0.42u w=0.62u m=1
M29 N_6 N_12 N_23 VDD mp5  l=0.42u w=0.62u m=1
M30 N_24 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 N_14 N_8 VDD mp5  l=0.42u w=0.62u m=1
M32 N_12 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M33 QN N_6 VDD VDD mp5  l=0.42u w=0.96u m=1
M34 N_15 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M35 N_14 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_18 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_27 D VDD VDD mp5  l=0.42u w=0.62u m=1
M38 N_4 SE N_27 VDD mp5  l=0.42u w=0.62u m=1
M39 N_4 N_18 N_26 VDD mp5  l=0.42u w=0.62u m=1
M40 N_26 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdcrn1
* SPICE INPUT		Mon Sep 24 12:49:09 2018	sdcrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrn2
.subckt sdcrn2 VDD QN GND RN SI SE D CK
M1 N_12 RN GND GND mn5  l=0.5u w=0.6u m=1
M2 QN N_6 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_18 SE GND GND mn5  l=0.5u w=0.6u m=1
M4 N_56 D GND GND mn5  l=0.5u w=0.6u m=1
M5 N_28 N_18 N_56 GND mn5  l=0.5u w=0.6u m=1
M6 N_28 SI N_55 GND mn5  l=0.5u w=0.6u m=1
M7 N_55 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M9 GND CK N_14 GND mn5  l=0.5u w=0.6u m=1
M10 N_3 N_14 N_28 GND mn5  l=0.5u w=0.6u m=1
M11 N_57 N_15 N_3 GND mn5  l=0.5u w=0.6u m=1
M12 N_57 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_2 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M14 N_2 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_8 N_15 N_58 GND mn5  l=0.5u w=0.6u m=1
M16 N_59 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M17 GND N_8 N_6 GND mn5  l=0.5u w=0.6u m=1
M18 N_6 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M19 N_58 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M20 N_59 N_14 N_8 GND mn5  l=0.5u w=0.6u m=1
M21 N_4 N_15 N_3 VDD mp5  l=0.42u w=0.62u m=1
M22 N_22 N_14 N_3 VDD mp5  l=0.42u w=0.6u m=1
M23 VDD N_2 N_22 VDD mp5  l=0.42u w=0.6u m=1
M24 VDD N_3 N_21 VDD mp5  l=0.42u w=0.62u m=1
M25 N_2 N_12 N_21 VDD mp5  l=0.42u w=0.62u m=1
M26 N_25 N_15 N_8 VDD mp5  l=0.42u w=0.6u m=1
M27 VDD N_6 N_25 VDD mp5  l=0.42u w=0.6u m=1
M28 VDD N_8 N_23 VDD mp5  l=0.42u w=0.62u m=1
M29 N_6 N_12 N_23 VDD mp5  l=0.42u w=0.62u m=1
M30 N_24 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 N_14 N_8 VDD mp5  l=0.42u w=0.62u m=1
M32 N_12 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M33 QN N_6 VDD VDD mp5  l=0.42u w=1.28u m=1
M34 N_15 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M35 N_14 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_18 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_27 D VDD VDD mp5  l=0.42u w=0.62u m=1
M38 N_4 SE N_27 VDD mp5  l=0.42u w=0.62u m=1
M39 N_4 N_18 N_26 VDD mp5  l=0.42u w=0.62u m=1
M40 N_26 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdcrn2
* SPICE INPUT		Mon Sep 24 12:49:17 2018	sdcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq1
.subckt sdcrq1 VDD Q GND RN SI SE D CK
M1 N_4 N_14 N_30 GND mn5  l=0.5u w=0.6u m=1
M2 N_36 N_15 N_4 GND mn5  l=0.5u w=0.6u m=1
M3 N_36 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_2 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_37 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_12 N_15 N_37 GND mn5  l=0.5u w=0.6u m=1
M8 N_38 N_14 N_12 GND mn5  l=0.5u w=0.6u m=1
M9 N_38 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_10 RN GND GND mn5  l=0.5u w=0.6u m=1
M11 N_18 SE GND GND mn5  l=0.5u w=0.6u m=1
M12 N_40 D GND GND mn5  l=0.5u w=0.6u m=1
M13 N_30 N_18 N_40 GND mn5  l=0.5u w=0.6u m=1
M14 N_30 SI N_39 GND mn5  l=0.5u w=0.6u m=1
M15 N_39 SE GND GND mn5  l=0.5u w=0.6u m=1
M16 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M17 GND CK N_14 GND mn5  l=0.5u w=0.6u m=1
M18 N_7 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M19 GND N_12 Q GND mn5  l=0.5u w=0.72u m=1
M20 N_7 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M21 GND N_10 Q GND mn5  l=0.5u w=0.72u m=1
M22 N_4 N_15 N_3 VDD mp5  l=0.42u w=0.62u m=1
M23 N_22 N_14 N_4 VDD mp5  l=0.42u w=0.6u m=1
M24 VDD N_2 N_22 VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_4 N_21 VDD mp5  l=0.42u w=0.62u m=1
M26 N_2 N_10 N_21 VDD mp5  l=0.42u w=0.62u m=1
M27 N_24 N_10 N_7 VDD mp5  l=0.42u w=0.62u m=1
M28 VDD N_12 N_23 VDD mp5  l=0.42u w=0.96u m=1
M29 VDD N_12 N_24 VDD mp5  l=0.42u w=0.62u m=1
M30 Q N_10 N_23 VDD mp5  l=0.42u w=0.96u m=1
M31 N_25 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_25 N_14 N_12 VDD mp5  l=0.42u w=0.62u m=1
M33 N_26 N_15 N_12 VDD mp5  l=0.42u w=0.6u m=1
M34 N_26 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M35 N_10 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_15 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_14 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M38 N_18 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M39 N_28 D VDD VDD mp5  l=0.42u w=0.62u m=1
M40 N_3 SE N_28 VDD mp5  l=0.42u w=0.62u m=1
M41 N_3 N_18 N_27 VDD mp5  l=0.42u w=0.62u m=1
M42 N_27 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdcrq1
* SPICE INPUT		Mon Sep 24 12:49:26 2018	sdcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq2
.subckt sdcrq2 VDD Q GND RN SI SE D CK
M1 N_4 N_14 N_30 GND mn5  l=0.5u w=0.6u m=1
M2 N_57 N_15 N_4 GND mn5  l=0.5u w=0.6u m=1
M3 N_57 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_2 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_2 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_58 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_12 N_15 N_58 GND mn5  l=0.5u w=0.6u m=1
M8 N_59 N_14 N_12 GND mn5  l=0.5u w=0.6u m=1
M9 N_59 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_10 RN GND GND mn5  l=0.5u w=0.6u m=1
M11 N_18 SE GND GND mn5  l=0.5u w=0.6u m=1
M12 N_61 D GND GND mn5  l=0.5u w=0.6u m=1
M13 N_30 N_18 N_61 GND mn5  l=0.5u w=0.6u m=1
M14 N_30 SI N_60 GND mn5  l=0.5u w=0.6u m=1
M15 N_60 SE GND GND mn5  l=0.5u w=0.6u m=1
M16 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M17 GND CK N_14 GND mn5  l=0.5u w=0.6u m=1
M18 N_7 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M19 GND N_12 Q GND mn5  l=0.5u w=0.98u m=1
M20 N_7 N_12 GND GND mn5  l=0.5u w=0.6u m=1
M21 GND N_10 Q GND mn5  l=0.5u w=0.98u m=1
M22 N_4 N_15 N_3 VDD mp5  l=0.42u w=0.62u m=1
M23 N_22 N_14 N_4 VDD mp5  l=0.42u w=0.6u m=1
M24 VDD N_2 N_22 VDD mp5  l=0.42u w=0.6u m=1
M25 VDD N_4 N_21 VDD mp5  l=0.42u w=0.62u m=1
M26 N_2 N_10 N_21 VDD mp5  l=0.42u w=0.62u m=1
M27 N_24 N_10 N_7 VDD mp5  l=0.42u w=0.62u m=1
M28 VDD N_12 N_23 VDD mp5  l=0.42u w=1.28u m=1
M29 VDD N_12 N_24 VDD mp5  l=0.42u w=0.62u m=1
M30 Q N_10 N_23 VDD mp5  l=0.42u w=1.28u m=1
M31 N_25 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_25 N_14 N_12 VDD mp5  l=0.42u w=0.62u m=1
M33 N_26 N_15 N_12 VDD mp5  l=0.42u w=0.6u m=1
M34 N_26 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M35 N_10 RN VDD VDD mp5  l=0.42u w=0.62u m=1
M36 N_15 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M37 N_14 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M38 N_18 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M39 N_28 D VDD VDD mp5  l=0.42u w=0.62u m=1
M40 N_3 SE N_28 VDD mp5  l=0.42u w=0.62u m=1
M41 N_3 N_18 N_27 VDD mp5  l=0.42u w=0.62u m=1
M42 N_27 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdcrq2
* SPICE INPUT		Mon Sep 24 12:49:33 2018	sdnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb1
.subckt sdnfb1 VDD QN Q GND SI SE D CKN
M1 Q N_5 GND GND mn5  l=0.5u w=0.72u m=1
M2 QN N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_51 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_52 N_14 N_5 GND mn5  l=0.5u w=0.6u m=1
M5 N_51 N_15 N_5 GND mn5  l=0.5u w=0.6u m=1
M6 N_52 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_3 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_11 N_14 N_26 GND mn5  l=0.5u w=0.6u m=1
M9 N_53 N_15 N_11 GND mn5  l=0.5u w=0.6u m=1
M10 N_53 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_10 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_15 CKN GND GND mn5  l=0.5u w=0.6u m=1
M13 GND N_15 N_14 GND mn5  l=0.5u w=0.6u m=1
M14 N_18 SE GND GND mn5  l=0.5u w=0.6u m=1
M15 N_55 D GND GND mn5  l=0.5u w=0.6u m=1
M16 N_26 N_18 N_55 GND mn5  l=0.5u w=0.6u m=1
M17 N_26 SI N_54 GND mn5  l=0.5u w=0.6u m=1
M18 N_54 SE GND GND mn5  l=0.5u w=0.6u m=1
M19 N_21 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_21 N_14 N_5 VDD mp5  l=0.42u w=0.62u m=1
M21 N_22 N_15 N_5 VDD mp5  l=0.42u w=0.6u m=1
M22 N_22 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M23 N_3 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M24 Q N_5 VDD VDD mp5  l=0.42u w=0.96u m=1
M25 QN N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M26 N_12 N_15 N_11 VDD mp5  l=0.42u w=0.62u m=1
M27 N_23 N_14 N_11 VDD mp5  l=0.42u w=0.6u m=1
M28 N_23 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M29 N_10 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_15 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_14 N_15 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_18 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_12 SE N_25 VDD mp5  l=0.42u w=0.62u m=1
M35 N_12 N_18 N_24 VDD mp5  l=0.42u w=0.62u m=1
M36 N_24 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdnfb1
* SPICE INPUT		Mon Sep 24 12:49:40 2018	sdnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb2
.subckt sdnfb2 VDD QN Q GND SI SE D CKN
M1 Q N_5 GND GND mn5  l=0.5u w=0.98u m=1
M2 QN N_3 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_51 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_52 N_14 N_5 GND mn5  l=0.5u w=0.6u m=1
M5 N_51 N_15 N_5 GND mn5  l=0.5u w=0.6u m=1
M6 N_52 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_3 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_11 N_14 N_26 GND mn5  l=0.5u w=0.6u m=1
M9 N_53 N_15 N_11 GND mn5  l=0.5u w=0.6u m=1
M10 N_53 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_10 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_15 CKN GND GND mn5  l=0.5u w=0.6u m=1
M13 GND N_15 N_14 GND mn5  l=0.5u w=0.6u m=1
M14 N_18 SE GND GND mn5  l=0.5u w=0.6u m=1
M15 N_55 D GND GND mn5  l=0.5u w=0.6u m=1
M16 N_26 N_18 N_55 GND mn5  l=0.5u w=0.6u m=1
M17 N_26 SI N_54 GND mn5  l=0.5u w=0.6u m=1
M18 N_54 SE GND GND mn5  l=0.5u w=0.6u m=1
M19 N_21 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_21 N_14 N_5 VDD mp5  l=0.42u w=0.62u m=1
M21 N_22 N_15 N_5 VDD mp5  l=0.42u w=0.6u m=1
M22 N_22 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M23 N_3 N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
M24 Q N_5 VDD VDD mp5  l=0.42u w=1.28u m=1
M25 QN N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M26 N_12 N_15 N_11 VDD mp5  l=0.42u w=0.62u m=1
M27 N_23 N_14 N_11 VDD mp5  l=0.42u w=0.6u m=1
M28 N_23 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M29 N_10 N_11 VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_15 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_14 N_15 VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_18 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_12 SE N_25 VDD mp5  l=0.42u w=0.62u m=1
M35 N_12 N_18 N_24 VDD mp5  l=0.42u w=0.62u m=1
M36 N_24 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdnfb2
* SPICE INPUT		Mon Sep 24 12:49:48 2018	sdnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb1
.subckt sdnrb1 VDD QN Q GND SI SE D CK
M1 QN N_7 GND GND mn5  l=0.5u w=0.72u m=1
M2 Q N_9 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_51 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_52 N_14 N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_51 N_15 N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_52 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_53 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_14 N_26 GND mn5  l=0.5u w=0.6u m=1
M11 N_53 N_15 N_4 GND mn5  l=0.5u w=0.6u m=1
M12 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M13 GND CK N_14 GND mn5  l=0.5u w=0.6u m=1
M14 N_18 SE GND GND mn5  l=0.5u w=0.6u m=1
M15 N_55 D GND GND mn5  l=0.5u w=0.6u m=1
M16 N_26 N_18 N_55 GND mn5  l=0.5u w=0.6u m=1
M17 N_26 SI N_54 GND mn5  l=0.5u w=0.6u m=1
M18 N_54 SE GND GND mn5  l=0.5u w=0.6u m=1
M19 N_5 N_15 N_4 VDD mp5  l=0.42u w=0.62u m=1
M20 N_21 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_14 N_4 VDD mp5  l=0.42u w=0.6u m=1
M23 N_22 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_22 N_14 N_9 VDD mp5  l=0.42u w=0.62u m=1
M25 N_23 N_15 N_9 VDD mp5  l=0.42u w=0.6u m=1
M26 N_23 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M27 N_7 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 QN N_7 VDD VDD mp5  l=0.42u w=0.96u m=1
M29 Q N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M30 N_15 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_14 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_18 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_5 SE N_25 VDD mp5  l=0.42u w=0.62u m=1
M35 N_5 N_18 N_24 VDD mp5  l=0.42u w=0.62u m=1
M36 N_24 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdnrb1
* SPICE INPUT		Mon Sep 24 12:49:55 2018	sdnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb2
.subckt sdnrb2 VDD QN Q GND SI SE D CK
M1 QN N_7 GND GND mn5  l=0.5u w=0.98u m=1
M2 Q N_9 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_51 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M4 N_52 N_14 N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_51 N_15 N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_52 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_53 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_4 N_14 N_26 GND mn5  l=0.5u w=0.6u m=1
M11 N_53 N_15 N_4 GND mn5  l=0.5u w=0.6u m=1
M12 N_15 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M13 GND CK N_14 GND mn5  l=0.5u w=0.6u m=1
M14 N_18 SE GND GND mn5  l=0.5u w=0.6u m=1
M15 N_55 D GND GND mn5  l=0.5u w=0.6u m=1
M16 N_26 N_18 N_55 GND mn5  l=0.5u w=0.6u m=1
M17 N_26 SI N_54 GND mn5  l=0.5u w=0.6u m=1
M18 N_54 SE GND GND mn5  l=0.5u w=0.6u m=1
M19 N_5 N_15 N_4 VDD mp5  l=0.42u w=0.62u m=1
M20 N_21 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_14 N_4 VDD mp5  l=0.42u w=0.6u m=1
M23 N_22 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_22 N_14 N_9 VDD mp5  l=0.42u w=0.62u m=1
M25 N_23 N_15 N_9 VDD mp5  l=0.42u w=0.6u m=1
M26 N_23 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M27 N_7 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 QN N_7 VDD VDD mp5  l=0.42u w=1.28u m=1
M29 Q N_9 VDD VDD mp5  l=0.42u w=1.28u m=1
M30 N_15 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_14 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_18 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_25 D VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_5 SE N_25 VDD mp5  l=0.42u w=0.62u m=1
M35 N_5 N_18 N_24 VDD mp5  l=0.42u w=0.62u m=1
M36 N_24 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdnrb2
* SPICE INPUT		Mon Sep 24 12:50:02 2018	sdnrn1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrn1
.subckt sdnrn1 SE SI D CK GND VDD QN
M1 QN N_14 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_27 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_28 N_8 N_13 GND mn5  l=0.5u w=0.6u m=1
M4 N_27 N_11 N_13 GND mn5  l=0.5u w=0.6u m=1
M5 N_28 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_9 N_8 N_25 GND mn5  l=0.5u w=0.6u m=1
M8 N_29 N_11 N_9 GND mn5  l=0.5u w=0.6u m=1
M9 N_29 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_10 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_11 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M12 GND CK N_8 GND mn5  l=0.5u w=0.6u m=1
M13 N_4 SE GND GND mn5  l=0.5u w=0.6u m=1
M14 N_31 D GND GND mn5  l=0.5u w=0.6u m=1
M15 N_25 N_4 N_31 GND mn5  l=0.5u w=0.6u m=1
M16 N_25 SI N_30 GND mn5  l=0.5u w=0.6u m=1
M17 N_30 SE GND GND mn5  l=0.5u w=0.6u m=1
M18 N_26 N_11 N_9 VDD mp5  l=0.42u w=0.62u m=1
M19 N_50 N_8 N_9 VDD mp5  l=0.42u w=0.6u m=1
M20 N_50 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_10 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_51 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_51 N_8 N_13 VDD mp5  l=0.42u w=0.62u m=1
M24 N_52 N_11 N_13 VDD mp5  l=0.42u w=0.6u m=1
M25 N_52 N_14 VDD VDD mp5  l=0.42u w=0.6u m=1
M26 N_14 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M27 QN N_14 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_11 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_8 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_4 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_54 D VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_26 SE N_54 VDD mp5  l=0.42u w=0.62u m=1
M33 N_26 N_4 N_53 VDD mp5  l=0.42u w=0.62u m=1
M34 N_53 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdnrn1
* SPICE INPUT		Mon Sep 24 12:50:09 2018	sdnrn2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrn2
.subckt sdnrn2 SE SI D CK GND VDD QN
M1 QN N_14 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_50 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_51 N_8 N_13 GND mn5  l=0.5u w=0.6u m=1
M4 N_50 N_11 N_13 GND mn5  l=0.5u w=0.6u m=1
M5 N_51 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_9 N_8 N_25 GND mn5  l=0.5u w=0.6u m=1
M8 N_52 N_11 N_9 GND mn5  l=0.5u w=0.6u m=1
M9 N_52 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_10 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_11 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M12 GND CK N_8 GND mn5  l=0.5u w=0.6u m=1
M13 N_4 SE GND GND mn5  l=0.5u w=0.6u m=1
M14 N_54 D GND GND mn5  l=0.5u w=0.6u m=1
M15 N_25 N_4 N_54 GND mn5  l=0.5u w=0.6u m=1
M16 N_25 SI N_53 GND mn5  l=0.5u w=0.6u m=1
M17 N_53 SE GND GND mn5  l=0.5u w=0.6u m=1
M18 N_26 N_11 N_9 VDD mp5  l=0.42u w=0.62u m=1
M19 N_27 N_8 N_9 VDD mp5  l=0.42u w=0.6u m=1
M20 N_27 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_10 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_28 N_10 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_28 N_8 N_13 VDD mp5  l=0.42u w=0.62u m=1
M24 N_29 N_11 N_13 VDD mp5  l=0.42u w=0.6u m=1
M25 N_29 N_14 VDD VDD mp5  l=0.42u w=0.6u m=1
M26 N_14 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M27 QN N_14 VDD VDD mp5  l=0.42u w=1.28u m=1
M28 N_11 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_8 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_4 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_31 D VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_26 SE N_31 VDD mp5  l=0.42u w=0.62u m=1
M33 N_26 N_4 N_30 VDD mp5  l=0.42u w=0.62u m=1
M34 N_30 SI VDD VDD mp5  l=0.42u w=0.62u m=1
.ends sdnrn2
* SPICE INPUT		Mon Sep 24 12:50:16 2018	sdnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq1
.subckt sdnrq1 VDD Q GND SI SE D CK
M1 Q N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_49 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_50 N_13 N_9 GND mn5  l=0.5u w=0.6u m=1
M4 N_49 N_14 N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_50 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_4 N_13 N_25 GND mn5  l=0.5u w=0.6u m=1
M8 N_51 N_14 N_4 GND mn5  l=0.5u w=0.6u m=1
M9 N_51 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_14 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M12 GND CK N_13 GND mn5  l=0.5u w=0.6u m=1
M13 N_17 SE GND GND mn5  l=0.5u w=0.6u m=1
M14 N_53 D GND GND mn5  l=0.5u w=0.6u m=1
M15 N_25 SI N_52 GND mn5  l=0.5u w=0.6u m=1
M16 N_52 SE GND GND mn5  l=0.5u w=0.6u m=1
M17 N_25 N_17 N_53 GND mn5  l=0.5u w=0.6u m=1
M18 N_5 N_14 N_4 VDD mp5  l=0.42u w=0.62u m=1
M19 N_20 N_13 N_4 VDD mp5  l=0.42u w=0.6u m=1
M20 N_20 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_21 N_13 N_9 VDD mp5  l=0.42u w=0.62u m=1
M24 N_22 N_14 N_9 VDD mp5  l=0.42u w=0.6u m=1
M25 N_22 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M26 N_7 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M27 Q N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M28 N_14 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_13 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_17 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 D VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_5 SE N_24 VDD mp5  l=0.42u w=0.62u m=1
M33 N_23 SI VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_5 N_17 N_23 VDD mp5  l=0.42u w=0.62u m=1
.ends sdnrq1
* SPICE INPUT		Mon Sep 24 12:50:24 2018	sdnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq2
.subckt sdnrq2 VDD Q GND SI SE D CK
M1 Q N_9 GND GND mn5  l=0.5u w=0.98u m=1
M2 N_49 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_50 N_13 N_9 GND mn5  l=0.5u w=0.6u m=1
M4 N_49 N_14 N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_50 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_7 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_4 N_13 N_25 GND mn5  l=0.5u w=0.6u m=1
M8 N_51 N_14 N_4 GND mn5  l=0.5u w=0.6u m=1
M9 N_51 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M10 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M11 N_14 N_13 GND GND mn5  l=0.5u w=0.6u m=1
M12 GND CK N_13 GND mn5  l=0.5u w=0.6u m=1
M13 N_17 SE GND GND mn5  l=0.5u w=0.6u m=1
M14 N_53 D GND GND mn5  l=0.5u w=0.6u m=1
M15 N_25 SI N_52 GND mn5  l=0.5u w=0.6u m=1
M16 N_52 SE GND GND mn5  l=0.5u w=0.6u m=1
M17 N_25 N_17 N_53 GND mn5  l=0.5u w=0.6u m=1
M18 N_5 N_14 N_4 VDD mp5  l=0.42u w=0.62u m=1
M19 N_20 N_13 N_4 VDD mp5  l=0.42u w=0.6u m=1
M20 N_20 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_21 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_21 N_13 N_9 VDD mp5  l=0.42u w=0.62u m=1
M24 N_22 N_14 N_9 VDD mp5  l=0.42u w=0.6u m=1
M25 N_22 N_7 VDD VDD mp5  l=0.42u w=0.6u m=1
M26 N_7 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M27 Q N_9 VDD VDD mp5  l=0.42u w=1.28u m=1
M28 N_14 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M29 N_13 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M30 N_17 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M31 N_24 D VDD VDD mp5  l=0.42u w=0.62u m=1
M32 N_5 SE N_24 VDD mp5  l=0.42u w=0.62u m=1
M33 N_23 SI VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_5 N_17 N_23 VDD mp5  l=0.42u w=0.62u m=1
.ends sdnrq2
* SPICE INPUT		Mon Sep 24 12:50:31 2018	sdpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb1
.subckt sdpfb1 VDD Q QN GND SN CKN SI D SE
M1 N_10 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M2 GND N_12 N_55 GND mn5  l=0.5u w=0.6u m=1
M3 N_14 SN N_55 GND mn5  l=0.5u w=0.6u m=1
M4 N_56 N_4 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_12 N_3 N_33 GND mn5  l=0.5u w=0.6u m=1
M6 N_56 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_33 SI N_57 GND mn5  l=0.5u w=0.6u m=1
M9 N_57 SE GND GND mn5  l=0.5u w=0.6u m=1
M10 N_33 N_7 N_58 GND mn5  l=0.5u w=0.6u m=1
M11 N_58 D GND GND mn5  l=0.5u w=0.6u m=1
M12 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_4 CKN GND GND mn5  l=0.5u w=0.6u m=1
M14 GND SN N_59 GND mn5  l=0.5u w=0.6u m=1
M15 N_60 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_16 N_4 N_60 GND mn5  l=0.5u w=0.6u m=1
M17 N_61 N_3 N_16 GND mn5  l=0.5u w=0.6u m=1
M18 N_18 N_16 N_59 GND mn5  l=0.5u w=0.6u m=1
M19 N_61 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M20 QN N_18 GND GND mn5  l=0.5u w=0.72u m=1
M21 Q N_10 GND GND mn5  l=0.5u w=0.72u m=1
M22 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_4 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_7 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_23 SI VDD VDD mp5  l=0.42u w=0.6u m=1
M26 N_8 N_7 N_23 VDD mp5  l=0.42u w=0.6u m=1
M27 N_24 D VDD VDD mp5  l=0.42u w=0.6u m=1
M28 N_8 SE N_24 VDD mp5  l=0.42u w=0.6u m=1
M29 N_14 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M30 N_18 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M31 N_26 N_3 N_16 VDD mp5  l=0.42u w=0.62u m=1
M32 N_26 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_27 N_4 N_16 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD SN N_14 VDD mp5  l=0.42u w=0.6u m=1
M35 N_18 N_16 VDD VDD mp5  l=0.42u w=0.6u m=1
M36 N_10 N_18 VDD VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_18 N_27 VDD mp5  l=0.42u w=0.6u m=1
M38 N_12 N_4 N_8 VDD mp5  l=0.42u w=0.6u m=1
M39 N_25 N_3 N_12 VDD mp5  l=0.42u w=0.6u m=1
M40 N_25 N_14 VDD VDD mp5  l=0.42u w=0.6u m=1
M41 QN N_18 VDD VDD mp5  l=0.42u w=0.96u m=1
M42 Q N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdpfb1
* SPICE INPUT		Mon Sep 24 12:50:38 2018	sdpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb2
.subckt sdpfb2 VDD Q QN GND SN CKN SI D SE
M1 N_10 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M2 GND N_12 N_55 GND mn5  l=0.5u w=0.6u m=1
M3 N_14 SN N_55 GND mn5  l=0.5u w=0.6u m=1
M4 N_56 N_4 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_12 N_3 N_33 GND mn5  l=0.5u w=0.6u m=1
M6 N_56 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_33 SI N_57 GND mn5  l=0.5u w=0.6u m=1
M9 N_57 SE GND GND mn5  l=0.5u w=0.6u m=1
M10 N_33 N_7 N_58 GND mn5  l=0.5u w=0.6u m=1
M11 N_58 D GND GND mn5  l=0.5u w=0.6u m=1
M12 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_4 CKN GND GND mn5  l=0.5u w=0.6u m=1
M14 GND SN N_59 GND mn5  l=0.5u w=0.6u m=1
M15 N_60 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_16 N_4 N_60 GND mn5  l=0.5u w=0.6u m=1
M17 N_61 N_3 N_16 GND mn5  l=0.5u w=0.6u m=1
M18 N_18 N_16 N_59 GND mn5  l=0.5u w=0.6u m=1
M19 N_61 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M20 QN N_18 GND GND mn5  l=0.5u w=0.98u m=1
M21 Q N_10 GND GND mn5  l=0.5u w=0.98u m=1
M22 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_4 CKN VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_7 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_23 SI VDD VDD mp5  l=0.42u w=0.6u m=1
M26 N_8 N_7 N_23 VDD mp5  l=0.42u w=0.6u m=1
M27 N_24 D VDD VDD mp5  l=0.42u w=0.6u m=1
M28 N_8 SE N_24 VDD mp5  l=0.42u w=0.6u m=1
M29 N_14 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M30 N_18 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M31 N_26 N_3 N_16 VDD mp5  l=0.42u w=0.62u m=1
M32 N_26 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_27 N_4 N_16 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD SN N_14 VDD mp5  l=0.42u w=0.6u m=1
M35 N_18 N_16 VDD VDD mp5  l=0.42u w=0.6u m=1
M36 N_10 N_18 VDD VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_18 N_27 VDD mp5  l=0.42u w=0.6u m=1
M38 N_12 N_4 N_8 VDD mp5  l=0.42u w=0.6u m=1
M39 N_25 N_3 N_12 VDD mp5  l=0.42u w=0.6u m=1
M40 N_25 N_14 VDD VDD mp5  l=0.42u w=0.6u m=1
M41 QN N_18 VDD VDD mp5  l=0.42u w=1.28u m=1
M42 Q N_10 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends sdpfb2
* SPICE INPUT		Mon Sep 24 12:50:46 2018	sdprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb1
.subckt sdprb1 VDD Q QN GND SN CK SI D SE
M1 N_10 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M2 GND N_12 N_55 GND mn5  l=0.5u w=0.6u m=1
M3 N_14 SN N_55 GND mn5  l=0.5u w=0.6u m=1
M4 N_56 N_3 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_12 N_4 N_33 GND mn5  l=0.5u w=0.6u m=1
M6 N_56 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_33 SI N_57 GND mn5  l=0.5u w=0.6u m=1
M9 N_57 SE GND GND mn5  l=0.5u w=0.6u m=1
M10 N_33 N_7 N_58 GND mn5  l=0.5u w=0.6u m=1
M11 N_58 D GND GND mn5  l=0.5u w=0.6u m=1
M12 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.6u m=1
M14 GND SN N_59 GND mn5  l=0.5u w=0.6u m=1
M15 N_60 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_16 N_3 N_60 GND mn5  l=0.5u w=0.6u m=1
M17 N_61 N_4 N_16 GND mn5  l=0.5u w=0.6u m=1
M18 N_18 N_16 N_59 GND mn5  l=0.5u w=0.6u m=1
M19 N_61 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M20 QN N_18 GND GND mn5  l=0.5u w=0.72u m=1
M21 Q N_10 GND GND mn5  l=0.5u w=0.72u m=1
M22 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_4 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_7 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_23 SI VDD VDD mp5  l=0.42u w=0.6u m=1
M26 N_8 N_7 N_23 VDD mp5  l=0.42u w=0.6u m=1
M27 N_24 D VDD VDD mp5  l=0.42u w=0.6u m=1
M28 N_8 SE N_24 VDD mp5  l=0.42u w=0.6u m=1
M29 N_14 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M30 N_18 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M31 N_26 N_4 N_16 VDD mp5  l=0.42u w=0.62u m=1
M32 N_26 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_27 N_3 N_16 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD SN N_14 VDD mp5  l=0.42u w=0.6u m=1
M35 N_18 N_16 VDD VDD mp5  l=0.42u w=0.6u m=1
M36 N_10 N_18 VDD VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_18 N_27 VDD mp5  l=0.42u w=0.6u m=1
M38 N_12 N_3 N_8 VDD mp5  l=0.42u w=0.6u m=1
M39 N_25 N_4 N_12 VDD mp5  l=0.42u w=0.6u m=1
M40 N_25 N_14 VDD VDD mp5  l=0.42u w=0.6u m=1
M41 QN N_18 VDD VDD mp5  l=0.42u w=0.96u m=1
M42 Q N_10 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends sdprb1
* SPICE INPUT		Mon Sep 24 12:50:53 2018	sdprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb2
.subckt sdprb2 VDD Q QN GND SN CK SI D SE
M1 N_10 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M2 GND N_12 N_55 GND mn5  l=0.5u w=0.6u m=1
M3 N_14 SN N_55 GND mn5  l=0.5u w=0.6u m=1
M4 N_56 N_3 N_12 GND mn5  l=0.5u w=0.6u m=1
M5 N_12 N_4 N_33 GND mn5  l=0.5u w=0.6u m=1
M6 N_56 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 SE GND GND mn5  l=0.5u w=0.6u m=1
M8 N_33 SI N_57 GND mn5  l=0.5u w=0.6u m=1
M9 N_57 SE GND GND mn5  l=0.5u w=0.6u m=1
M10 N_33 N_7 N_58 GND mn5  l=0.5u w=0.6u m=1
M11 N_58 D GND GND mn5  l=0.5u w=0.6u m=1
M12 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_4 CK GND GND mn5  l=0.5u w=0.6u m=1
M14 GND SN N_59 GND mn5  l=0.5u w=0.6u m=1
M15 N_60 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_16 N_3 N_60 GND mn5  l=0.5u w=0.6u m=1
M17 N_61 N_4 N_16 GND mn5  l=0.5u w=0.6u m=1
M18 N_18 N_16 N_59 GND mn5  l=0.5u w=0.6u m=1
M19 N_61 N_18 GND GND mn5  l=0.5u w=0.6u m=1
M20 QN N_18 GND GND mn5  l=0.5u w=0.98u m=1
M21 Q N_10 GND GND mn5  l=0.5u w=0.98u m=1
M22 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_4 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_7 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M25 N_23 SI VDD VDD mp5  l=0.42u w=0.6u m=1
M26 N_8 N_7 N_23 VDD mp5  l=0.42u w=0.6u m=1
M27 N_24 D VDD VDD mp5  l=0.42u w=0.6u m=1
M28 N_8 SE N_24 VDD mp5  l=0.42u w=0.6u m=1
M29 N_14 N_12 VDD VDD mp5  l=0.42u w=0.6u m=1
M30 N_18 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M31 N_26 N_4 N_16 VDD mp5  l=0.42u w=0.62u m=1
M32 N_26 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M33 N_27 N_3 N_16 VDD mp5  l=0.42u w=0.6u m=1
M34 VDD SN N_14 VDD mp5  l=0.42u w=0.6u m=1
M35 N_18 N_16 VDD VDD mp5  l=0.42u w=0.6u m=1
M36 N_10 N_18 VDD VDD mp5  l=0.42u w=0.62u m=1
M37 VDD N_18 N_27 VDD mp5  l=0.42u w=0.6u m=1
M38 N_12 N_3 N_8 VDD mp5  l=0.42u w=0.6u m=1
M39 N_25 N_4 N_12 VDD mp5  l=0.42u w=0.6u m=1
M40 N_25 N_14 VDD VDD mp5  l=0.42u w=0.6u m=1
M41 QN N_18 VDD VDD mp5  l=0.42u w=1.28u m=1
M42 Q N_10 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends sdprb2
* SPICE INPUT		Mon Sep 24 12:51:01 2018	sdprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq1
.subckt sdprq1 GND Q VDD SN SE SI D CK
M1 Q N_17 N_20 GND mn5  l=0.5u w=0.72u m=1
M2 GND SN N_20 GND mn5  l=0.5u w=0.72u m=1
M3 N_6 N_14 N_5 GND mn5  l=0.5u w=0.6u m=1
M4 N_22 N_13 N_6 GND mn5  l=0.5u w=0.6u m=1
M5 N_22 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M6 GND N_6 N_21 GND mn5  l=0.5u w=0.6u m=1
M7 N_4 SN N_21 GND mn5  l=0.5u w=0.6u m=1
M8 N_10 SE GND GND mn5  l=0.5u w=0.6u m=1
M9 N_24 D GND GND mn5  l=0.5u w=0.6u m=1
M10 N_5 N_10 N_24 GND mn5  l=0.5u w=0.6u m=1
M11 N_5 SI N_23 GND mn5  l=0.5u w=0.6u m=1
M12 N_23 SE GND GND mn5  l=0.5u w=0.6u m=1
M13 N_14 CK GND GND mn5  l=0.5u w=0.6u m=1
M14 N_13 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_26 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_17 N_13 N_26 GND mn5  l=0.5u w=0.6u m=1
M17 N_27 N_14 N_17 GND mn5  l=0.5u w=0.6u m=1
M18 N_27 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M19 GND SN N_25 GND mn5  l=0.5u w=0.6u m=1
M20 N_15 N_17 N_25 GND mn5  l=0.5u w=0.6u m=1
M21 N_14 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_13 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_10 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_54 D VDD VDD mp5  l=0.42u w=0.6u m=1
M25 N_29 SE N_54 VDD mp5  l=0.42u w=0.6u m=1
M26 N_29 N_10 N_53 VDD mp5  l=0.42u w=0.6u m=1
M27 N_53 SI VDD VDD mp5  l=0.42u w=0.6u m=1
M28 N_6 N_13 N_29 VDD mp5  l=0.42u w=0.6u m=1
M29 N_55 N_14 N_6 VDD mp5  l=0.42u w=0.6u m=1
M30 N_55 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M31 N_4 N_6 VDD VDD mp5  l=0.42u w=0.6u m=1
M32 VDD SN N_4 VDD mp5  l=0.42u w=0.6u m=1
M33 N_56 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_17 N_14 N_56 VDD mp5  l=0.42u w=0.62u m=1
M35 N_57 N_13 N_17 VDD mp5  l=0.42u w=0.6u m=1
M36 VDD N_15 N_57 VDD mp5  l=0.42u w=0.6u m=1
M37 N_15 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M38 VDD N_17 Q VDD mp5  l=0.42u w=0.96u m=1
M39 VDD N_17 N_15 VDD mp5  l=0.42u w=0.6u m=1
M40 VDD SN Q VDD mp5  l=0.42u w=0.96u m=1
.ends sdprq1
* SPICE INPUT		Mon Sep 24 12:51:08 2018	sdprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq2
.subckt sdprq2 GND Q VDD SN SE SI D CK
M1 Q N_17 N_20 GND mn5  l=0.5u w=0.98u m=1
M2 GND SN N_20 GND mn5  l=0.5u w=0.98u m=1
M3 N_6 N_14 N_5 GND mn5  l=0.5u w=0.6u m=1
M4 N_22 N_13 N_6 GND mn5  l=0.5u w=0.6u m=1
M5 N_22 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M6 GND N_6 N_21 GND mn5  l=0.5u w=0.6u m=1
M7 N_4 SN N_21 GND mn5  l=0.5u w=0.6u m=1
M8 N_10 SE GND GND mn5  l=0.5u w=0.6u m=1
M9 N_24 D GND GND mn5  l=0.5u w=0.6u m=1
M10 N_5 N_10 N_24 GND mn5  l=0.5u w=0.6u m=1
M11 N_5 SI N_23 GND mn5  l=0.5u w=0.6u m=1
M12 N_23 SE GND GND mn5  l=0.5u w=0.6u m=1
M13 N_14 CK GND GND mn5  l=0.5u w=0.6u m=1
M14 N_13 N_14 GND GND mn5  l=0.5u w=0.6u m=1
M15 N_26 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M16 N_17 N_13 N_26 GND mn5  l=0.5u w=0.6u m=1
M17 N_27 N_14 N_17 GND mn5  l=0.5u w=0.6u m=1
M18 N_27 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M19 GND SN N_25 GND mn5  l=0.5u w=0.6u m=1
M20 N_15 N_17 N_25 GND mn5  l=0.5u w=0.6u m=1
M21 N_14 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_13 N_14 VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_10 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_54 D VDD VDD mp5  l=0.42u w=0.6u m=1
M25 N_29 SE N_54 VDD mp5  l=0.42u w=0.6u m=1
M26 N_29 N_10 N_53 VDD mp5  l=0.42u w=0.6u m=1
M27 N_53 SI VDD VDD mp5  l=0.42u w=0.6u m=1
M28 N_6 N_13 N_29 VDD mp5  l=0.42u w=0.6u m=1
M29 N_55 N_14 N_6 VDD mp5  l=0.42u w=0.6u m=1
M30 N_55 N_4 VDD VDD mp5  l=0.42u w=0.6u m=1
M31 N_4 N_6 VDD VDD mp5  l=0.42u w=0.6u m=1
M32 VDD SN N_4 VDD mp5  l=0.42u w=0.6u m=1
M33 N_56 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M34 N_17 N_14 N_56 VDD mp5  l=0.42u w=0.62u m=1
M35 N_57 N_13 N_17 VDD mp5  l=0.42u w=0.6u m=1
M36 VDD N_15 N_57 VDD mp5  l=0.42u w=0.6u m=1
M37 N_15 SN VDD VDD mp5  l=0.42u w=0.6u m=1
M38 VDD N_17 Q VDD mp5  l=0.42u w=1.28u m=1
M39 VDD N_17 N_15 VDD mp5  l=0.42u w=0.6u m=1
M40 VDD SN Q VDD mp5  l=0.42u w=1.28u m=1
.ends sdprq2
* SPICE INPUT		Mon Sep 24 12:51:15 2018	tiehi
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tiehi
.subckt tiehi VDD Y GND
M1 N_5 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_5 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends tiehi
* SPICE INPUT		Mon Sep 24 12:51:23 2018	tielo
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tielo
.subckt tielo VDD GND Y
M1 Y N_3 GND GND mn5  l=0.5u w=0.6u m=1
M2 N_3 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends tielo
* SPICE INPUT		Mon Sep 24 12:51:30 2018	tlatncad1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad1
.subckt tlatncad1 VDD ECK GND CK E
M1 ECK N_9 GND GND mn5  l=0.5u w=0.72u m=1
M2 ECK N_3 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M4 N_27 N_7 N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_7 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_26 E GND GND mn5  l=0.5u w=0.6u m=1
M7 N_26 N_3 N_9 GND mn5  l=0.5u w=0.6u m=1
M8 N_27 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M9 GND N_9 N_6 GND mn5  l=0.5u w=0.6u m=1
M10 N_11 N_9 ECK VDD mp5  l=0.42u w=0.96u m=1
M11 N_11 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M12 N_3 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_12 N_7 N_9 VDD mp5  l=0.42u w=0.62u m=1
M14 VDD N_3 N_7 VDD mp5  l=0.42u w=0.62u m=1
M15 N_12 E VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_13 N_3 N_9 VDD mp5  l=0.42u w=0.6u m=1
M17 N_13 N_6 VDD VDD mp5  l=0.42u w=0.6u m=1
M18 N_6 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends tlatncad1
* SPICE INPUT		Mon Sep 24 12:51:37 2018	tlatncad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad2
.subckt tlatncad2 VDD ECK GND CK E
M1 ECK N_9 GND GND mn5  l=0.5u w=0.98u m=1
M2 ECK N_3 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M4 N_27 N_7 N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_7 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_26 E GND GND mn5  l=0.5u w=0.6u m=1
M7 N_26 N_3 N_9 GND mn5  l=0.5u w=0.6u m=1
M8 N_27 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M9 GND N_9 N_6 GND mn5  l=0.5u w=0.6u m=1
M10 N_11 N_9 ECK VDD mp5  l=0.42u w=1.28u m=1
M11 N_11 N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
M12 N_3 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_12 N_7 N_9 VDD mp5  l=0.42u w=0.62u m=1
M14 VDD N_3 N_7 VDD mp5  l=0.42u w=0.62u m=1
M15 N_12 E VDD VDD mp5  l=0.42u w=0.62u m=1
M16 N_13 N_3 N_9 VDD mp5  l=0.42u w=0.6u m=1
M17 N_13 N_6 VDD VDD mp5  l=0.42u w=0.6u m=1
M18 N_6 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends tlatncad2
* SPICE INPUT		Mon Sep 24 12:51:45 2018	tlatncad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad4
.subckt tlatncad4 CK E GND VDD ECK
M1 N_2 N_9 N_15 GND mn5  l=0.5u w=0.6u m=1
M2 N_15 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_16 E GND GND mn5  l=0.5u w=0.6u m=1
M4 N_2 N_3 N_16 GND mn5  l=0.5u w=0.6u m=1
M5 N_3 CK GND GND mn5  l=0.5u w=0.6u m=1
M6 N_9 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M7 GND N_3 ECK GND mn5  l=0.5u w=0.735u m=1
M8 GND N_3 ECK GND mn5  l=0.5u w=0.735u m=1
M9 ECK N_2 GND GND mn5  l=0.5u w=0.735u m=1
M10 ECK N_2 GND GND mn5  l=0.5u w=0.735u m=1
M11 N_8 N_2 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_3 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M13 N_9 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M14 N_8 N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_31 N_8 VDD VDD mp5  l=0.42u w=0.6u m=1
M16 N_32 E VDD VDD mp5  l=0.42u w=0.62u m=1
M17 N_32 N_9 N_2 VDD mp5  l=0.42u w=0.62u m=1
M18 N_2 N_3 N_31 VDD mp5  l=0.42u w=0.6u m=1
M19 N_14 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_14 N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
M21 ECK N_2 N_14 VDD mp5  l=0.42u w=0.96u m=1
M22 N_14 N_2 ECK VDD mp5  l=0.42u w=0.96u m=1
.ends tlatncad4
* SPICE INPUT		Mon Sep 24 12:51:52 2018	tlatntscad1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad1
.subckt tlatntscad1 VDD ECK GND CK E SE
M1 ECK N_11 GND GND mn5  l=0.5u w=0.72u m=1
M2 N_11 CK GND GND mn5  l=0.5u w=0.6u m=1
M3 ECK N_6 GND GND mn5  l=0.5u w=0.72u m=1
M4 N_8 N_9 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_9 SE GND GND mn5  l=0.5u w=0.6u m=1
M6 N_9 E GND GND mn5  l=0.5u w=0.6u m=1
M7 N_35 N_11 N_6 GND mn5  l=0.5u w=0.6u m=1
M8 N_36 N_4 N_6 GND mn5  l=0.5u w=0.6u m=1
M9 N_36 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M10 GND N_6 N_3 GND mn5  l=0.5u w=0.6u m=1
M11 N_4 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_35 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M13 N_15 N_11 N_6 VDD mp5  l=0.42u w=0.6u m=1
M14 N_14 N_4 N_6 VDD mp5  l=0.42u w=0.62u m=1
M15 N_15 N_3 VDD VDD mp5  l=0.42u w=0.6u m=1
M16 N_3 N_6 VDD VDD mp5  l=0.42u w=0.62u m=1
M17 VDD N_11 N_4 VDD mp5  l=0.42u w=0.62u m=1
M18 N_14 N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_8 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_16 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_16 E N_9 VDD mp5  l=0.42u w=0.62u m=1
M22 N_17 N_11 VDD VDD mp5  l=0.42u w=0.96u m=1
M23 N_11 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M24 N_17 N_6 ECK VDD mp5  l=0.42u w=0.96u m=1
.ends tlatntscad1
* SPICE INPUT		Mon Sep 24 12:51:59 2018	tlatntscad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad2
.subckt tlatntscad2 VDD ECK GND CK SE E
M1 N_11 CK GND GND mn5  l=0.5u w=0.6u m=1
M2 ECK N_11 GND GND mn5  l=0.5u w=0.98u m=1
M3 ECK N_9 GND GND mn5  l=0.5u w=0.98u m=1
M4 N_4 E GND GND mn5  l=0.5u w=0.6u m=1
M5 N_4 SE GND GND mn5  l=0.5u w=0.6u m=1
M6 N_3 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_7 N_11 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_35 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_35 N_11 N_9 GND mn5  l=0.5u w=0.6u m=1
M10 N_36 N_7 N_9 GND mn5  l=0.5u w=0.6u m=1
M11 N_36 N_6 GND GND mn5  l=0.5u w=0.6u m=1
M12 GND N_9 N_6 GND mn5  l=0.5u w=0.6u m=1
M13 N_14 E N_4 VDD mp5  l=0.42u w=0.62u m=1
M14 N_14 SE VDD VDD mp5  l=0.42u w=0.62u m=1
M15 N_3 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M16 VDD N_11 N_7 VDD mp5  l=0.42u w=0.62u m=1
M17 N_15 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M18 N_16 N_11 N_9 VDD mp5  l=0.42u w=0.6u m=1
M19 N_15 N_7 N_9 VDD mp5  l=0.42u w=0.62u m=1
M20 N_16 N_6 VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_6 N_9 VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_11 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M23 N_17 N_11 VDD VDD mp5  l=0.42u w=1.28u m=1
M24 N_17 N_9 ECK VDD mp5  l=0.42u w=1.28u m=1
.ends tlatntscad2
* SPICE INPUT		Mon Sep 24 12:52:07 2018	tlatntscad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad4
.subckt tlatntscad4 VDD ECK GND CK E SE
M1 N_16 E GND GND mn5  l=0.5u w=0.6u m=1
M2 N_15 N_16 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_16 SE GND GND mn5  l=0.5u w=0.6u m=1
M4 GND N_13 N_10 GND mn5  l=0.5u w=0.6u m=1
M5 N_41 N_10 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_41 N_11 N_13 GND mn5  l=0.5u w=0.6u m=1
M7 N_40 N_8 N_13 GND mn5  l=0.5u w=0.6u m=1
M8 N_40 N_15 GND GND mn5  l=0.5u w=0.6u m=1
M9 N_11 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M10 ECK N_8 GND GND mn5  l=0.5u w=0.735u m=1
M11 ECK N_8 GND GND mn5  l=0.5u w=0.735u m=1
M12 N_8 CK GND GND mn5  l=0.5u w=0.6u m=1
M13 ECK N_13 GND GND mn5  l=0.5u w=0.735u m=1
M14 ECK N_13 GND GND mn5  l=0.5u w=0.735u m=1
M15 N_3 N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M16 N_3 N_8 VDD VDD mp5  l=0.42u w=0.96u m=1
M17 N_3 N_13 ECK VDD mp5  l=0.42u w=0.96u m=1
M18 N_3 N_13 ECK VDD mp5  l=0.42u w=0.96u m=1
M19 N_8 CK VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_10 N_13 VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_19 N_10 VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_18 N_11 N_13 VDD mp5  l=0.42u w=0.62u m=1
M23 N_19 N_8 N_13 VDD mp5  l=0.42u w=0.6u m=1
M24 N_18 N_15 VDD VDD mp5  l=0.42u w=0.62u m=1
M25 VDD N_8 N_11 VDD mp5  l=0.42u w=0.62u m=1
M26 N_20 E N_16 VDD mp5  l=0.42u w=0.62u m=1
M27 N_15 N_16 VDD VDD mp5  l=0.42u w=0.62u m=1
M28 N_20 SE VDD VDD mp5  l=0.42u w=0.62u m=1
.ends tlatntscad4
* SPICE INPUT		Mon Sep 24 12:52:14 2018	xn02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d0
.subckt xn02d0 VDD Y GND A B
M1 N_4 B GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A N_3 GND mn5  l=0.5u w=0.6u m=1
M3 N_8 A N_4 GND mn5  l=0.5u w=0.6u m=1
M4 N_8 N_3 N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_9 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M6 Y N_8 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_3 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_8 N_3 N_4 VDD mp5  l=0.42u w=0.62u m=1
M10 N_9 A N_8 VDD mp5  l=0.42u w=0.62u m=1
M11 N_9 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Y N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends xn02d0
* SPICE INPUT		Mon Sep 24 12:52:21 2018	xn02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d1
.subckt xn02d1 A B GND VDD Y
M1 N_4 B GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A N_5 GND mn5  l=0.5u w=0.6u m=1
M3 N_3 N_5 N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_11 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_3 GND GND mn5  l=0.5u w=0.72u m=1
M6 N_3 A N_4 GND mn5  l=0.5u w=0.6u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_3 N_5 N_4 VDD mp5  l=0.42u w=0.62u m=1
M10 N_11 A N_3 VDD mp5  l=0.42u w=0.62u m=1
M11 N_11 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Y N_3 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends xn02d1
* SPICE INPUT		Mon Sep 24 12:52:28 2018	xn02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d2
.subckt xn02d2 A B GND VDD Y
M1 N_4 B GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A N_5 GND mn5  l=0.5u w=0.6u m=1
M3 N_3 N_5 N_11 GND mn5  l=0.5u w=0.6u m=1
M4 N_11 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M5 Y N_3 GND GND mn5  l=0.5u w=0.98u m=1
M6 N_3 A N_4 GND mn5  l=0.5u w=0.6u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_3 N_5 N_4 VDD mp5  l=0.42u w=0.62u m=1
M10 N_11 A N_3 VDD mp5  l=0.42u w=0.62u m=1
M11 N_11 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Y N_3 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends xn02d2
* SPICE INPUT		Mon Sep 24 12:52:36 2018	xn03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d0
.subckt xn03d0 VDD Y GND C B A
M1 N_6 N_14 N_5 GND mn5  l=0.5u w=0.6u m=1
M2 N_3 N_14 N_2 GND mn5  l=0.5u w=0.6u m=1
M3 N_6 B N_2 GND mn5  l=0.5u w=0.6u m=1
M4 N_5 B N_3 GND mn5  l=0.5u w=0.6u m=1
M5 N_2 C N_7 GND mn5  l=0.5u w=0.6u m=1
M6 N_5 N_12 N_7 GND mn5  l=0.5u w=0.6u m=1
M7 Y N_7 GND GND mn5  l=0.5u w=0.6u m=1
M8 N_12 C GND GND mn5  l=0.5u w=0.6u m=1
M9 N_14 B GND GND mn5  l=0.5u w=0.6u m=1
M10 N_3 A GND GND mn5  l=0.5u w=0.6u m=1
M11 N_6 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_5 N_14 N_3 VDD mp5  l=0.42u w=0.62u m=1
M13 N_6 N_14 N_2 VDD mp5  l=0.42u w=0.62u m=1
M14 N_6 B N_5 VDD mp5  l=0.42u w=0.62u m=1
M15 N_3 B N_2 VDD mp5  l=0.42u w=0.62u m=1
M16 N_5 C N_7 VDD mp5  l=0.42u w=0.62u m=1
M17 N_2 N_12 N_7 VDD mp5  l=0.42u w=0.62u m=1
M18 Y N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
M19 N_12 C VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_14 B VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_3 A VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_6 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends xn03d0
* SPICE INPUT		Mon Sep 24 12:52:43 2018	xn03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d1
.subckt xn03d1 C B A VDD Y GND
M1 N_14 N_6 N_13 GND mn5  l=0.5u w=0.6u m=1
M2 N_7 N_6 N_10 GND mn5  l=0.5u w=0.6u m=1
M3 N_14 B N_10 GND mn5  l=0.5u w=0.6u m=1
M4 N_13 B N_7 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 C N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_13 N_2 N_9 GND mn5  l=0.5u w=0.6u m=1
M7 Y N_9 GND GND mn5  l=0.5u w=0.72u m=1
M8 N_2 C GND GND mn5  l=0.5u w=0.6u m=1
M9 N_6 B GND GND mn5  l=0.5u w=0.6u m=1
M10 N_7 A GND GND mn5  l=0.5u w=0.6u m=1
M11 N_14 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_13 N_6 N_7 VDD mp5  l=0.42u w=0.62u m=1
M13 N_14 N_6 N_10 VDD mp5  l=0.42u w=0.62u m=1
M14 N_14 B N_13 VDD mp5  l=0.42u w=0.62u m=1
M15 N_7 B N_10 VDD mp5  l=0.42u w=0.62u m=1
M16 N_13 C N_9 VDD mp5  l=0.42u w=0.62u m=1
M17 N_10 N_2 N_9 VDD mp5  l=0.42u w=0.62u m=1
M18 Y N_9 VDD VDD mp5  l=0.42u w=0.96u m=1
M19 N_2 C VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_6 B VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_7 A VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_14 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends xn03d1
* SPICE INPUT		Mon Sep 24 12:52:51 2018	xn03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d2
.subckt xn03d2 C B A VDD Y GND
M1 N_14 N_6 N_13 GND mn5  l=0.5u w=0.6u m=1
M2 N_7 N_6 N_10 GND mn5  l=0.5u w=0.6u m=1
M3 N_14 B N_10 GND mn5  l=0.5u w=0.6u m=1
M4 N_13 B N_7 GND mn5  l=0.5u w=0.6u m=1
M5 N_10 C N_9 GND mn5  l=0.5u w=0.6u m=1
M6 N_13 N_2 N_9 GND mn5  l=0.5u w=0.6u m=1
M7 Y N_9 GND GND mn5  l=0.5u w=0.98u m=1
M8 N_2 C GND GND mn5  l=0.5u w=0.6u m=1
M9 N_6 B GND GND mn5  l=0.5u w=0.6u m=1
M10 N_7 A GND GND mn5  l=0.5u w=0.6u m=1
M11 N_14 N_7 GND GND mn5  l=0.5u w=0.6u m=1
M12 N_13 N_6 N_7 VDD mp5  l=0.42u w=0.62u m=1
M13 N_14 N_6 N_10 VDD mp5  l=0.42u w=0.62u m=1
M14 N_14 B N_13 VDD mp5  l=0.42u w=0.62u m=1
M15 N_7 B N_10 VDD mp5  l=0.42u w=0.62u m=1
M16 N_13 C N_9 VDD mp5  l=0.42u w=0.62u m=1
M17 N_10 N_2 N_9 VDD mp5  l=0.42u w=0.62u m=1
M18 Y N_9 VDD VDD mp5  l=0.42u w=1.28u m=1
M19 N_2 C VDD VDD mp5  l=0.42u w=0.62u m=1
M20 N_6 B VDD VDD mp5  l=0.42u w=0.62u m=1
M21 N_7 A VDD VDD mp5  l=0.42u w=0.62u m=1
M22 N_14 N_7 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends xn03d2
* SPICE INPUT		Mon Sep 24 12:52:58 2018	xr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d0
.subckt xr02d0 VDD Y GND A B
M1 N_4 B GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A N_3 GND mn5  l=0.5u w=0.6u m=1
M3 N_8 N_3 N_4 GND mn5  l=0.5u w=0.6u m=1
M4 N_8 A N_9 GND mn5  l=0.5u w=0.6u m=1
M5 N_9 N_4 GND GND mn5  l=0.5u w=0.6u m=1
M6 Y N_8 GND GND mn5  l=0.5u w=0.6u m=1
M7 N_4 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_3 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_8 A N_4 VDD mp5  l=0.42u w=0.62u m=1
M10 N_9 N_3 N_8 VDD mp5  l=0.42u w=0.62u m=1
M11 N_9 N_4 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Y N_8 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends xr02d0
* SPICE INPUT		Mon Sep 24 12:53:05 2018	xr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d1
.subckt xr02d1 A B GND VDD Y
M1 N_3 B GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A N_5 GND mn5  l=0.5u w=0.6u m=1
M3 N_2 N_5 N_3 GND mn5  l=0.5u w=0.6u m=1
M4 N_2 A N_11 GND mn5  l=0.5u w=0.6u m=1
M5 N_11 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M7 N_3 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_2 A N_3 VDD mp5  l=0.42u w=0.62u m=1
M10 N_11 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M11 N_11 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
.ends xr02d1
* SPICE INPUT		Mon Sep 24 12:53:12 2018	xr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d2
.subckt xr02d2 A B GND VDD Y
M1 N_3 B GND GND mn5  l=0.5u w=0.6u m=1
M2 GND A N_5 GND mn5  l=0.5u w=0.6u m=1
M3 N_2 N_5 N_3 GND mn5  l=0.5u w=0.6u m=1
M4 N_2 A N_11 GND mn5  l=0.5u w=0.6u m=1
M5 N_11 N_3 GND GND mn5  l=0.5u w=0.6u m=1
M6 Y N_2 GND GND mn5  l=0.5u w=0.98u m=1
M7 N_3 B VDD VDD mp5  l=0.42u w=0.62u m=1
M8 N_5 A VDD VDD mp5  l=0.42u w=0.62u m=1
M9 N_2 A N_3 VDD mp5  l=0.42u w=0.62u m=1
M10 N_11 N_5 N_2 VDD mp5  l=0.42u w=0.62u m=1
M11 N_11 N_3 VDD VDD mp5  l=0.42u w=0.62u m=1
M12 Y N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
.ends xr02d2
* SPICE INPUT		Mon Sep 24 12:53:19 2018	xr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d0
.subckt xr03d0 A C B VDD Y GND
M1 N_4 C GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_2 GND GND mn5  l=0.5u w=0.6u m=1
M3 N_6 B GND GND mn5  l=0.5u w=0.6u m=1
M4 N_16 N_5 GND GND mn5  l=0.5u w=0.6u m=1
M5 N_5 A GND GND mn5  l=0.5u w=0.6u m=1
M6 N_16 B N_12 GND mn5  l=0.5u w=0.6u m=1
M7 N_11 B N_5 GND mn5  l=0.5u w=0.6u m=1
M8 N_16 N_6 N_11 GND mn5  l=0.5u w=0.6u m=1
M9 N_5 N_6 N_12 GND mn5  l=0.5u w=0.6u m=1
M10 N_11 C N_2 GND mn5  l=0.5u w=0.6u m=1
M11 N_12 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M12 N_12 C N_2 VDD mp5  l=0.42u w=0.6u m=1
M13 N_11 N_4 N_2 VDD mp5  l=0.42u w=0.6u m=1
M14 N_6 B VDD VDD mp5  l=0.42u w=0.6u m=1
M15 N_16 N_5 VDD VDD mp5  l=0.42u w=0.6u m=1
M16 N_5 A VDD VDD mp5  l=0.42u w=0.6u m=1
M17 N_16 B N_11 VDD mp5  l=0.42u w=0.6u m=1
M18 N_5 B N_12 VDD mp5  l=0.42u w=0.6u m=1
M19 N_11 N_6 N_5 VDD mp5  l=0.42u w=0.6u m=1
M20 N_16 N_6 N_12 VDD mp5  l=0.42u w=0.6u m=1
M21 N_4 C VDD VDD mp5  l=0.42u w=0.6u m=1
M22 Y N_2 VDD VDD mp5  l=0.42u w=0.62u m=1
.ends xr03d0
* SPICE INPUT		Mon Sep 24 12:53:26 2018	xr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d1
.subckt xr03d1 C B A VDD Y GND
M1 N_4 C GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_2 GND GND mn5  l=0.5u w=0.72u m=1
M3 N_7 B GND GND mn5  l=0.5u w=0.6u m=1
M4 N_8 A GND GND mn5  l=0.5u w=0.6u m=1
M5 N_14 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_7 N_13 GND mn5  l=0.5u w=0.6u m=1
M7 N_8 N_7 N_10 GND mn5  l=0.5u w=0.6u m=1
M8 N_14 B N_10 GND mn5  l=0.5u w=0.6u m=1
M9 N_13 B N_8 GND mn5  l=0.5u w=0.6u m=1
M10 N_10 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M11 N_13 C N_2 GND mn5  l=0.5u w=0.6u m=1
M12 N_13 N_7 N_8 VDD mp5  l=0.42u w=0.6u m=1
M13 N_14 N_7 N_10 VDD mp5  l=0.42u w=0.6u m=1
M14 N_14 B N_13 VDD mp5  l=0.42u w=0.6u m=1
M15 N_8 B N_10 VDD mp5  l=0.42u w=0.6u m=1
M16 N_13 N_4 N_2 VDD mp5  l=0.42u w=0.6u m=1
M17 N_10 C N_2 VDD mp5  l=0.42u w=0.6u m=1
M18 N_4 C VDD VDD mp5  l=0.42u w=0.6u m=1
M19 Y N_2 VDD VDD mp5  l=0.42u w=0.96u m=1
M20 N_7 B VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_8 A VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_14 N_8 VDD VDD mp5  l=0.42u w=0.6u m=1
.ends xr03d1
* SPICE INPUT		Mon Sep 24 12:53:34 2018	xr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d2
.subckt xr03d2 C B A VDD Y GND
M1 N_4 C GND GND mn5  l=0.5u w=0.6u m=1
M2 Y N_2 GND GND mn5  l=0.5u w=0.98u m=1
M3 N_7 B GND GND mn5  l=0.5u w=0.6u m=1
M4 N_8 A GND GND mn5  l=0.5u w=0.6u m=1
M5 N_14 N_8 GND GND mn5  l=0.5u w=0.6u m=1
M6 N_14 N_7 N_13 GND mn5  l=0.5u w=0.6u m=1
M7 N_8 N_7 N_10 GND mn5  l=0.5u w=0.6u m=1
M8 N_14 B N_10 GND mn5  l=0.5u w=0.6u m=1
M9 N_13 B N_8 GND mn5  l=0.5u w=0.6u m=1
M10 N_10 N_4 N_2 GND mn5  l=0.5u w=0.6u m=1
M11 N_13 C N_2 GND mn5  l=0.5u w=0.6u m=1
M12 N_13 N_7 N_8 VDD mp5  l=0.42u w=0.6u m=1
M13 N_14 N_7 N_10 VDD mp5  l=0.42u w=0.6u m=1
M14 N_14 B N_13 VDD mp5  l=0.42u w=0.6u m=1
M15 N_8 B N_10 VDD mp5  l=0.42u w=0.6u m=1
M16 N_13 N_4 N_2 VDD mp5  l=0.42u w=0.6u m=1
M17 N_10 C N_2 VDD mp5  l=0.42u w=0.6u m=1
M18 N_4 C VDD VDD mp5  l=0.42u w=0.6u m=1
M19 Y N_2 VDD VDD mp5  l=0.42u w=1.28u m=1
M20 N_7 B VDD VDD mp5  l=0.42u w=0.6u m=1
M21 N_8 A VDD VDD mp5  l=0.42u w=0.6u m=1
M22 N_14 N_8 VDD VDD mp5  l=0.42u w=0.6u m=1
.ends xr03d2
