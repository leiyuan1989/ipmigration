* SPICE INPUT		Tue Jul 31 18:28:43 2018	ad01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d0
.subckt ad01d0 VDD CO S GND CI B A
M1 S N_15 GND GND mn15  l=0.13u w=0.26u m=1
M2 CO N_12 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.27u m=1
M4 N_69 N_6 GND GND mn15  l=0.13u w=0.27u m=1
M5 N_69 N_11 N_5 GND mn15  l=0.13u w=0.27u m=1
M6 N_5 B N_6 GND mn15  l=0.13u w=0.27u m=1
M7 N_11 B GND GND mn15  l=0.13u w=0.27u m=1
M8 GND N_5 N_10 GND mn15  l=0.13u w=0.27u m=1
M9 N_13 N_5 N_12 GND mn15  l=0.13u w=0.27u m=1
M10 N_11 N_10 N_12 GND mn15  l=0.13u w=0.27u m=1
M11 N_10 N_13 N_15 GND mn15  l=0.13u w=0.27u m=1
M12 N_5 CI N_15 GND mn15  l=0.13u w=0.27u m=1
M13 N_13 CI GND GND mn15  l=0.13u w=0.27u m=1
M14 S N_15 VDD VDD mp15  l=0.13u w=0.4u m=1
M15 CO N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_20 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_6 N_11 N_5 VDD mp15  l=0.13u w=0.27u m=1
M19 N_20 B N_5 VDD mp15  l=0.13u w=0.4u m=1
M20 N_11 B VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_10 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 N_11 N_5 N_12 VDD mp15  l=0.13u w=0.27u m=1
M23 N_13 N_10 N_12 VDD mp15  l=0.13u w=0.27u m=1
M24 N_5 N_13 N_15 VDD mp15  l=0.13u w=0.27u m=1
M25 N_10 CI N_15 VDD mp15  l=0.13u w=0.27u m=1
M26 N_13 CI VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ad01d0
* SPICE INPUT		Tue Jul 31 18:28:58 2018	ad01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d1
.subckt ad01d1 GND S CO CI VDD B A
M1 N_2 A GND GND mn15  l=0.13u w=0.38u m=1
M2 N_20 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_20 N_8 N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B N_2 GND mn15  l=0.13u w=0.33u m=1
M5 N_8 B GND GND mn15  l=0.13u w=0.38u m=1
M6 GND N_3 N_6 GND mn15  l=0.13u w=0.38u m=1
M7 N_10 N_3 N_9 GND mn15  l=0.13u w=0.27u m=1
M8 N_8 N_6 N_9 GND mn15  l=0.13u w=0.27u m=1
M9 N_6 N_10 N_12 GND mn15  l=0.13u w=0.27u m=1
M10 N_3 CI N_12 GND mn15  l=0.13u w=0.27u m=1
M11 GND CI N_10 GND mn15  l=0.13u w=0.37u m=1
M12 S N_12 GND GND mn15  l=0.13u w=0.43u m=1
M13 CO N_9 GND GND mn15  l=0.13u w=0.46u m=1
M14 VDD A N_2 VDD mp15  l=0.13u w=0.53u m=1
M15 N_73 N_2 VDD VDD mp15  l=0.13u w=0.66u m=1
M16 N_2 N_8 N_3 VDD mp15  l=0.13u w=0.315u m=1
M17 N_73 B N_3 VDD mp15  l=0.13u w=0.66u m=1
M18 N_8 B VDD VDD mp15  l=0.13u w=0.53u m=1
M19 N_6 N_3 VDD VDD mp15  l=0.13u w=0.53u m=1
M20 N_8 N_3 N_9 VDD mp15  l=0.13u w=0.27u m=1
M21 N_10 N_6 N_9 VDD mp15  l=0.13u w=0.27u m=1
M22 N_3 N_10 N_12 VDD mp15  l=0.13u w=0.27u m=1
M23 N_6 CI N_12 VDD mp15  l=0.13u w=0.27u m=1
M24 N_10 CI VDD VDD mp15  l=0.13u w=0.27u m=1
M25 VDD CI N_10 VDD mp15  l=0.13u w=0.26u m=1
M26 S N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 CO N_9 VDD VDD mp15  l=0.13u w=0.35u m=1
M28 CO N_9 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends ad01d1
* SPICE INPUT		Tue Jul 31 18:29:15 2018	ad01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d2
.subckt ad01d2 VDD S CO GND CI B A
M1 N_3 B N_2 GND mn15  l=0.13u w=0.36u m=1
M2 N_29 N_9 N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.4u m=1
M4 N_29 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_9 N_8 N_19 GND mn15  l=0.13u w=0.36u m=1
M6 N_19 N_3 N_15 GND mn15  l=0.13u w=0.36u m=1
M7 N_8 N_15 N_11 GND mn15  l=0.13u w=0.18u m=1
M8 N_11 N_15 N_8 GND mn15  l=0.13u w=0.18u m=1
M9 N_3 CI N_11 GND mn15  l=0.13u w=0.35u m=1
M10 GND CI N_15 GND mn15  l=0.13u w=0.2u m=1
M11 N_15 CI GND GND mn15  l=0.13u w=0.2u m=1
M12 GND N_11 S GND mn15  l=0.13u w=0.46u m=1
M13 GND N_11 S GND mn15  l=0.13u w=0.46u m=1
M14 GND N_19 CO GND mn15  l=0.13u w=0.46u m=1
M15 CO N_19 GND GND mn15  l=0.13u w=0.46u m=1
M16 N_8 N_3 GND GND mn15  l=0.13u w=0.41u m=1
M17 N_9 B GND GND mn15  l=0.13u w=0.4u m=1
M18 N_23 B N_3 VDD mp15  l=0.13u w=0.66u m=1
M19 N_3 N_9 N_2 VDD mp15  l=0.13u w=0.27u m=1
M20 N_3 N_9 N_2 VDD mp15  l=0.13u w=0.26u m=1
M21 VDD A N_2 VDD mp15  l=0.13u w=0.59u m=1
M22 N_23 N_2 VDD VDD mp15  l=0.13u w=0.66u m=1
M23 N_8 N_3 VDD VDD mp15  l=0.13u w=0.56u m=1
M24 N_9 B VDD VDD mp15  l=0.13u w=0.56u m=1
M25 N_11 CI N_8 VDD mp15  l=0.13u w=0.53u m=1
M26 N_15 CI VDD VDD mp15  l=0.13u w=0.59u m=1
M27 VDD N_11 S VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_11 S VDD mp15  l=0.13u w=0.69u m=1
M29 CO N_19 VDD VDD mp15  l=0.13u w=0.68u m=1
M30 VDD N_19 CO VDD mp15  l=0.13u w=0.69u m=1
M31 N_9 N_3 N_19 VDD mp15  l=0.13u w=0.53u m=1
M32 N_19 N_8 N_15 VDD mp15  l=0.13u w=0.53u m=1
M33 N_3 N_15 N_11 VDD mp15  l=0.13u w=0.49u m=1
.ends ad01d2
* SPICE INPUT		Tue Jul 31 18:29:28 2018	ad01d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01d3
.subckt ad01d3 VDD S CO GND CI B A
M1 N_2 A GND GND mn15  l=0.13u w=0.4u m=1
M2 N_92 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_92 N_9 N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B N_2 GND mn15  l=0.13u w=0.36u m=1
M5 N_9 B GND GND mn15  l=0.13u w=0.4u m=1
M6 N_8 N_3 GND GND mn15  l=0.13u w=0.45u m=1
M7 S N_18 GND GND mn15  l=0.13u w=0.46u m=1
M8 S N_18 GND GND mn15  l=0.13u w=0.46u m=1
M9 S N_18 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_14 N_3 N_15 GND mn15  l=0.13u w=0.36u m=1
M11 N_9 N_8 N_14 GND mn15  l=0.13u w=0.36u m=1
M12 N_3 CI N_18 GND mn15  l=0.13u w=0.35u m=1
M13 N_8 N_15 N_18 GND mn15  l=0.13u w=0.19u m=1
M14 N_18 N_15 N_8 GND mn15  l=0.13u w=0.17u m=1
M15 CO N_14 GND GND mn15  l=0.13u w=0.46u m=1
M16 CO N_14 GND GND mn15  l=0.13u w=0.46u m=1
M17 CO N_14 GND GND mn15  l=0.13u w=0.46u m=1
M18 GND CI N_15 GND mn15  l=0.13u w=0.21u m=1
M19 N_15 CI GND GND mn15  l=0.13u w=0.19u m=1
M20 VDD A N_2 VDD mp15  l=0.13u w=0.58u m=1
M21 N_26 N_2 VDD VDD mp15  l=0.13u w=0.66u m=1
M22 N_3 N_9 N_2 VDD mp15  l=0.13u w=0.27u m=1
M23 N_3 N_9 N_2 VDD mp15  l=0.13u w=0.26u m=1
M24 N_26 B N_3 VDD mp15  l=0.13u w=0.66u m=1
M25 N_9 B VDD VDD mp15  l=0.13u w=0.56u m=1
M26 N_8 N_3 VDD VDD mp15  l=0.13u w=0.56u m=1
M27 S N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 S N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 S N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 N_9 N_3 N_14 VDD mp15  l=0.13u w=0.53u m=1
M31 N_15 N_8 N_14 VDD mp15  l=0.13u w=0.53u m=1
M32 N_18 N_15 N_3 VDD mp15  l=0.13u w=0.49u m=1
M33 N_18 CI N_8 VDD mp15  l=0.13u w=0.53u m=1
M34 CO N_14 VDD VDD mp15  l=0.13u w=0.71u m=1
M35 CO N_14 VDD VDD mp15  l=0.13u w=0.71u m=1
M36 CO N_14 VDD VDD mp15  l=0.13u w=0.65u m=1
M37 N_15 CI VDD VDD mp15  l=0.13u w=0.59u m=1
.ends ad01d3
* SPICE INPUT		Tue Jul 31 18:29:41 2018	ad01dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ad01dm
.subckt ad01dm GND S CO CI VDD B A
M1 S N_17 GND GND mn15  l=0.13u w=0.35u m=1
M2 CO N_14 GND GND mn15  l=0.13u w=0.35u m=1
M3 N_6 CI GND GND mn15  l=0.13u w=0.31u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.31u m=1
M5 N_20 N_7 GND GND mn15  l=0.13u w=0.31u m=1
M6 N_20 N_13 N_8 GND mn15  l=0.13u w=0.31u m=1
M7 N_8 B N_7 GND mn15  l=0.13u w=0.29u m=1
M8 N_13 B GND GND mn15  l=0.13u w=0.31u m=1
M9 GND N_8 N_11 GND mn15  l=0.13u w=0.31u m=1
M10 N_6 N_8 N_14 GND mn15  l=0.13u w=0.29u m=1
M11 N_13 N_11 N_14 GND mn15  l=0.13u w=0.29u m=1
M12 N_11 N_6 N_17 GND mn15  l=0.13u w=0.29u m=1
M13 N_8 CI N_17 GND mn15  l=0.13u w=0.29u m=1
M14 S N_17 VDD VDD mp15  l=0.13u w=0.53u m=1
M15 CO N_14 VDD VDD mp15  l=0.13u w=0.52u m=1
M16 N_6 CI VDD VDD mp15  l=0.13u w=0.48u m=1
M17 N_7 A VDD VDD mp15  l=0.13u w=0.48u m=1
M18 N_27 N_7 VDD VDD mp15  l=0.13u w=0.45u m=1
M19 N_7 N_13 N_8 VDD mp15  l=0.13u w=0.31u m=1
M20 N_27 B N_8 VDD mp15  l=0.13u w=0.45u m=1
M21 N_13 B VDD VDD mp15  l=0.13u w=0.48u m=1
M22 N_11 N_8 VDD VDD mp15  l=0.13u w=0.48u m=1
M23 N_13 N_8 N_14 VDD mp15  l=0.13u w=0.35u m=1
M24 N_6 N_11 N_14 VDD mp15  l=0.13u w=0.35u m=1
M25 N_8 N_6 N_17 VDD mp15  l=0.13u w=0.29u m=1
M26 N_11 CI N_17 VDD mp15  l=0.13u w=0.29u m=1
.ends ad01dm
* SPICE INPUT		Tue Jul 31 18:29:53 2018	adfh01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=adfh01d0
.subckt adfh01d0 GND S CO A B CI VDD
M1 CO N_13 GND GND mn15  l=0.13u w=0.26u m=1
M2 S N_8 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND CI N_5 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M5 N_8 N_14 N_7 GND mn15  l=0.13u w=0.28u m=1
M6 N_13 N_20 N_11 GND mn15  l=0.13u w=0.28u m=1
M7 N_8 N_20 N_5 GND mn15  l=0.13u w=0.28u m=1
M8 N_13 N_14 N_5 GND mn15  l=0.13u w=0.28u m=1
M9 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M10 N_15 N_11 N_14 GND mn15  l=0.13u w=0.3u m=1
M11 N_20 B N_15 GND mn15  l=0.13u w=0.3u m=1
M12 N_14 B N_16 GND mn15  l=0.13u w=0.28u m=1
M13 N_20 N_11 N_16 GND mn15  l=0.13u w=0.28u m=1
M14 N_15 N_21 GND GND mn15  l=0.13u w=0.36u m=1
M15 N_16 A GND GND mn15  l=0.13u w=0.3u m=1
M16 GND A N_21 GND mn15  l=0.13u w=0.18u m=1
M17 CO N_13 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 S N_8 VDD VDD mp15  l=0.13u w=0.4u m=1
M19 VDD CI N_5 VDD mp15  l=0.13u w=0.35u m=1
M20 VDD N_5 N_7 VDD mp15  l=0.13u w=0.35u m=1
M21 N_5 N_14 N_8 VDD mp15  l=0.13u w=0.28u m=1
M22 N_13 N_14 N_11 VDD mp15  l=0.13u w=0.28u m=1
M23 N_7 N_20 N_8 VDD mp15  l=0.13u w=0.28u m=1
M24 N_5 N_20 N_13 VDD mp15  l=0.13u w=0.28u m=1
M25 N_11 B VDD VDD mp15  l=0.13u w=0.35u m=1
M26 VDD B N_11 VDD mp15  l=0.13u w=0.35u m=1
M27 N_16 B N_20 VDD mp15  l=0.13u w=0.4u m=1
M28 N_14 B N_15 VDD mp15  l=0.13u w=0.4u m=1
M29 N_14 N_11 N_16 VDD mp15  l=0.13u w=0.57u m=1
M30 N_20 N_11 N_15 VDD mp15  l=0.13u w=0.56u m=1
M31 N_15 N_21 VDD VDD mp15  l=0.13u w=0.53u m=1
M32 N_21 A VDD VDD mp15  l=0.13u w=0.3u m=1
M33 N_16 A VDD VDD mp15  l=0.13u w=0.46u m=1
.ends adfh01d0
* SPICE INPUT		Tue Jul 31 18:30:06 2018	adfh01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=adfh01d1
.subckt adfh01d1 GND S CO A B CI VDD
M1 N_4 A GND GND mn15  l=0.13u w=0.41u m=1
M2 N_3 A GND GND mn15  l=0.13u w=0.27u m=1
M3 N_8 N_3 GND GND mn15  l=0.13u w=0.41u m=1
M4 N_9 B N_8 GND mn15  l=0.13u w=0.27u m=1
M5 N_6 B N_4 GND mn15  l=0.13u w=0.27u m=1
M6 N_9 N_19 N_4 GND mn15  l=0.13u w=0.27u m=1
M7 CO N_21 GND GND mn15  l=0.13u w=0.46u m=1
M8 S N_16 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND CI N_13 GND mn15  l=0.13u w=0.41u m=1
M10 N_15 N_13 GND GND mn15  l=0.13u w=0.41u m=1
M11 N_16 N_6 N_15 GND mn15  l=0.13u w=0.27u m=1
M12 N_21 N_9 N_19 GND mn15  l=0.13u w=0.27u m=1
M13 N_16 N_9 N_13 GND mn15  l=0.13u w=0.27u m=1
M14 N_21 N_6 N_13 GND mn15  l=0.13u w=0.27u m=1
M15 GND B N_19 GND mn15  l=0.13u w=0.46u m=1
M16 N_8 N_19 N_6 GND mn15  l=0.13u w=0.27u m=1
M17 CO N_21 VDD VDD mp15  l=0.13u w=0.35u m=1
M18 CO N_21 VDD VDD mp15  l=0.13u w=0.35u m=1
M19 S N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_4 A VDD VDD mp15  l=0.13u w=0.59u m=1
M21 N_3 A VDD VDD mp15  l=0.13u w=0.35u m=1
M22 VDD CI N_13 VDD mp15  l=0.13u w=0.59u m=1
M23 VDD N_13 N_15 VDD mp15  l=0.13u w=0.59u m=1
M24 N_13 N_6 N_16 VDD mp15  l=0.13u w=0.4u m=1
M25 N_21 N_6 N_19 VDD mp15  l=0.13u w=0.4u m=1
M26 N_15 N_9 N_16 VDD mp15  l=0.13u w=0.4u m=1
M27 N_13 N_9 N_21 VDD mp15  l=0.13u w=0.4u m=1
M28 N_19 B VDD VDD mp15  l=0.13u w=0.35u m=1
M29 VDD B N_19 VDD mp15  l=0.13u w=0.35u m=1
M30 N_8 N_3 VDD VDD mp15  l=0.13u w=0.59u m=1
M31 N_4 B N_9 VDD mp15  l=0.13u w=0.4u m=1
M32 N_6 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M33 N_6 N_19 N_4 VDD mp15  l=0.13u w=0.4u m=1
M34 N_9 N_19 N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends adfh01d1
* SPICE INPUT		Tue Jul 31 18:30:19 2018	adfh01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=adfh01d2
.subckt adfh01d2 S GND CO VDD CI B A
M1 CO N_26 GND GND mn15  l=0.13u w=0.46u m=1
M2 GND N_26 CO GND mn15  l=0.13u w=0.46u m=1
M3 GND N_10 S GND mn15  l=0.13u w=0.46u m=1
M4 GND N_10 S GND mn15  l=0.13u w=0.46u m=1
M5 GND CI N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_10 N_14 N_9 GND mn15  l=0.13u w=0.41u m=1
M7 N_9 N_7 GND GND mn15  l=0.13u w=0.4u m=1
M8 N_13 A GND GND mn15  l=0.13u w=0.38u m=1
M9 N_12 A GND GND mn15  l=0.13u w=0.27u m=1
M10 N_17 N_12 GND GND mn15  l=0.13u w=0.4u m=1
M11 N_18 B N_17 GND mn15  l=0.13u w=0.41u m=1
M12 N_13 B N_14 GND mn15  l=0.13u w=0.41u m=1
M13 N_18 N_23 N_13 GND mn15  l=0.13u w=0.41u m=1
M14 N_14 N_23 N_17 GND mn15  l=0.13u w=0.41u m=1
M15 GND B N_23 GND mn15  l=0.13u w=0.235u m=1
M16 N_23 B GND GND mn15  l=0.13u w=0.225u m=1
M17 N_26 N_14 N_7 GND mn15  l=0.13u w=0.41u m=1
M18 N_7 N_18 N_10 GND mn15  l=0.13u w=0.41u m=1
M19 N_26 N_18 N_23 GND mn15  l=0.13u w=0.41u m=1
M20 N_13 A VDD VDD mp15  l=0.13u w=0.56u m=1
M21 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M22 VDD N_26 CO VDD mp15  l=0.13u w=0.47u m=1
M23 CO N_26 VDD VDD mp15  l=0.13u w=0.47u m=1
M24 VDD N_26 CO VDD mp15  l=0.13u w=0.46u m=1
M25 VDD N_10 S VDD mp15  l=0.13u w=0.69u m=1
M26 VDD N_10 S VDD mp15  l=0.13u w=0.69u m=1
M27 N_17 N_12 VDD VDD mp15  l=0.13u w=0.59u m=1
M28 N_17 N_23 N_18 VDD mp15  l=0.13u w=0.31u m=1
M29 N_17 N_23 N_18 VDD mp15  l=0.13u w=0.31u m=1
M30 N_18 B N_13 VDD mp15  l=0.13u w=0.62u m=1
M31 N_13 N_23 N_14 VDD mp15  l=0.13u w=0.62u m=1
M32 N_17 B N_14 VDD mp15  l=0.13u w=0.62u m=1
M33 VDD B N_23 VDD mp15  l=0.13u w=0.35u m=1
M34 VDD B N_23 VDD mp15  l=0.13u w=0.35u m=1
M35 N_23 N_14 N_26 VDD mp15  l=0.13u w=0.31u m=1
M36 N_23 N_14 N_26 VDD mp15  l=0.13u w=0.31u m=1
M37 N_7 N_18 N_26 VDD mp15  l=0.13u w=0.62u m=1
M38 N_10 N_18 N_9 VDD mp15  l=0.13u w=0.62u m=1
M39 N_7 N_14 N_10 VDD mp15  l=0.13u w=0.62u m=1
M40 N_7 CI VDD VDD mp15  l=0.13u w=0.59u m=1
M41 N_9 N_7 VDD VDD mp15  l=0.13u w=0.59u m=1
.ends adfh01d2
* SPICE INPUT		Tue Jul 31 18:30:31 2018	ah01d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d0
.subckt ah01d0 GND CO S VDD A B
M1 N_12 B GND GND mn15  l=0.13u w=0.26u m=1
M2 CO N_4 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_12 A N_4 GND mn15  l=0.13u w=0.26u m=1
M4 N_11 B N_9 GND mn15  l=0.13u w=0.26u m=1
M5 N_6 B GND GND mn15  l=0.13u w=0.26u m=1
M6 N_9 N_10 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_11 N_6 N_10 GND mn15  l=0.13u w=0.26u m=1
M8 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M9 GND N_11 S GND mn15  l=0.13u w=0.26u m=1
M10 N_4 B VDD VDD mp15  l=0.13u w=0.4u m=1
M11 CO N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_10 B N_11 VDD mp15  l=0.13u w=0.4u m=1
M14 N_6 B VDD VDD mp15  l=0.13u w=0.4u m=1
M15 N_9 N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_9 N_6 N_11 VDD mp15  l=0.13u w=0.4u m=1
M17 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M18 S N_11 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ah01d0
* SPICE INPUT		Tue Jul 31 18:30:44 2018	ah01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d1
.subckt ah01d1 GND S CO A VDD B
M1 S N_8 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_8 B N_6 GND mn15  l=0.13u w=0.28u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.26u m=1
M4 N_6 N_7 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 N_3 N_7 GND mn15  l=0.13u w=0.28u m=1
M6 N_7 A GND GND mn15  l=0.13u w=0.31u m=1
M7 CO N_11 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_12 B GND GND mn15  l=0.13u w=0.28u m=1
M9 N_12 A N_11 GND mn15  l=0.13u w=0.28u m=1
M10 S N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_7 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M12 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_6 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_8 N_3 N_6 VDD mp15  l=0.13u w=0.38u m=1
M15 N_7 A VDD VDD mp15  l=0.13u w=0.46u m=1
M16 CO N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_11 B VDD VDD mp15  l=0.13u w=0.28u m=1
M18 N_11 A VDD VDD mp15  l=0.13u w=0.28u m=1
.ends ah01d1
* SPICE INPUT		Tue Jul 31 18:31:00 2018	ah01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d2
.subckt ah01d2 GND S CO VDD A B
M1 N_3 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_8 B N_7 GND mn15  l=0.13u w=0.31u m=1
M3 S N_8 GND GND mn15  l=0.13u w=0.46u m=1
M4 S N_8 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_9 N_3 N_8 GND mn15  l=0.13u w=0.36u m=1
M6 N_9 A GND GND mn15  l=0.13u w=0.33u m=1
M7 N_7 N_9 GND GND mn15  l=0.13u w=0.31u m=1
M8 N_14 B GND GND mn15  l=0.13u w=0.47u m=1
M9 N_14 A N_12 GND mn15  l=0.13u w=0.47u m=1
M10 GND N_12 CO GND mn15  l=0.13u w=0.46u m=1
M11 GND N_12 CO GND mn15  l=0.13u w=0.46u m=1
M12 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_9 B N_8 VDD mp15  l=0.13u w=0.52u m=1
M14 S N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 S N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_9 A VDD VDD mp15  l=0.13u w=0.51u m=1
M17 N_7 N_9 VDD VDD mp15  l=0.13u w=0.48u m=1
M18 N_8 N_3 N_7 VDD mp15  l=0.13u w=0.48u m=1
M19 VDD B N_12 VDD mp15  l=0.13u w=0.52u m=1
M20 N_12 A VDD VDD mp15  l=0.13u w=0.26u m=1
M21 N_12 A VDD VDD mp15  l=0.13u w=0.26u m=1
M22 VDD N_12 CO VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_12 CO VDD mp15  l=0.13u w=0.69u m=1
.ends ah01d2
* SPICE INPUT		Tue Jul 31 18:31:18 2018	ah01d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01d3
.subckt ah01d3 GND CO S VDD A B
M1 GND B N_25 GND mn15  l=0.13u w=0.45u m=1
M2 N_24 B GND GND mn15  l=0.13u w=0.21u m=1
M3 GND B N_4 GND mn15  l=0.13u w=0.28u m=1
M4 N_6 A N_25 GND mn15  l=0.13u w=0.36u m=1
M5 N_6 A N_24 GND mn15  l=0.13u w=0.36u m=1
M6 CO N_6 GND GND mn15  l=0.13u w=0.46u m=1
M7 CO N_6 GND GND mn15  l=0.13u w=0.46u m=1
M8 CO N_6 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_13 S GND mn15  l=0.13u w=0.46u m=1
M10 GND N_13 S GND mn15  l=0.13u w=0.46u m=1
M11 GND N_13 S GND mn15  l=0.13u w=0.46u m=1
M12 N_14 B N_13 GND mn15  l=0.13u w=0.27u m=1
M13 N_13 B N_14 GND mn15  l=0.13u w=0.27u m=1
M14 GND N_20 N_14 GND mn15  l=0.13u w=0.25u m=1
M15 N_14 N_20 GND GND mn15  l=0.13u w=0.24u m=1
M16 N_20 N_4 N_13 GND mn15  l=0.13u w=0.27u m=1
M17 N_13 N_4 N_20 GND mn15  l=0.13u w=0.27u m=1
M18 N_20 A GND GND mn15  l=0.13u w=0.3u m=1
M19 N_20 A GND GND mn15  l=0.13u w=0.3u m=1
M20 VDD N_13 S VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_13 S VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_13 S VDD mp15  l=0.13u w=0.69u m=1
M23 VDD B N_6 VDD mp15  l=0.13u w=0.41u m=1
M24 N_6 B VDD VDD mp15  l=0.13u w=0.41u m=1
M25 VDD B N_4 VDD mp15  l=0.13u w=0.4u m=1
M26 N_6 A VDD VDD mp15  l=0.13u w=0.41u m=1
M27 VDD A N_6 VDD mp15  l=0.13u w=0.39u m=1
M28 CO N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 CO N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 CO N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 N_13 N_4 N_14 VDD mp15  l=0.13u w=0.37u m=1
M32 N_13 N_4 N_14 VDD mp15  l=0.13u w=0.325u m=1
M33 N_14 N_20 VDD VDD mp15  l=0.13u w=0.33u m=1
M34 VDD N_20 N_14 VDD mp15  l=0.13u w=0.33u m=1
M35 N_20 B N_13 VDD mp15  l=0.13u w=0.36u m=1
M36 N_20 B N_13 VDD mp15  l=0.13u w=0.34u m=1
M37 VDD A N_20 VDD mp15  l=0.13u w=0.5u m=1
M38 N_20 A VDD VDD mp15  l=0.13u w=0.5u m=1
.ends ah01d3
* SPICE INPUT		Tue Jul 31 18:31:30 2018	ah01dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ah01dm
.subckt ah01dm GND S CO A VDD B
M1 S N_8 GND GND mn15  l=0.13u w=0.35u m=1
M2 N_8 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.26u m=1
M4 N_6 N_7 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 N_3 N_7 GND mn15  l=0.13u w=0.26u m=1
M6 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M7 CO N_11 GND GND mn15  l=0.13u w=0.35u m=1
M8 N_12 B GND GND mn15  l=0.13u w=0.26u m=1
M9 N_12 A N_11 GND mn15  l=0.13u w=0.26u m=1
M10 S N_8 VDD VDD mp15  l=0.13u w=0.53u m=1
M11 N_7 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M12 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_6 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_8 N_3 N_6 VDD mp15  l=0.13u w=0.4u m=1
M15 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M16 CO N_11 VDD VDD mp15  l=0.13u w=0.53u m=1
M17 N_11 B VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_11 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ah01dm
* SPICE INPUT		Tue Jul 31 18:31:43 2018	an02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d0
.subckt an02d0 GND Y VDD A B
M1 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 B N_4 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M5 N_4 B VDD VDD mp15  l=0.13u w=0.325u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.325u m=1
.ends an02d0
* SPICE INPUT		Tue Jul 31 18:31:57 2018	an02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d1
.subckt an02d1 GND Y VDD A B
M1 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_5 B N_4 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M5 N_4 B VDD VDD mp15  l=0.13u w=0.325u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.325u m=1
.ends an02d1
* SPICE INPUT		Tue Jul 31 18:32:10 2018	an02d1p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d1p5
.subckt an02d1p5 GND Y VDD A B
M1 N_5 B N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an02d1p5
* SPICE INPUT		Tue Jul 31 18:32:22 2018	an02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d2
.subckt an02d2 Y GND VDD A B
M1 GND A N_6 GND mn15  l=0.13u w=0.46u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 N_6 B N_4 GND mn15  l=0.13u w=0.46u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.57u m=1
M6 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M8 N_4 B VDD VDD mp15  l=0.13u w=0.57u m=1
.ends an02d2
* SPICE INPUT		Tue Jul 31 18:32:34 2018	an02d2p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d2p5
.subckt an02d2p5 Y GND VDD A B
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_8 B N_5 GND mn15  l=0.13u w=0.46u m=1
M6 N_5 B N_7 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an02d2p5
* SPICE INPUT		Tue Jul 31 18:32:46 2018	an02d3p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d3p5
.subckt an02d3p5 Y GND VDD A B
M1 N_10 B N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_12 B N_4 GND mn15  l=0.13u w=0.46u m=1
M5 N_4 B N_11 GND mn15  l=0.13u w=0.46u m=1
M6 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M14 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD B N_4 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an02d3p5
* SPICE INPUT		Tue Jul 31 18:32:58 2018	an02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02d4
.subckt an02d4 Y GND VDD A B
M1 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_10 B N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_5 B N_9 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_10 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD B N_5 VDD mp15  l=0.13u w=0.345u m=1
M12 VDD A N_5 VDD mp15  l=0.13u w=0.345u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an02d4
* SPICE INPUT		Tue Jul 31 18:33:10 2018	an02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an02dm
.subckt an02dm GND Y VDD A B
M1 N_5 B N_4 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_4 B VDD VDD mp15  l=0.13u w=0.325u m=1
M5 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.325u m=1
.ends an02dm
* SPICE INPUT		Tue Jul 31 18:33:22 2018	an03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d0
.subckt an03d0 GND Y VDD A B C
M1 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_5 C N_4 GND mn15  l=0.13u w=0.26u m=1
M5 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.29u m=1
M7 N_4 B VDD VDD mp15  l=0.13u w=0.29u m=1
M8 N_4 C VDD VDD mp15  l=0.13u w=0.29u m=1
.ends an03d0
* SPICE INPUT		Tue Jul 31 18:33:35 2018	an03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d1
.subckt an03d1 GND Y VDD A B C
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C N_4 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.29u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.29u m=1
M7 N_4 C VDD VDD mp15  l=0.13u w=0.29u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an03d1
* SPICE INPUT		Tue Jul 31 18:33:47 2018	an03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d2
.subckt an03d2 Y GND VDD A B C
M1 N_6 C N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 VDD C N_4 VDD mp15  l=0.13u w=0.51u m=1
M7 N_4 B VDD VDD mp15  l=0.13u w=0.51u m=1
M8 VDD A N_4 VDD mp15  l=0.13u w=0.51u m=1
M9 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends an03d2
* SPICE INPUT		Tue Jul 31 18:34:01 2018	an03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03d4
.subckt an03d4 Y GND VDD A B C
M1 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_10 B N_9 GND mn15  l=0.13u w=0.46u m=1
M3 N_11 C N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_5 C N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_12 B N_11 GND mn15  l=0.13u w=0.46u m=1
M6 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_5 A VDD VDD mp15  l=0.13u w=0.505u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.505u m=1
M13 N_5 C VDD VDD mp15  l=0.13u w=0.505u m=1
M14 N_5 C VDD VDD mp15  l=0.13u w=0.505u m=1
M15 N_5 B VDD VDD mp15  l=0.13u w=0.505u m=1
M16 VDD A N_5 VDD mp15  l=0.13u w=0.505u m=1
M17 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an03d4
* SPICE INPUT		Tue Jul 31 18:34:17 2018	an03dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an03dm
.subckt an03dm GND Y VDD A B C
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C N_4 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.29u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.29u m=1
M7 N_4 C VDD VDD mp15  l=0.13u w=0.29u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends an03dm
* SPICE INPUT		Tue Jul 31 18:34:33 2018	an04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d0
.subckt an04d0 GND Y D C B A VDD
M1 N_5 D N_4 GND mn15  l=0.13u w=0.26u m=1
M2 N_6 C N_5 GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M5 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M6 N_4 D VDD VDD mp15  l=0.13u w=0.26u m=1
M7 VDD C N_4 VDD mp15  l=0.13u w=0.26u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_4 B VDD VDD mp15  l=0.13u w=0.26u m=1
M10 N_4 A VDD VDD mp15  l=0.13u w=0.26u m=1
.ends an04d0
* SPICE INPUT		Tue Jul 31 18:34:47 2018	an04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d1
.subckt an04d1 GND Y VDD A B C D
M1 N_5 D N_4 GND mn15  l=0.13u w=0.36u m=1
M2 N_6 C N_5 GND mn15  l=0.13u w=0.36u m=1
M3 N_7 B N_6 GND mn15  l=0.13u w=0.36u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.36u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_4 D VDD VDD mp15  l=0.13u w=0.36u m=1
M7 N_4 C VDD VDD mp15  l=0.13u w=0.36u m=1
M8 N_4 B VDD VDD mp15  l=0.13u w=0.36u m=1
M9 N_4 A VDD VDD mp15  l=0.13u w=0.36u m=1
M10 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends an04d1
* SPICE INPUT		Tue Jul 31 18:35:00 2018	an04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d2
.subckt an04d2 Y GND VDD A B C D
M1 N_6 D N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 C N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_8 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_4 D VDD VDD mp15  l=0.13u w=0.46u m=1
M8 VDD C N_4 VDD mp15  l=0.13u w=0.46u m=1
M9 N_4 B VDD VDD mp15  l=0.13u w=0.46u m=1
M10 VDD A N_4 VDD mp15  l=0.13u w=0.46u m=1
M11 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends an04d2
* SPICE INPUT		Tue Jul 31 18:35:12 2018	an04d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04d4
.subckt an04d4 Y GND VDD D C B A
M1 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_8 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_8 GND mn15  l=0.13u w=0.46u m=1
M7 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M8 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 C N_7 GND mn15  l=0.13u w=0.46u m=1
M10 N_7 C N_12 GND mn15  l=0.13u w=0.46u m=1
M11 N_13 D N_12 GND mn15  l=0.13u w=0.46u m=1
M12 N_12 D N_13 GND mn15  l=0.13u w=0.46u m=1
M13 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_13 A VDD VDD mp15  l=0.13u w=0.46u m=1
M18 N_13 A VDD VDD mp15  l=0.13u w=0.46u m=1
M19 N_13 B VDD VDD mp15  l=0.13u w=0.46u m=1
M20 N_13 B VDD VDD mp15  l=0.13u w=0.46u m=1
M21 N_13 C VDD VDD mp15  l=0.13u w=0.46u m=1
M22 N_13 C VDD VDD mp15  l=0.13u w=0.46u m=1
M23 VDD D N_13 VDD mp15  l=0.13u w=0.46u m=1
M24 VDD D N_13 VDD mp15  l=0.13u w=0.46u m=1
.ends an04d4
* SPICE INPUT		Tue Jul 31 18:35:25 2018	an04dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=an04dm
.subckt an04dm GND Y VDD A B C D
M1 N_7 B N_6 GND mn15  l=0.13u w=0.3u m=1
M2 N_5 D N_4 GND mn15  l=0.13u w=0.3u m=1
M3 N_6 C N_5 GND mn15  l=0.13u w=0.3u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.3u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.3u m=1
M7 N_4 D VDD VDD mp15  l=0.13u w=0.3u m=1
M8 VDD C N_4 VDD mp15  l=0.13u w=0.3u m=1
M9 N_4 A VDD VDD mp15  l=0.13u w=0.3u m=1
M10 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends an04dm
* SPICE INPUT		Wed Aug  1 08:15:11 2018	antenna
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR


* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d0
.subckt aoi211d0 GND Y VDD D C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y D GND GND mn15  l=0.13u w=0.26u m=1
M4 Y C GND GND mn15  l=0.13u w=0.26u m=1
M5 N_11 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_11 B VDD VDD mp15  l=0.13u w=0.4u m=1
M7 Y D N_14 VDD mp15  l=0.13u w=0.4u m=1
M8 N_11 C N_14 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi211d0
* SPICE INPUT		Tue Jul 31 18:35:58 2018	aoi211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d1
.subckt aoi211d1 Y VDD GND D C B A
M1 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y C GND GND mn15  l=0.13u w=0.26u m=1
M4 Y D GND GND mn15  l=0.13u w=0.26u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_4 C N_6 VDD mp15  l=0.13u w=0.69u m=1
M8 Y D N_6 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi211d1
* SPICE INPUT		Tue Jul 31 18:36:12 2018	aoi211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d2
.subckt aoi211d2 GND Y VDD C D A B
M1 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_8 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND C Y GND mn15  l=0.13u w=0.46u m=1
M6 Y D GND GND mn15  l=0.13u w=0.46u m=1
M7 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_12 B VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_12 B VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_18 C N_12 VDD mp15  l=0.13u w=0.69u m=1
M12 Y D N_17 VDD mp15  l=0.13u w=0.69u m=1
M13 Y D N_18 VDD mp15  l=0.13u w=0.69u m=1
M14 N_12 C N_17 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi211d2
* SPICE INPUT		Tue Jul 31 18:36:31 2018	aoi211d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi211d4
.subckt aoi211d4 GND Y VDD C D A B
M1 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_11 GND mn15  l=0.13u w=0.46u m=1
M4 GND D Y GND mn15  l=0.13u w=0.46u m=1
M5 Y D GND GND mn15  l=0.13u w=0.46u m=1
M6 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_14 B Y GND mn15  l=0.13u w=0.46u m=1
M9 Y B N_13 GND mn15  l=0.13u w=0.46u m=1
M10 Y C GND GND mn15  l=0.13u w=0.46u m=1
M11 Y C GND GND mn15  l=0.13u w=0.46u m=1
M12 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M13 N_20 C N_70 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD B N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_72 D Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y D N_71 VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M20 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD B N_20 VDD mp15  l=0.13u w=0.69u m=1
M22 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_71 C N_20 VDD mp15  l=0.13u w=0.69u m=1
M24 N_73 C N_20 VDD mp15  l=0.13u w=0.69u m=1
M25 N_20 C N_72 VDD mp15  l=0.13u w=0.69u m=1
M26 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 Y D N_70 VDD mp15  l=0.13u w=0.69u m=1
M28 Y D N_73 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi211d4
* SPICE INPUT		Tue Jul 31 18:36:45 2018	aoi21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d0
.subckt aoi21d0 Y VDD GND C B A
M1 N_19 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_19 B Y GND mn15  l=0.13u w=0.26u m=1
M3 Y C GND GND mn15  l=0.13u w=0.26u m=1
M4 VDD A N_2 VDD mp15  l=0.13u w=0.4u m=1
M5 VDD B N_2 VDD mp15  l=0.13u w=0.4u m=1
M6 Y C N_2 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi21d0
* SPICE INPUT		Tue Jul 31 18:36:57 2018	aoi21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d1
.subckt aoi21d1 Y VDD GND C B A
M1 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_19 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y C GND GND mn15  l=0.13u w=0.26u m=1
M4 VDD A N_2 VDD mp15  l=0.13u w=0.69u m=1
M5 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M6 Y C N_2 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21d1
* SPICE INPUT		Tue Jul 31 18:37:09 2018	aoi21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d2
.subckt aoi21d2 GND Y VDD C A B
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M5 Y C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_12 B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_12 B VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21d2
* SPICE INPUT		Tue Jul 31 18:37:22 2018	aoi21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21d4
.subckt aoi21d4 GND Y VDD C A B
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_11 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_13 B Y GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_12 GND mn15  l=0.13u w=0.46u m=1
M8 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M9 Y C GND GND mn15  l=0.13u w=0.31u m=1
M10 Y C GND GND mn15  l=0.13u w=0.31u m=1
M11 Y C GND GND mn15  l=0.13u w=0.31u m=1
M12 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD B N_20 VDD mp15  l=0.13u w=0.69u m=1
M14 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD B N_20 VDD mp15  l=0.13u w=0.69u m=1
M18 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Y C N_20 VDD mp15  l=0.13u w=0.85u m=1
M21 Y C N_20 VDD mp15  l=0.13u w=0.69u m=1
M22 Y C N_20 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21d4
* SPICE INPUT		Tue Jul 31 18:37:34 2018	aoi21dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21dm
.subckt aoi21dm Y VDD GND C B A
M1 N_19 A GND GND mn15  l=0.13u w=0.36u m=1
M2 N_19 B Y GND mn15  l=0.13u w=0.36u m=1
M3 Y C GND GND mn15  l=0.13u w=0.26u m=1
M4 VDD A N_2 VDD mp15  l=0.13u w=0.55u m=1
M5 VDD B N_2 VDD mp15  l=0.13u w=0.55u m=1
M6 Y C N_2 VDD mp15  l=0.13u w=0.55u m=1
.ends aoi21dm
* SPICE INPUT		Tue Jul 31 18:37:46 2018	aoi21md0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21md0
.subckt aoi21md0 GND Y VDD A B CN
M1 GND CN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 GND A N_6 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_3 CN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_10 B VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_10 N_3 Y VDD mp15  l=0.13u w=0.4u m=1
.ends aoi21md0
* SPICE INPUT		Tue Jul 31 18:37:57 2018	aoi21md1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21md1
.subckt aoi21md1 GND Y VDD A B CN
M1 N_3 CN GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_7 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 CN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_11 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M7 N_11 B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21md1
* SPICE INPUT		Tue Jul 31 18:38:09 2018	aoi21md2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21md2
.subckt aoi21md2 GND Y VDD A B CN
M1 N_3 CN GND GND mn15  l=0.13u w=0.3u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M4 Y B N_8 GND mn15  l=0.13u w=0.46u m=1
M5 Y B N_9 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_8 GND mn15  l=0.13u w=0.46u m=1
M7 VDD CN N_3 VDD mp15  l=0.13u w=0.45u m=1
M8 N_13 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M9 Y N_3 N_13 VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_13 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21md2
* SPICE INPUT		Tue Jul 31 18:38:21 2018	aoi21md3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi21md3
.subckt aoi21md3 GND Y VDD B A CN
M1 N_3 CN GND GND mn15  l=0.13u w=0.46u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.31u m=1
M3 Y N_3 GND GND mn15  l=0.13u w=0.31u m=1
M4 Y N_3 GND GND mn15  l=0.13u w=0.31u m=1
M5 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_14 B Y GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_13 GND mn15  l=0.13u w=0.46u m=1
M8 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M10 Y B N_12 GND mn15  l=0.13u w=0.46u m=1
M11 Y B N_15 GND mn15  l=0.13u w=0.46u m=1
M12 GND A N_12 GND mn15  l=0.13u w=0.46u m=1
M13 N_3 CN VDD VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_3 N_22 VDD mp15  l=0.13u w=0.85u m=1
M15 N_22 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M16 N_22 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_22 VDD mp15  l=0.13u w=0.69u m=1
M18 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD B N_22 VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_22 VDD mp15  l=0.13u w=0.69u m=1
M21 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi21md3
* SPICE INPUT		Tue Jul 31 18:38:33 2018	aoi221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d0
.subckt aoi221d0 GND Y VDD E D C A B
M1 N_6 B Y GND mn15  l=0.13u w=0.26u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_7 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 D Y GND mn15  l=0.13u w=0.26u m=1
M5 Y E GND GND mn15  l=0.13u w=0.26u m=1
M6 N_14 B VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_14 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_12 C N_14 VDD mp15  l=0.13u w=0.4u m=1
M9 N_14 D N_12 VDD mp15  l=0.13u w=0.4u m=1
M10 Y E N_12 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi221d0
* SPICE INPUT		Tue Jul 31 18:38:45 2018	aoi221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d1
.subckt aoi221d1 VDD Y GND E D C A B
M1 N_15 B Y GND mn15  l=0.13u w=0.46u m=1
M2 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_16 D Y GND mn15  l=0.13u w=0.46u m=1
M5 Y E GND GND mn15  l=0.13u w=0.26u m=1
M6 N_3 B VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_3 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_3 C N_5 VDD mp15  l=0.13u w=0.69u m=1
M9 N_3 D N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 Y E N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi221d1
* SPICE INPUT		Tue Jul 31 18:38:57 2018	aoi221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d2
.subckt aoi221d2 GND Y VDD E C D A B
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_9 GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_11 D Y GND mn15  l=0.13u w=0.46u m=1
M6 N_12 C GND GND mn15  l=0.13u w=0.46u m=1
M7 N_11 C GND GND mn15  l=0.13u w=0.46u m=1
M8 N_12 D Y GND mn15  l=0.13u w=0.46u m=1
M9 GND E Y GND mn15  l=0.13u w=0.46u m=1
M10 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD B N_22 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD B N_22 VDD mp15  l=0.13u w=0.69u m=1
M13 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_22 D N_19 VDD mp15  l=0.13u w=0.69u m=1
M15 N_22 C N_19 VDD mp15  l=0.13u w=0.69u m=1
M16 N_19 C N_22 VDD mp15  l=0.13u w=0.69u m=1
M17 N_19 D N_22 VDD mp15  l=0.13u w=0.69u m=1
M18 N_19 E Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_19 E Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi221d2
* SPICE INPUT		Tue Jul 31 18:39:09 2018	aoi221d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi221d4
.subckt aoi221d4 Y GND VDD E C D A B
M1 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_14 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_13 GND mn15  l=0.13u w=0.46u m=1
M4 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_16 B Y GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_15 GND mn15  l=0.13u w=0.46u m=1
M8 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND E Y GND mn15  l=0.13u w=0.46u m=1
M10 GND E Y GND mn15  l=0.13u w=0.46u m=1
M11 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M12 N_18 D Y GND mn15  l=0.13u w=0.46u m=1
M13 Y D N_17 GND mn15  l=0.13u w=0.46u m=1
M14 N_19 C GND GND mn15  l=0.13u w=0.46u m=1
M15 N_18 C GND GND mn15  l=0.13u w=0.46u m=1
M16 N_20 D Y GND mn15  l=0.13u w=0.46u m=1
M17 Y D N_19 GND mn15  l=0.13u w=0.46u m=1
M18 N_20 C GND GND mn15  l=0.13u w=0.46u m=1
M19 N_33 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_33 B VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD B N_33 VDD mp15  l=0.13u w=0.69u m=1
M22 N_33 A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 VDD A N_33 VDD mp15  l=0.13u w=0.69u m=1
M24 VDD B N_33 VDD mp15  l=0.13u w=0.69u m=1
M25 VDD B N_33 VDD mp15  l=0.13u w=0.69u m=1
M26 VDD A N_33 VDD mp15  l=0.13u w=0.69u m=1
M27 N_30 E Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y E N_30 VDD mp15  l=0.13u w=0.69u m=1
M29 N_30 E Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_30 E Y VDD mp15  l=0.13u w=0.69u m=1
M31 N_33 C N_30 VDD mp15  l=0.13u w=0.69u m=1
M32 N_33 D N_30 VDD mp15  l=0.13u w=0.69u m=1
M33 N_30 D N_33 VDD mp15  l=0.13u w=0.69u m=1
M34 N_33 C N_30 VDD mp15  l=0.13u w=0.69u m=1
M35 N_30 C N_33 VDD mp15  l=0.13u w=0.69u m=1
M36 N_33 D N_30 VDD mp15  l=0.13u w=0.69u m=1
M37 N_30 D N_33 VDD mp15  l=0.13u w=0.69u m=1
M38 N_30 C N_33 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi221d4
* SPICE INPUT		Tue Jul 31 18:39:23 2018	aoi222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi222d0
.subckt aoi222d0 Y GND VDD F E C D B A
M1 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y F N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y B N_7 GND mn15  l=0.13u w=0.26u m=1
M4 N_8 D Y GND mn15  l=0.13u w=0.26u m=1
M5 N_8 C GND GND mn15  l=0.13u w=0.26u m=1
M6 GND E N_6 GND mn15  l=0.13u w=0.26u m=1
M7 VDD A N_17 VDD mp15  l=0.13u w=0.4u m=1
M8 VDD B N_17 VDD mp15  l=0.13u w=0.4u m=1
M9 N_14 F Y VDD mp15  l=0.13u w=0.4u m=1
M10 N_17 D N_14 VDD mp15  l=0.13u w=0.4u m=1
M11 N_14 C N_17 VDD mp15  l=0.13u w=0.4u m=1
M12 N_14 E Y VDD mp15  l=0.13u w=0.4u m=1
.ends aoi222d0
* SPICE INPUT		Tue Jul 31 18:39:38 2018	aoi222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi222d1
.subckt aoi222d1 Y GND VDD F E C D B A
M1 Y F N_6 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 D Y GND mn15  l=0.13u w=0.46u m=1
M5 N_8 C GND GND mn15  l=0.13u w=0.46u m=1
M6 GND E N_6 GND mn15  l=0.13u w=0.46u m=1
M7 VDD A N_17 VDD mp15  l=0.13u w=0.69u m=1
M8 VDD B N_17 VDD mp15  l=0.13u w=0.69u m=1
M9 N_14 F Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_17 D N_14 VDD mp15  l=0.13u w=0.69u m=1
M11 N_14 C N_17 VDD mp15  l=0.13u w=0.69u m=1
M12 N_14 E Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi222d1
* SPICE INPUT		Tue Jul 31 18:39:53 2018	aoi222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi222d2
.subckt aoi222d2 GND Y VDD E F C D A B
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_11 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_12 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_13 D Y GND mn15  l=0.13u w=0.46u m=1
M7 Y D N_12 GND mn15  l=0.13u w=0.46u m=1
M8 N_13 C GND GND mn15  l=0.13u w=0.46u m=1
M9 N_14 E GND GND mn15  l=0.13u w=0.46u m=1
M10 GND E N_9 GND mn15  l=0.13u w=0.46u m=1
M11 Y F N_9 GND mn15  l=0.13u w=0.46u m=1
M12 Y F N_14 GND mn15  l=0.13u w=0.46u m=1
M13 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD B N_26 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD B N_26 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD A N_26 VDD mp15  l=0.13u w=0.69u m=1
M17 N_26 C N_22 VDD mp15  l=0.13u w=0.69u m=1
M18 N_26 D N_22 VDD mp15  l=0.13u w=0.69u m=1
M19 N_22 D N_26 VDD mp15  l=0.13u w=0.69u m=1
M20 N_22 C N_26 VDD mp15  l=0.13u w=0.69u m=1
M21 Y E N_22 VDD mp15  l=0.13u w=0.69u m=1
M22 N_22 E Y VDD mp15  l=0.13u w=0.69u m=1
M23 N_22 F Y VDD mp15  l=0.13u w=0.69u m=1
M24 N_22 F Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi222d2
* SPICE INPUT		Tue Jul 31 18:40:08 2018	aoi222d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi222d4
.subckt aoi222d4 GND Y A D C B VDD F E
M1 GND E N_15 GND mn15  l=0.13u w=0.46u m=1
M2 Y F N_15 GND mn15  l=0.13u w=0.46u m=1
M3 Y F N_26 GND mn15  l=0.13u w=0.46u m=1
M4 N_26 E GND GND mn15  l=0.13u w=0.46u m=1
M5 N_25 E GND GND mn15  l=0.13u w=0.46u m=1
M6 N_25 F Y GND mn15  l=0.13u w=0.46u m=1
M7 Y F N_24 GND mn15  l=0.13u w=0.46u m=1
M8 N_24 E GND GND mn15  l=0.13u w=0.46u m=1
M9 N_23 C GND GND mn15  l=0.13u w=0.46u m=1
M10 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M11 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M12 Y D N_22 GND mn15  l=0.13u w=0.46u m=1
M13 N_22 C GND GND mn15  l=0.13u w=0.46u m=1
M14 N_21 C GND GND mn15  l=0.13u w=0.46u m=1
M15 N_21 D Y GND mn15  l=0.13u w=0.46u m=1
M16 Y D N_20 GND mn15  l=0.13u w=0.46u m=1
M17 N_20 C GND GND mn15  l=0.13u w=0.46u m=1
M18 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M19 N_19 B Y GND mn15  l=0.13u w=0.46u m=1
M20 Y B N_18 GND mn15  l=0.13u w=0.46u m=1
M21 N_18 A GND GND mn15  l=0.13u w=0.46u m=1
M22 N_17 A GND GND mn15  l=0.13u w=0.46u m=1
M23 N_17 B Y GND mn15  l=0.13u w=0.46u m=1
M24 Y B N_16 GND mn15  l=0.13u w=0.46u m=1
M25 N_47 E Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_47 F Y VDD mp15  l=0.13u w=0.69u m=1
M27 N_47 F Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y E N_47 VDD mp15  l=0.13u w=0.69u m=1
M29 N_47 E Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y F N_47 VDD mp15  l=0.13u w=0.69u m=1
M31 N_47 F Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y E N_47 VDD mp15  l=0.13u w=0.69u m=1
M33 N_47 C N_41 VDD mp15  l=0.13u w=0.69u m=1
M34 N_41 D N_47 VDD mp15  l=0.13u w=0.69u m=1
M35 N_47 D N_41 VDD mp15  l=0.13u w=0.69u m=1
M36 N_41 C N_47 VDD mp15  l=0.13u w=0.69u m=1
M37 N_47 C N_41 VDD mp15  l=0.13u w=0.69u m=1
M38 N_41 D N_47 VDD mp15  l=0.13u w=0.69u m=1
M39 N_47 D N_41 VDD mp15  l=0.13u w=0.69u m=1
M40 N_41 C N_47 VDD mp15  l=0.13u w=0.69u m=1
M41 N_41 A VDD VDD mp15  l=0.13u w=0.69u m=1
M42 VDD A N_41 VDD mp15  l=0.13u w=0.69u m=1
M43 VDD B N_41 VDD mp15  l=0.13u w=0.69u m=1
M44 VDD B N_41 VDD mp15  l=0.13u w=0.69u m=1
M45 N_41 A VDD VDD mp15  l=0.13u w=0.69u m=1
M46 VDD A N_41 VDD mp15  l=0.13u w=0.69u m=1
M47 N_41 B VDD VDD mp15  l=0.13u w=0.69u m=1
M48 VDD B N_41 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi222d4
* SPICE INPUT		Tue Jul 31 18:40:20 2018	aoi22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d0
.subckt aoi22d0 GND Y VDD C D B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y D N_5 GND mn15  l=0.13u w=0.26u m=1
M4 GND C N_5 GND mn15  l=0.13u w=0.26u m=1
M5 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_10 B VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_10 D Y VDD mp15  l=0.13u w=0.4u m=1
M8 Y C N_10 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi22d0
* SPICE INPUT		Tue Jul 31 18:40:33 2018	aoi22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d1
.subckt aoi22d1 GND Y VDD C D B A
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 Y D N_5 GND mn15  l=0.13u w=0.46u m=1
M4 GND C N_5 GND mn15  l=0.13u w=0.46u m=1
M5 VDD A N_10 VDD mp15  l=0.13u w=0.69u m=1
M6 N_10 B VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_10 D Y VDD mp15  l=0.13u w=0.69u m=1
M8 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi22d1
* SPICE INPUT		Tue Jul 31 18:40:46 2018	aoi22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d2
.subckt aoi22d2 GND Y VDD D C A B
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_9 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_8 GND mn15  l=0.13u w=0.46u m=1
M4 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_10 C GND GND mn15  l=0.13u w=0.46u m=1
M6 Y D N_7 GND mn15  l=0.13u w=0.46u m=1
M7 Y D N_10 GND mn15  l=0.13u w=0.46u m=1
M8 N_7 C GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M10 VDD B N_16 VDD mp15  l=0.13u w=0.69u m=1
M11 N_16 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y C N_16 VDD mp15  l=0.13u w=0.69u m=1
M14 N_16 D Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_16 D Y VDD mp15  l=0.13u w=0.69u m=1
M16 N_16 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi22d2
* SPICE INPUT		Tue Jul 31 18:40:59 2018	aoi22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22d4
.subckt aoi22d4 GND Y VDD D C A B
M1 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_12 GND mn15  l=0.13u w=0.46u m=1
M4 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_15 B Y GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_14 GND mn15  l=0.13u w=0.46u m=1
M8 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M10 N_17 D Y GND mn15  l=0.13u w=0.46u m=1
M11 Y D N_16 GND mn15  l=0.13u w=0.46u m=1
M12 N_18 C GND GND mn15  l=0.13u w=0.46u m=1
M13 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M14 Y D N_11 GND mn15  l=0.13u w=0.46u m=1
M15 Y D N_18 GND mn15  l=0.13u w=0.46u m=1
M16 N_11 C GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD A N_28 VDD mp15  l=0.13u w=0.69u m=1
M18 VDD B N_28 VDD mp15  l=0.13u w=0.69u m=1
M19 N_28 B VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_28 VDD mp15  l=0.13u w=0.69u m=1
M21 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD B N_28 VDD mp15  l=0.13u w=0.69u m=1
M23 N_28 B VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 Y C N_28 VDD mp15  l=0.13u w=0.69u m=1
M26 Y D N_28 VDD mp15  l=0.13u w=0.69u m=1
M27 N_28 D Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y C N_28 VDD mp15  l=0.13u w=0.69u m=1
M29 N_28 C Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_28 D Y VDD mp15  l=0.13u w=0.69u m=1
M31 N_28 D Y VDD mp15  l=0.13u w=0.69u m=1
M32 N_28 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi22d4
* SPICE INPUT		Tue Jul 31 18:41:11 2018	aoi22dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi22dm
.subckt aoi22dm GND Y VDD C D B A
M1 N_6 A GND GND mn15  l=0.13u w=0.36u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.36u m=1
M3 Y D N_5 GND mn15  l=0.13u w=0.36u m=1
M4 GND C N_5 GND mn15  l=0.13u w=0.36u m=1
M5 N_10 A VDD VDD mp15  l=0.13u w=0.55u m=1
M6 N_10 B VDD VDD mp15  l=0.13u w=0.55u m=1
M7 N_10 D Y VDD mp15  l=0.13u w=0.55u m=1
M8 N_10 C Y VDD mp15  l=0.13u w=0.55u m=1
.ends aoi22dm
* SPICE INPUT		Tue Jul 31 18:41:24 2018	aoi2m1d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi2m1d0
.subckt aoi2m1d0 Y GND VDD C A BN
M1 N_5 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 N_5 Y GND mn15  l=0.13u w=0.26u m=1
M4 GND C Y GND mn15  l=0.13u w=0.26u m=1
M5 VDD BN N_5 VDD mp15  l=0.13u w=0.4u m=1
M6 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 VDD N_5 N_10 VDD mp15  l=0.13u w=0.4u m=1
M8 Y C N_10 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi2m1d0
* SPICE INPUT		Tue Jul 31 18:41:39 2018	aoi2m1d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi2m1d1
.subckt aoi2m1d1 GND Y VDD C A BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_7 N_3 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND C Y GND mn15  l=0.13u w=0.26u m=1
M5 N_3 BN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 VDD A N_11 VDD mp15  l=0.13u w=0.69u m=1
M7 VDD N_3 N_11 VDD mp15  l=0.13u w=0.69u m=1
M8 Y C N_11 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi2m1d1
* SPICE INPUT		Tue Jul 31 18:41:58 2018	aoi2m1d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi2m1d2
.subckt aoi2m1d2 GND Y VDD C A BN
M1 GND BN N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_8 N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_4 N_7 GND mn15  l=0.13u w=0.46u m=1
M5 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M6 Y C GND GND mn15  l=0.13u w=0.46u m=1
M7 VDD BN N_4 VDD mp15  l=0.13u w=0.69u m=1
M8 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_4 N_13 VDD mp15  l=0.13u w=0.69u m=1
M10 N_13 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
M13 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi2m1d2
* SPICE INPUT		Tue Jul 31 18:42:12 2018	aoi2m1d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi2m1d4
.subckt aoi2m1d4 Y GND VDD C A BN
M1 N_6 BN GND GND mn15  l=0.13u w=0.46u m=1
M2 N_6 BN GND GND mn15  l=0.13u w=0.46u m=1
M3 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_12 N_6 Y GND mn15  l=0.13u w=0.46u m=1
M5 Y N_6 N_11 GND mn15  l=0.13u w=0.46u m=1
M6 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_14 N_6 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_6 N_13 GND mn15  l=0.13u w=0.46u m=1
M10 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M11 GND C Y GND mn15  l=0.13u w=0.46u m=1
M12 GND C Y GND mn15  l=0.13u w=0.46u m=1
M13 VDD BN N_6 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD BN N_6 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_6 N_20 VDD mp15  l=0.13u w=0.69u m=1
M17 N_20 N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M19 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_6 N_20 VDD mp15  l=0.13u w=0.69u m=1
M21 N_20 N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_20 C Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y C N_20 VDD mp15  l=0.13u w=0.69u m=1
M25 N_20 C Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_20 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi2m1d4
* SPICE INPUT		Tue Jul 31 18:42:24 2018	aoi31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d0
.subckt aoi31d0 GND Y VDD D C B A
M1 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y D GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 C Y GND mn15  l=0.13u w=0.26u m=1
M5 N_11 A VDD VDD mp15  l=0.13u w=0.35u m=1
M6 Y D N_11 VDD mp15  l=0.13u w=0.4u m=1
M7 VDD B N_11 VDD mp15  l=0.13u w=0.38u m=1
M8 VDD C N_11 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi31d0
* SPICE INPUT		Tue Jul 31 18:42:36 2018	aoi31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d1
.subckt aoi31d1 GND Y VDD D C B A
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_6 B N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M4 Y D GND GND mn15  l=0.13u w=0.26u m=1
M5 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 VDD B N_11 VDD mp15  l=0.13u w=0.69u m=1
M7 VDD C N_11 VDD mp15  l=0.13u w=0.69u m=1
M8 Y D N_11 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi31d1
* SPICE INPUT		Tue Jul 31 18:42:48 2018	aoi31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d2
.subckt aoi31d2 GND Y C B A D VDD
M1 Y D GND GND mn15  l=0.13u w=0.46u m=1
M2 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_9 B N_8 GND mn15  l=0.13u w=0.46u m=1
M4 Y C N_7 GND mn15  l=0.13u w=0.46u m=1
M5 N_8 C Y GND mn15  l=0.13u w=0.46u m=1
M6 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M7 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_18 D Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_18 D Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_18 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_18 C VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_18 C VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_18 B VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi31d2
* SPICE INPUT		Tue Jul 31 18:43:00 2018	aoi31d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31d4
.subckt aoi31d4 GND Y VDD D C B A
M1 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_2 B N_3 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M9 Y C N_3 GND mn15  l=0.13u w=0.46u m=1
M10 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M11 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M12 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M13 Y D GND GND mn15  l=0.13u w=0.46u m=1
M14 Y D GND GND mn15  l=0.13u w=0.46u m=1
M15 N_19 A VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_19 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_19 VDD mp15  l=0.13u w=0.69u m=1
M18 N_19 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_19 B VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_19 B VDD VDD mp15  l=0.13u w=0.61u m=1
M21 N_19 B VDD VDD mp15  l=0.13u w=0.61u m=1
M22 VDD B N_19 VDD mp15  l=0.13u w=0.61u m=1
M23 VDD C N_19 VDD mp15  l=0.13u w=0.575u m=1
M24 VDD C N_19 VDD mp15  l=0.13u w=0.575u m=1
M25 N_19 C VDD VDD mp15  l=0.13u w=0.575u m=1
M26 VDD C N_19 VDD mp15  l=0.13u w=0.575u m=1
M27 N_19 C VDD VDD mp15  l=0.13u w=0.575u m=1
M28 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M29 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M31 Y D N_19 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi31d4
* SPICE INPUT		Tue Jul 31 18:43:11 2018	aoi31dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi31dm
.subckt aoi31dm GND Y VDD D C B A
M1 N_5 A GND GND mn15  l=0.13u w=0.36u m=1
M2 N_6 B N_5 GND mn15  l=0.13u w=0.36u m=1
M3 N_6 C Y GND mn15  l=0.13u w=0.36u m=1
M4 Y D GND GND mn15  l=0.13u w=0.26u m=1
M5 N_11 A VDD VDD mp15  l=0.13u w=0.55u m=1
M6 VDD B N_11 VDD mp15  l=0.13u w=0.55u m=1
M7 VDD C N_11 VDD mp15  l=0.13u w=0.55u m=1
M8 Y D N_11 VDD mp15  l=0.13u w=0.55u m=1
.ends aoi31dm
* SPICE INPUT		Tue Jul 31 18:43:23 2018	aoi32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d0
.subckt aoi32d0 GND Y VDD D E C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y C N_7 GND mn15  l=0.13u w=0.26u m=1
M4 Y E N_5 GND mn15  l=0.13u w=0.26u m=1
M5 GND D N_5 GND mn15  l=0.13u w=0.26u m=1
M6 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_13 B VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_13 C VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_13 E Y VDD mp15  l=0.13u w=0.4u m=1
M10 N_13 D Y VDD mp15  l=0.13u w=0.4u m=1
.ends aoi32d0
* SPICE INPUT		Tue Jul 31 18:43:36 2018	aoi32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d1
.subckt aoi32d1 GND Y VDD D E C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_7 C Y GND mn15  l=0.13u w=0.46u m=1
M4 Y E N_5 GND mn15  l=0.13u w=0.36u m=1
M5 GND D N_5 GND mn15  l=0.13u w=0.36u m=1
M6 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 VDD B N_13 VDD mp15  l=0.13u w=0.69u m=1
M8 N_13 C VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_13 E Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_13 D Y VDD mp15  l=0.13u w=0.69u m=1
.ends aoi32d1
* SPICE INPUT		Tue Jul 31 18:43:47 2018	aoi32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d2
.subckt aoi32d2 GND Y VDD D E A B C
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_9 B N_8 GND mn15  l=0.13u w=0.46u m=1
M3 GND D N_7 GND mn15  l=0.13u w=0.36u m=1
M4 Y E N_7 GND mn15  l=0.13u w=0.36u m=1
M5 Y E N_12 GND mn15  l=0.13u w=0.36u m=1
M6 N_12 D GND GND mn15  l=0.13u w=0.36u m=1
M7 N_10 C Y GND mn15  l=0.13u w=0.46u m=1
M8 Y C N_9 GND mn15  l=0.13u w=0.46u m=1
M9 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M10 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M11 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_21 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_21 D Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_21 E Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_21 E Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y D N_21 VDD mp15  l=0.13u w=0.69u m=1
M17 N_21 C VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_21 C VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD B N_21 VDD mp15  l=0.13u w=0.69u m=1
M20 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi32d2
* SPICE INPUT		Tue Jul 31 18:43:59 2018	aoi32d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32d4
.subckt aoi32d4 GND Y D E C VDD B A
M1 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_2 B N_3 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 D GND GND mn15  l=0.13u w=0.36u m=1
M10 N_12 D GND GND mn15  l=0.13u w=0.36u m=1
M11 N_12 D GND GND mn15  l=0.13u w=0.36u m=1
M12 GND D N_12 GND mn15  l=0.13u w=0.36u m=1
M13 Y C N_3 GND mn15  l=0.13u w=0.46u m=1
M14 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M15 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M16 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M17 N_12 E Y GND mn15  l=0.13u w=0.48u m=1
M18 N_12 E Y GND mn15  l=0.13u w=0.48u m=1
M19 N_12 E Y GND mn15  l=0.13u w=0.48u m=1
M20 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD A N_24 VDD mp15  l=0.13u w=0.69u m=1
M23 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_24 B VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_24 B VDD VDD mp15  l=0.13u w=0.61u m=1
M26 N_24 B VDD VDD mp15  l=0.13u w=0.61u m=1
M27 VDD B N_24 VDD mp15  l=0.13u w=0.61u m=1
M28 N_24 D Y VDD mp15  l=0.13u w=0.69u m=1
M29 N_24 D Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_24 D Y VDD mp15  l=0.13u w=0.69u m=1
M31 Y D N_24 VDD mp15  l=0.13u w=0.69u m=1
M32 N_24 C VDD VDD mp15  l=0.13u w=0.575u m=1
M33 VDD C N_24 VDD mp15  l=0.13u w=0.575u m=1
M34 N_24 C VDD VDD mp15  l=0.13u w=0.575u m=1
M35 VDD C N_24 VDD mp15  l=0.13u w=0.575u m=1
M36 N_24 C VDD VDD mp15  l=0.13u w=0.575u m=1
M37 N_24 E Y VDD mp15  l=0.13u w=0.605u m=1
M38 Y E N_24 VDD mp15  l=0.13u w=0.605u m=1
M39 N_24 E Y VDD mp15  l=0.13u w=0.605u m=1
M40 N_24 E Y VDD mp15  l=0.13u w=0.645u m=1
.ends aoi32d4
* SPICE INPUT		Tue Jul 31 18:44:11 2018	aoi32dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi32dm
.subckt aoi32dm GND Y VDD D E C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.36u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.36u m=1
M3 N_7 C Y GND mn15  l=0.13u w=0.36u m=1
M4 Y E N_5 GND mn15  l=0.13u w=0.3u m=1
M5 GND D N_5 GND mn15  l=0.13u w=0.3u m=1
M6 N_13 A VDD VDD mp15  l=0.13u w=0.55u m=1
M7 N_13 B VDD VDD mp15  l=0.13u w=0.55u m=1
M8 N_13 C VDD VDD mp15  l=0.13u w=0.55u m=1
M9 N_13 E Y VDD mp15  l=0.13u w=0.55u m=1
M10 N_13 D Y VDD mp15  l=0.13u w=0.55u m=1
.ends aoi32dm
* SPICE INPUT		Tue Jul 31 18:44:23 2018	aoi33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d0
.subckt aoi33d0 GND Y VDD D E F C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y C N_7 GND mn15  l=0.13u w=0.26u m=1
M4 N_8 F Y GND mn15  l=0.13u w=0.26u m=1
M5 N_8 E N_5 GND mn15  l=0.13u w=0.26u m=1
M6 GND D N_5 GND mn15  l=0.13u w=0.26u m=1
M7 N_15 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_15 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_15 C VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y F N_15 VDD mp15  l=0.13u w=0.4u m=1
M11 Y E N_15 VDD mp15  l=0.13u w=0.4u m=1
M12 Y D N_15 VDD mp15  l=0.13u w=0.4u m=1
.ends aoi33d0
* SPICE INPUT		Tue Jul 31 18:44:36 2018	aoi33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d1
.subckt aoi33d1 GND Y VDD D E F C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 Y C N_7 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 F Y GND mn15  l=0.13u w=0.46u m=1
M5 N_8 E N_5 GND mn15  l=0.13u w=0.46u m=1
M6 GND D N_5 GND mn15  l=0.13u w=0.46u m=1
M7 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_15 B VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_15 C VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y F N_15 VDD mp15  l=0.13u w=0.69u m=1
M11 Y E N_15 VDD mp15  l=0.13u w=0.69u m=1
M12 Y D N_15 VDD mp15  l=0.13u w=0.69u m=1
.ends aoi33d1
* SPICE INPUT		Tue Jul 31 18:44:51 2018	aoi33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d2
.subckt aoi33d2 Y GND A C D E VDD B F
M1 Y F N_10 GND mn15  l=0.13u w=0.46u m=1
M2 N_11 F Y GND mn15  l=0.13u w=0.46u m=1
M3 N_11 E N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 E N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_2 D GND GND mn15  l=0.13u w=0.46u m=1
M7 GND D N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_13 B N_12 GND mn15  l=0.13u w=0.46u m=1
M9 GND A N_15 GND mn15  l=0.13u w=0.46u m=1
M10 N_15 B N_14 GND mn15  l=0.13u w=0.46u m=1
M11 Y C N_13 GND mn15  l=0.13u w=0.46u m=1
M12 N_14 C Y GND mn15  l=0.13u w=0.46u m=1
M13 Y F N_28 VDD mp15  l=0.13u w=0.565u m=1
M14 Y F N_28 VDD mp15  l=0.13u w=0.405u m=1
M15 N_28 F Y VDD mp15  l=0.13u w=0.41u m=1
M16 VDD A N_28 VDD mp15  l=0.13u w=0.69u m=1
M17 N_28 E Y VDD mp15  l=0.13u w=0.69u m=1
M18 N_28 D Y VDD mp15  l=0.13u w=0.69u m=1
M19 Y D N_28 VDD mp15  l=0.13u w=0.69u m=1
M20 N_28 B VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 Y E N_28 VDD mp15  l=0.13u w=0.69u m=1
M23 VDD B N_28 VDD mp15  l=0.13u w=0.69u m=1
M24 N_28 C VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_28 C VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi33d2
* SPICE INPUT		Tue Jul 31 18:45:05 2018	aoi33d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoi33d4
.subckt aoi33d4 GND Y VDD A B C F E D
M1 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 B N_3 GND mn15  l=0.13u w=0.46u m=1
M5 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_12 F Y GND mn15  l=0.13u w=0.46u m=1
M10 Y F N_12 GND mn15  l=0.13u w=0.46u m=1
M11 N_12 F Y GND mn15  l=0.13u w=0.46u m=1
M12 N_12 F Y GND mn15  l=0.13u w=0.46u m=1
M13 Y C N_3 GND mn15  l=0.13u w=0.46u m=1
M14 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M15 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M16 N_3 C Y GND mn15  l=0.13u w=0.46u m=1
M17 N_21 D GND GND mn15  l=0.13u w=0.46u m=1
M18 N_21 D GND GND mn15  l=0.13u w=0.46u m=1
M19 N_21 D GND GND mn15  l=0.13u w=0.46u m=1
M20 N_21 D GND GND mn15  l=0.13u w=0.46u m=1
M21 N_21 E N_12 GND mn15  l=0.13u w=0.46u m=1
M22 N_12 E N_21 GND mn15  l=0.13u w=0.46u m=1
M23 N_12 E N_21 GND mn15  l=0.13u w=0.46u m=1
M24 N_12 E N_21 GND mn15  l=0.13u w=0.46u m=1
M25 Y D N_35 VDD mp15  l=0.13u w=0.69u m=1
M26 N_35 D Y VDD mp15  l=0.13u w=0.69u m=1
M27 N_35 D Y VDD mp15  l=0.13u w=0.69u m=1
M28 N_35 D Y VDD mp15  l=0.13u w=0.69u m=1
M29 N_35 E Y VDD mp15  l=0.13u w=0.575u m=1
M30 N_35 E Y VDD mp15  l=0.13u w=0.55u m=1
M31 Y E N_35 VDD mp15  l=0.13u w=0.545u m=1
M32 N_35 E Y VDD mp15  l=0.13u w=0.545u m=1
M33 Y E N_35 VDD mp15  l=0.13u w=0.545u m=1
M34 N_35 F Y VDD mp15  l=0.13u w=0.56u m=1
M35 N_35 F Y VDD mp15  l=0.13u w=0.565u m=1
M36 N_35 F Y VDD mp15  l=0.13u w=0.545u m=1
M37 Y F N_35 VDD mp15  l=0.13u w=0.545u m=1
M38 N_35 F Y VDD mp15  l=0.13u w=0.545u m=1
M39 N_35 C VDD VDD mp15  l=0.13u w=0.545u m=1
M40 N_35 C VDD VDD mp15  l=0.13u w=0.555u m=1
M41 N_35 C VDD VDD mp15  l=0.13u w=0.555u m=1
M42 VDD C N_35 VDD mp15  l=0.13u w=0.555u m=1
M43 N_35 C VDD VDD mp15  l=0.13u w=0.555u m=1
M44 N_35 B VDD VDD mp15  l=0.13u w=0.6u m=1
M45 N_35 B VDD VDD mp15  l=0.13u w=0.6u m=1
M46 VDD B N_35 VDD mp15  l=0.13u w=0.6u m=1
M47 N_35 B VDD VDD mp15  l=0.13u w=0.69u m=1
M48 N_35 B VDD VDD mp15  l=0.13u w=0.265u m=1
M49 N_35 A VDD VDD mp15  l=0.13u w=0.69u m=1
M50 VDD A N_35 VDD mp15  l=0.13u w=0.69u m=1
M51 VDD A N_35 VDD mp15  l=0.13u w=0.69u m=1
M52 N_35 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoi33d4
* SPICE INPUT		Tue Jul 31 18:45:20 2018	aoim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d0
.subckt aoim21d0 Y VDD AN C GND BN
M1 GND BN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 GND N_3 Y GND mn15  l=0.13u w=0.26u m=1
M3 GND C Y GND mn15  l=0.13u w=0.26u m=1
M4 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M5 N_8 BN N_3 VDD mp15  l=0.13u w=0.4u m=1
M6 VDD N_3 N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 Y C N_7 VDD mp15  l=0.13u w=0.4u m=1
M8 VDD AN N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends aoim21d0
* SPICE INPUT		Tue Jul 31 18:45:34 2018	aoim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d1
.subckt aoim21d1 Y VDD GND C AN BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_3 Y GND mn15  l=0.13u w=0.35u m=1
M4 GND C Y GND mn15  l=0.13u w=0.35u m=1
M5 N_6 BN N_3 VDD mp15  l=0.13u w=0.52u m=1
M6 VDD AN N_6 VDD mp15  l=0.13u w=0.52u m=1
M7 VDD N_3 N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 Y C N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends aoim21d1
* SPICE INPUT		Tue Jul 31 18:45:47 2018	aoim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d2
.subckt aoim21d2 VDD Y GND C AN BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.36u m=1
M2 GND AN N_3 GND mn15  l=0.13u w=0.36u m=1
M3 Y N_3 GND GND mn15  l=0.13u w=0.36u m=1
M4 GND C Y GND mn15  l=0.13u w=0.36u m=1
M5 GND C Y GND mn15  l=0.13u w=0.36u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.36u m=1
M7 N_7 BN N_3 VDD mp15  l=0.13u w=0.69u m=1
M8 VDD AN N_7 VDD mp15  l=0.13u w=0.69u m=1
M9 N_8 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y C N_6 VDD mp15  l=0.13u w=0.69u m=1
M11 Y C N_8 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_3 N_6 VDD mp15  l=0.13u w=0.69u m=1
.ends aoim21d2
* SPICE INPUT		Tue Jul 31 18:45:59 2018	aoim21d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21d3
.subckt aoim21d3 VDD Y GND C AN BN
M1 N_4 AN GND GND mn15  l=0.13u w=0.35u m=1
M2 N_4 BN GND GND mn15  l=0.13u w=0.35u m=1
M3 N_4 BN GND GND mn15  l=0.13u w=0.33u m=1
M4 GND AN N_4 GND mn15  l=0.13u w=0.33u m=1
M5 Y C GND GND mn15  l=0.13u w=0.46u m=1
M6 Y C GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND C Y GND mn15  l=0.13u w=0.46u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M11 N_10 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_11 BN N_4 VDD mp15  l=0.13u w=0.69u m=1
M13 N_4 BN N_10 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD AN N_11 VDD mp15  l=0.13u w=0.69u m=1
M15 N_12 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
M17 N_13 C Y VDD mp15  l=0.13u w=0.62u m=1
M18 N_14 N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
M19 VDD N_4 N_13 VDD mp15  l=0.13u w=0.62u m=1
M20 Y C N_9 VDD mp15  l=0.13u w=0.685u m=1
M21 N_14 C Y VDD mp15  l=0.13u w=0.695u m=1
M22 N_9 N_4 VDD VDD mp15  l=0.13u w=0.685u m=1
.ends aoim21d3
* SPICE INPUT		Tue Jul 31 18:46:11 2018	aoim21dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim21dm
.subckt aoim21dm Y VDD GND C AN BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_3 Y GND mn15  l=0.13u w=0.28u m=1
M4 GND C Y GND mn15  l=0.13u w=0.28u m=1
M5 N_8 BN N_3 VDD mp15  l=0.13u w=0.4u m=1
M6 VDD AN N_8 VDD mp15  l=0.13u w=0.4u m=1
M7 VDD N_3 N_7 VDD mp15  l=0.13u w=0.55u m=1
M8 Y C N_7 VDD mp15  l=0.13u w=0.55u m=1
.ends aoim21dm
* SPICE INPUT		Tue Jul 31 18:46:24 2018	aoim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d0
.subckt aoim22d0 GND Y VDD C D BN AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 BN GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M4 Y D N_7 GND mn15  l=0.13u w=0.26u m=1
M5 GND C N_7 GND mn15  l=0.13u w=0.26u m=1
M6 VDD AN N_32 VDD mp15  l=0.13u w=0.4u m=1
M7 N_5 BN N_32 VDD mp15  l=0.13u w=0.4u m=1
M8 N_11 N_5 Y VDD mp15  l=0.13u w=0.4u m=1
M9 N_11 D VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_11 C VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aoim22d0
* SPICE INPUT		Tue Jul 31 18:46:36 2018	aoim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d1
.subckt aoim22d1 GND Y C D VDD BN AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 BN GND GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_7 GND mn15  l=0.13u w=0.46u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M5 Y D N_7 GND mn15  l=0.13u w=0.46u m=1
M6 VDD AN N_32 VDD mp15  l=0.13u w=0.52u m=1
M7 N_32 BN N_5 VDD mp15  l=0.13u w=0.52u m=1
M8 N_11 C VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_11 N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M10 N_11 D VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoim22d1
* SPICE INPUT		Tue Jul 31 18:46:50 2018	aoim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d2
.subckt aoim22d2 GND Y VDD C D BN AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.36u m=1
M2 N_5 BN GND GND mn15  l=0.13u w=0.36u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M4 GND C N_9 GND mn15  l=0.13u w=0.47u m=1
M5 N_10 C GND GND mn15  l=0.13u w=0.45u m=1
M6 Y D N_9 GND mn15  l=0.13u w=0.47u m=1
M7 Y D N_10 GND mn15  l=0.13u w=0.45u m=1
M8 VDD AN N_20 VDD mp15  l=0.13u w=0.69u m=1
M9 N_20 BN N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 N_14 C VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_14 N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
M13 N_14 C VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_14 D VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_14 D VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoim22d2
* SPICE INPUT		Tue Jul 31 18:47:10 2018	aoim22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22d4
.subckt aoim22d4 GND Y VDD AN BN C D
M1 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M2 N_15 D Y GND mn15  l=0.13u w=0.46u m=1
M3 Y D N_14 GND mn15  l=0.13u w=0.46u m=1
M4 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_15 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_17 D Y GND mn15  l=0.13u w=0.46u m=1
M7 Y D N_16 GND mn15  l=0.13u w=0.46u m=1
M8 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M10 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_3 AN GND GND mn15  l=0.13u w=0.35u m=1
M12 GND AN N_3 GND mn15  l=0.13u w=0.35u m=1
M13 N_3 BN GND GND mn15  l=0.13u w=0.35u m=1
M14 GND BN N_3 GND mn15  l=0.13u w=0.35u m=1
M15 VDD C N_25 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD D N_25 VDD mp15  l=0.13u w=0.69u m=1
M17 N_25 D VDD VDD mp15  l=0.13u w=0.69u m=1
M18 VDD C N_25 VDD mp15  l=0.13u w=0.69u m=1
M19 N_25 C VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD D N_25 VDD mp15  l=0.13u w=0.69u m=1
M21 N_25 D VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_25 C VDD VDD mp15  l=0.13u w=0.69u m=1
M23 Y N_3 N_25 VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_3 N_25 VDD mp15  l=0.13u w=0.69u m=1
M25 N_25 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_25 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M27 N_31 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M28 N_3 BN N_30 VDD mp15  l=0.13u w=0.69u m=1
M29 N_3 BN N_31 VDD mp15  l=0.13u w=0.69u m=1
M30 N_30 AN VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aoim22d4
* SPICE INPUT		Tue Jul 31 18:47:24 2018	aoim22dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aoim22dm
.subckt aoim22dm GND Y C D VDD BN AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 BN GND GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_7 GND mn15  l=0.13u w=0.36u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M5 Y D N_7 GND mn15  l=0.13u w=0.36u m=1
M6 VDD AN N_32 VDD mp15  l=0.13u w=0.34u m=1
M7 N_32 BN N_5 VDD mp15  l=0.13u w=0.34u m=1
M8 N_11 C VDD VDD mp15  l=0.13u w=0.55u m=1
M9 N_11 N_5 Y VDD mp15  l=0.13u w=0.55u m=1
M10 N_11 D VDD VDD mp15  l=0.13u w=0.55u m=1
.ends aoim22dm
* SPICE INPUT		Tue Jul 31 18:47:36 2018	aor211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d0
.subckt aor211d0 Y GND VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 C GND GND mn15  l=0.13u w=0.26u m=1
M3 N_7 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.26u m=1
M6 N_16 D N_5 VDD mp15  l=0.13u w=0.38u m=1
M7 N_16 C N_11 VDD mp15  l=0.13u w=0.38u m=1
M8 N_11 B VDD VDD mp15  l=0.13u w=0.38u m=1
M9 N_11 A VDD VDD mp15  l=0.13u w=0.38u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor211d0
* SPICE INPUT		Tue Jul 31 18:47:47 2018	aor211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d1
.subckt aor211d1 GND Y VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 C GND GND mn15  l=0.13u w=0.26u m=1
M3 N_7 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_16 D N_5 VDD mp15  l=0.13u w=0.38u m=1
M7 N_16 C N_11 VDD mp15  l=0.13u w=0.38u m=1
M8 N_11 B VDD VDD mp15  l=0.13u w=0.38u m=1
M9 N_11 A VDD VDD mp15  l=0.13u w=0.38u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor211d1
* SPICE INPUT		Tue Jul 31 18:47:59 2018	aor211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d2
.subckt aor211d2 Y GND A B C D VDD
M1 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_6 D GND GND mn15  l=0.13u w=0.26u m=1
M4 N_6 C GND GND mn15  l=0.13u w=0.26u m=1
M5 N_9 B N_6 GND mn15  l=0.13u w=0.46u m=1
M6 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M7 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_6 D N_37 VDD mp15  l=0.13u w=0.69u m=1
M10 N_13 C N_37 VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
.ends aor211d2
* SPICE INPUT		Tue Jul 31 18:48:13 2018	aor211d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor211d4
.subckt aor211d4 GND Y VDD C D A B
M1 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 B N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B N_12 GND mn15  l=0.13u w=0.46u m=1
M4 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND C N_3 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 D GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M10 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M11 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_17 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_17 B VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_25 C N_17 VDD mp15  l=0.13u w=0.69u m=1
M16 N_3 D N_24 VDD mp15  l=0.13u w=0.69u m=1
M17 N_3 D N_25 VDD mp15  l=0.13u w=0.69u m=1
M18 N_17 C N_24 VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor211d4
* SPICE INPUT		Tue Jul 31 18:48:25 2018	aor21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d0
.subckt aor21d0 GND Y VDD C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_10 A VDD VDD mp15  l=0.13u w=0.38u m=1
M6 VDD B N_10 VDD mp15  l=0.13u w=0.38u m=1
M7 N_5 C N_10 VDD mp15  l=0.13u w=0.38u m=1
M8 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor21d0
* SPICE INPUT		Tue Jul 31 18:48:36 2018	aor21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d1
.subckt aor21d1 GND Y VDD C B A
M1 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 B N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_10 A VDD VDD mp15  l=0.13u w=0.38u m=1
M6 VDD B N_10 VDD mp15  l=0.13u w=0.38u m=1
M7 N_5 C N_10 VDD mp15  l=0.13u w=0.38u m=1
M8 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor21d1
* SPICE INPUT		Tue Jul 31 18:48:48 2018	aor21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d2
.subckt aor21d2 GND Y VDD C B A
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_8 B N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 C GND GND mn15  l=0.13u w=0.26u m=1
M4 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M6 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M7 VDD B N_12 VDD mp15  l=0.13u w=0.69u m=1
M8 N_3 C N_12 VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor21d2
* SPICE INPUT		Tue Jul 31 18:49:02 2018	aor21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor21d4
.subckt aor21d4 GND Y VDD C A B
M1 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 B N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B N_11 GND mn15  l=0.13u w=0.46u m=1
M4 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M7 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M8 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M10 VDD A N_17 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD B N_17 VDD mp15  l=0.13u w=0.69u m=1
M12 N_17 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_17 C N_3 VDD mp15  l=0.13u w=0.69u m=1
M15 N_17 C N_3 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M19 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor21d4
* SPICE INPUT		Tue Jul 31 18:49:17 2018	aor221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d0
.subckt aor221d0 GND Y VDD E D C A B
M1 N_8 B N_3 GND mn15  l=0.13u w=0.26u m=1
M2 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_9 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_9 D N_3 GND mn15  l=0.13u w=0.26u m=1
M5 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_15 B VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_15 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_15 C N_14 VDD mp15  l=0.13u w=0.4u m=1
M10 N_14 D N_15 VDD mp15  l=0.13u w=0.4u m=1
M11 N_3 E N_14 VDD mp15  l=0.13u w=0.4u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor221d0
* SPICE INPUT		Tue Jul 31 18:49:31 2018	aor221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d1
.subckt aor221d1 GND Y VDD E D C A B
M1 N_8 B N_3 GND mn15  l=0.13u w=0.26u m=1
M2 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_9 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_9 D N_3 GND mn15  l=0.13u w=0.26u m=1
M5 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_15 B VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_15 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_15 C N_14 VDD mp15  l=0.13u w=0.4u m=1
M10 N_14 D N_15 VDD mp15  l=0.13u w=0.4u m=1
M11 N_3 E N_14 VDD mp15  l=0.13u w=0.4u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor221d1
* SPICE INPUT		Tue Jul 31 18:49:44 2018	aor221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d2
.subckt aor221d2 GND Y VDD E C D B A
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 B N_10 GND mn15  l=0.13u w=0.46u m=1
M3 N_4 D N_9 GND mn15  l=0.13u w=0.46u m=1
M4 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_4 E GND GND mn15  l=0.13u w=0.26u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M9 N_16 B VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_16 D N_15 VDD mp15  l=0.13u w=0.69u m=1
M11 N_15 C N_16 VDD mp15  l=0.13u w=0.69u m=1
M12 N_4 E N_15 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor221d2
* SPICE INPUT		Tue Jul 31 18:50:00 2018	aor221d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor221d4
.subckt aor221d4 Y GND D C B E A VDD
M1 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M2 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M5 N_8 E GND GND mn15  l=0.13u w=0.46u m=1
M6 N_16 D N_8 GND mn15  l=0.13u w=0.46u m=1
M7 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M8 N_15 C GND GND mn15  l=0.13u w=0.46u m=1
M9 N_15 D N_8 GND mn15  l=0.13u w=0.46u m=1
M10 N_8 B N_14 GND mn15  l=0.13u w=0.46u m=1
M11 N_13 B N_8 GND mn15  l=0.13u w=0.46u m=1
M12 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M13 N_13 A GND GND mn15  l=0.13u w=0.46u m=1
M14 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M17 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_8 E N_27 VDD mp15  l=0.13u w=0.69u m=1
M19 N_27 E N_8 VDD mp15  l=0.13u w=0.69u m=1
M20 N_27 D N_22 VDD mp15  l=0.13u w=0.69u m=1
M21 N_22 C N_27 VDD mp15  l=0.13u w=0.69u m=1
M22 N_22 C N_27 VDD mp15  l=0.13u w=0.69u m=1
M23 N_27 D N_22 VDD mp15  l=0.13u w=0.69u m=1
M24 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor221d4
* SPICE INPUT		Tue Jul 31 18:50:15 2018	aor222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor222d0
.subckt aor222d0 GND Y A D B VDD C E F
M1 N_9 F N_2 GND mn15  l=0.13u w=0.26u m=1
M2 N_9 E GND GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_8 GND mn15  l=0.13u w=0.26u m=1
M4 N_2 D N_8 GND mn15  l=0.13u w=0.26u m=1
M5 N_10 B N_2 GND mn15  l=0.13u w=0.26u m=1
M6 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_2 F N_19 VDD mp15  l=0.13u w=0.4u m=1
M9 N_19 E N_2 VDD mp15  l=0.13u w=0.4u m=1
M10 N_19 C N_15 VDD mp15  l=0.13u w=0.4u m=1
M11 N_15 D N_19 VDD mp15  l=0.13u w=0.4u m=1
M12 N_15 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_15 A VDD VDD mp15  l=0.13u w=0.4u m=1
M14 Y N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor222d0
* SPICE INPUT		Tue Jul 31 18:50:26 2018	aor222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor222d1
.subckt aor222d1 GND Y VDD B A D C E F
M1 N_9 F N_2 GND mn15  l=0.13u w=0.26u m=1
M2 N_9 E GND GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_8 GND mn15  l=0.13u w=0.26u m=1
M4 N_2 D N_8 GND mn15  l=0.13u w=0.26u m=1
M5 N_10 B N_2 GND mn15  l=0.13u w=0.26u m=1
M6 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_2 F N_19 VDD mp15  l=0.13u w=0.4u m=1
M9 N_19 E N_2 VDD mp15  l=0.13u w=0.4u m=1
M10 N_19 C N_17 VDD mp15  l=0.13u w=0.4u m=1
M11 N_17 D N_19 VDD mp15  l=0.13u w=0.4u m=1
M12 N_17 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_17 A VDD VDD mp15  l=0.13u w=0.4u m=1
M14 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor222d1
* SPICE INPUT		Tue Jul 31 18:50:37 2018	aor222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor222d2
.subckt aor222d2 GND Y VDD A B D C E F
M1 N_10 F N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_10 E GND GND mn15  l=0.13u w=0.46u m=1
M3 GND C N_9 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 D N_9 GND mn15  l=0.13u w=0.46u m=1
M5 N_11 B N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_2 F N_19 VDD mp15  l=0.13u w=0.69u m=1
M10 N_19 E N_2 VDD mp15  l=0.13u w=0.69u m=1
M11 N_19 C N_17 VDD mp15  l=0.13u w=0.69u m=1
M12 N_19 D N_17 VDD mp15  l=0.13u w=0.69u m=1
M13 N_17 B VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_17 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor222d2
* SPICE INPUT		Tue Jul 31 18:50:50 2018	aor222d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor222d4
.subckt aor222d4 Y GND VDD A B D C E F
M1 N_13 E GND GND mn15  l=0.13u w=0.46u m=1
M2 N_14 F N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_5 F N_13 GND mn15  l=0.13u w=0.46u m=1
M4 N_14 E GND GND mn15  l=0.13u w=0.46u m=1
M5 N_15 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_16 D N_5 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 D N_15 GND mn15  l=0.13u w=0.46u m=1
M8 N_16 C GND GND mn15  l=0.13u w=0.46u m=1
M9 N_17 A GND GND mn15  l=0.13u w=0.46u m=1
M10 N_18 B N_5 GND mn15  l=0.13u w=0.46u m=1
M11 N_5 B N_17 GND mn15  l=0.13u w=0.46u m=1
M12 N_18 A GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M15 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M16 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M17 N_5 E N_30 VDD mp15  l=0.13u w=0.69u m=1
M18 N_5 F N_30 VDD mp15  l=0.13u w=0.69u m=1
M19 N_30 F N_5 VDD mp15  l=0.13u w=0.69u m=1
M20 N_30 E N_5 VDD mp15  l=0.13u w=0.69u m=1
M21 N_27 C N_30 VDD mp15  l=0.13u w=0.69u m=1
M22 N_30 D N_27 VDD mp15  l=0.13u w=0.69u m=1
M23 N_30 D N_27 VDD mp15  l=0.13u w=0.69u m=1
M24 N_30 C N_27 VDD mp15  l=0.13u w=0.69u m=1
M25 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_27 B VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_27 B VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD A N_27 VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor222d4
* SPICE INPUT		Tue Jul 31 18:51:01 2018	aor22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d0
.subckt aor22d0 GND Y VDD A B D C
M1 GND C N_7 GND mn15  l=0.13u w=0.26u m=1
M2 N_2 D N_7 GND mn15  l=0.13u w=0.26u m=1
M3 N_8 B N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_2 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_13 C N_2 VDD mp15  l=0.13u w=0.4u m=1
M7 N_13 D N_2 VDD mp15  l=0.13u w=0.4u m=1
M8 N_13 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor22d0
* SPICE INPUT		Tue Jul 31 18:51:13 2018	aor22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d1
.subckt aor22d1 GND Y VDD A B D C
M1 GND C N_7 GND mn15  l=0.13u w=0.26u m=1
M2 N_2 D N_7 GND mn15  l=0.13u w=0.26u m=1
M3 N_8 B N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_13 C N_2 VDD mp15  l=0.13u w=0.4u m=1
M7 N_13 D N_2 VDD mp15  l=0.13u w=0.4u m=1
M8 N_13 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor22d1
* SPICE INPUT		Tue Jul 31 18:51:26 2018	aor22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d2
.subckt aor22d2 Y GND VDD A B D C
M1 N_8 B N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND C N_9 GND mn15  l=0.13u w=0.46u m=1
M6 N_4 D N_9 GND mn15  l=0.13u w=0.46u m=1
M7 N_14 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M8 N_4 D N_14 VDD mp15  l=0.13u w=0.69u m=1
M9 N_14 B VDD VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_14 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor22d2
* SPICE INPUT		Tue Jul 31 18:51:37 2018	aor22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor22d4
.subckt aor22d4 GND Y VDD A B C D
M1 N_13 C GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 D N_12 GND mn15  l=0.13u w=0.46u m=1
M3 N_4 D N_13 GND mn15  l=0.13u w=0.46u m=1
M4 N_12 C GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M10 N_15 B N_4 GND mn15  l=0.13u w=0.46u m=1
M11 N_4 B N_14 GND mn15  l=0.13u w=0.46u m=1
M12 N_15 A GND GND mn15  l=0.13u w=0.46u m=1
M13 N_4 C N_22 VDD mp15  l=0.13u w=0.69u m=1
M14 N_22 D N_4 VDD mp15  l=0.13u w=0.69u m=1
M15 N_22 D N_4 VDD mp15  l=0.13u w=0.69u m=1
M16 N_22 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_22 B VDD VDD mp15  l=0.13u w=0.69u m=1
M24 VDD A N_22 VDD mp15  l=0.13u w=0.69u m=1
.ends aor22d4
* SPICE INPUT		Tue Jul 31 18:51:50 2018	aor31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d0
.subckt aor31d0 GND Y VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 C N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_12 D N_5 VDD mp15  l=0.13u w=0.4u m=1
M7 N_12 C VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_12 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends aor31d0
* SPICE INPUT		Tue Jul 31 18:52:02 2018	aor31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d1
.subckt aor31d1 GND Y VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 C N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_12 D N_5 VDD mp15  l=0.13u w=0.4u m=1
M7 N_12 C VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_12 B VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor31d1
* SPICE INPUT		Tue Jul 31 18:52:15 2018	aor31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d2
.subckt aor31d2 Y GND VDD A B C D
M1 N_5 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_7 C N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_13 D N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_13 C VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_13 B VDD VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
.ends aor31d2
* SPICE INPUT		Tue Jul 31 18:52:29 2018	aor31d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=aor31d4
.subckt aor31d4 GND Y VDD D A B C
M1 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 B N_11 GND mn15  l=0.13u w=0.46u m=1
M3 N_13 C N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C N_12 GND mn15  l=0.13u w=0.46u m=1
M5 N_14 B N_13 GND mn15  l=0.13u w=0.46u m=1
M6 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_3 D GND GND mn15  l=0.13u w=0.46u m=1
M8 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M11 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_20 C VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_20 C VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 B VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_3 D N_20 VDD mp15  l=0.13u w=0.69u m=1
M19 N_20 D N_3 VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M23 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends aor31d4
* SPICE INPUT		Tue Jul 31 18:52:45 2018	bh01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=bh01d1
.subckt bh01d1 VDD Y GND
M1 GND Y N_4 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 N_6 GND mn15  l=0.13u w=0.26u m=1
M3 GND N_4 N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_4 Y VDD VDD mp15  l=0.13u w=0.4u m=1
M5 Y N_4 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends bh01d1
* SPICE INPUT		Tue Jul 31 18:52:59 2018	buffd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd0
.subckt buffd0 GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends buffd0
* SPICE INPUT		Tue Jul 31 18:53:12 2018	buffd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd1
.subckt buffd1 GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd1
* SPICE INPUT		Tue Jul 31 18:53:29 2018	buffd12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd12
.subckt buffd12 Y GND VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M16 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M18 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M20 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd12
* SPICE INPUT		Tue Jul 31 18:53:41 2018	buffd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd16
.subckt buffd16 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M6 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M16 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M17 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M18 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M19 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M20 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M21 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M22 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M23 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M24 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M26 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M28 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M33 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M34 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M36 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M37 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M38 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M40 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M42 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M43 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M44 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd16
* SPICE INPUT		Tue Jul 31 18:53:53 2018	buffd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd2
.subckt buffd2 Y GND VDD A
M1 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M6 VDD A N_4 VDD mp15  l=0.13u w=0.55u m=1
.ends buffd2
* SPICE INPUT		Tue Jul 31 18:54:05 2018	buffd20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd20
.subckt buffd20 Y GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M4 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M6 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M11 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M12 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M13 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M14 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M15 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M16 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M17 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M18 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M19 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M20 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M21 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M22 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M23 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M24 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M25 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M26 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M27 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M28 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M29 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M30 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M31 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M32 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M33 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M34 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M36 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M37 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M38 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M40 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M42 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M43 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M44 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M45 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M46 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M47 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M48 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M49 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M50 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M51 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M52 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M53 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M54 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd20
* SPICE INPUT		Tue Jul 31 18:54:17 2018	buffd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd3
.subckt buffd3 GND Y VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd3
* SPICE INPUT		Tue Jul 31 18:54:29 2018	buffd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd4
.subckt buffd4 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.35u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.34u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M7 VDD A N_5 VDD mp15  l=0.13u w=0.54u m=1
M8 N_5 A VDD VDD mp15  l=0.13u w=0.54u m=1
M9 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd4
* SPICE INPUT		Tue Jul 31 18:54:40 2018	buffd5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd5
.subckt buffd5 GND Y VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M8 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M9 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd5
* SPICE INPUT		Tue Jul 31 18:54:52 2018	buffd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd6
.subckt buffd6 Y GND VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd6
* SPICE INPUT		Tue Jul 31 18:55:04 2018	buffd7
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd7
.subckt buffd7 GND Y VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.4u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.39u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.39u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 VDD A N_5 VDD mp15  l=0.13u w=0.6u m=1
M12 N_5 A VDD VDD mp15  l=0.13u w=0.6u m=1
M13 VDD A N_5 VDD mp15  l=0.13u w=0.6u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd7
* SPICE INPUT		Tue Jul 31 18:55:15 2018	buffd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffd8
.subckt buffd8 Y GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M11 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M12 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M13 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buffd8
* SPICE INPUT		Tue Jul 31 18:55:27 2018	buffdm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buffdm
.subckt buffdm VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends buffdm
* SPICE INPUT		Tue Jul 31 18:55:40 2018	buftd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd0
.subckt buftd0 GND Y VDD E A
M1 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_6 N_7 GND mn15  l=0.13u w=0.5u m=1
M4 Y E N_7 GND mn15  l=0.13u w=0.5u m=1
M5 VDD A N_6 VDD mp15  l=0.13u w=0.4u m=1
M6 N_14 N_6 VDD VDD mp15  l=0.13u w=0.53u m=1
M7 N_15 N_3 Y VDD mp15  l=0.13u w=0.27u m=1
M8 N_14 N_3 Y VDD mp15  l=0.13u w=0.53u m=1
M9 N_15 N_6 VDD VDD mp15  l=0.13u w=0.27u m=1
M10 N_3 E VDD VDD mp15  l=0.13u w=0.4u m=1
.ends buftd0
* SPICE INPUT		Tue Jul 31 18:55:54 2018	buftd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd1
.subckt buftd1 VDD Y GND E A
M1 N_4 A GND GND mn15  l=0.13u w=0.32u m=1
M2 N_14 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_15 E Y GND mn15  l=0.13u w=0.46u m=1
M4 Y E N_14 GND mn15  l=0.13u w=0.46u m=1
M5 N_15 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 E GND GND mn15  l=0.13u w=0.32u m=1
M7 VDD A N_4 VDD mp15  l=0.13u w=0.48u m=1
M8 N_7 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_8 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y N_3 N_7 VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_3 E VDD VDD mp15  l=0.13u w=0.48u m=1
.ends buftd1
* SPICE INPUT		Tue Jul 31 18:56:09 2018	buftd12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd12
.subckt buftd12 GND Y VDD A E
M1 N_5 E GND GND mn15  l=0.13u w=0.42u m=1
M2 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 A GND GND mn15  l=0.13u w=0.42u m=1
M7 N_2 E N_3 GND mn15  l=0.13u w=0.4u m=1
M8 N_2 E N_3 GND mn15  l=0.13u w=0.4u m=1
M9 N_3 E N_2 GND mn15  l=0.13u w=0.4u m=1
M10 N_3 N_5 GND GND mn15  l=0.13u w=0.38u m=1
M11 N_3 N_5 GND GND mn15  l=0.13u w=0.38u m=1
M12 N_3 N_5 GND GND mn15  l=0.13u w=0.38u m=1
M13 Y N_3 GND GND mn15  l=0.13u w=0.425u m=1
M14 Y N_3 GND GND mn15  l=0.13u w=0.425u m=1
M15 Y N_3 GND GND mn15  l=0.13u w=0.425u m=1
M16 GND N_3 Y GND mn15  l=0.13u w=0.425u m=1
M17 Y N_3 GND GND mn15  l=0.13u w=0.405u m=1
M18 Y N_3 GND GND mn15  l=0.13u w=0.455u m=1
M19 Y N_3 GND GND mn15  l=0.13u w=0.455u m=1
M20 Y N_3 GND GND mn15  l=0.13u w=0.455u m=1
M21 Y N_3 GND GND mn15  l=0.13u w=0.455u m=1
M22 Y N_3 GND GND mn15  l=0.13u w=0.4u m=1
M23 Y N_3 GND GND mn15  l=0.13u w=0.4u m=1
M24 GND N_3 Y GND mn15  l=0.13u w=0.4u m=1
M25 Y N_3 GND GND mn15  l=0.13u w=0.365u m=1
M26 VDD E N_5 VDD mp15  l=0.13u w=0.315u m=1
M27 N_5 E VDD VDD mp15  l=0.13u w=0.315u m=1
M28 N_2 A VDD VDD mp15  l=0.13u w=0.685u m=1
M29 N_2 A VDD VDD mp15  l=0.13u w=0.685u m=1
M30 N_2 A VDD VDD mp15  l=0.13u w=0.685u m=1
M31 N_2 A VDD VDD mp15  l=0.13u w=0.685u m=1
M32 N_2 A VDD VDD mp15  l=0.13u w=0.56u m=1
M33 N_2 E VDD VDD mp15  l=0.13u w=0.605u m=1
M34 N_2 E VDD VDD mp15  l=0.13u w=0.605u m=1
M35 VDD E N_2 VDD mp15  l=0.13u w=0.465u m=1
M36 N_2 N_5 N_3 VDD mp15  l=0.13u w=0.79u m=1
M37 N_3 N_5 N_2 VDD mp15  l=0.13u w=0.8u m=1
M38 N_3 N_5 N_2 VDD mp15  l=0.13u w=0.79u m=1
M39 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M40 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M41 Y N_2 VDD VDD mp15  l=0.13u w=0.71u m=1
M42 Y N_2 VDD VDD mp15  l=0.13u w=0.71u m=1
M43 VDD N_2 Y VDD mp15  l=0.13u w=0.71u m=1
M44 Y N_2 VDD VDD mp15  l=0.13u w=0.71u m=1
M45 VDD N_2 Y VDD mp15  l=0.13u w=0.71u m=1
M46 Y N_2 VDD VDD mp15  l=0.13u w=0.71u m=1
M47 VDD N_2 Y VDD mp15  l=0.13u w=0.71u m=1
M48 Y N_2 VDD VDD mp15  l=0.13u w=0.68u m=1
M49 VDD N_2 Y VDD mp15  l=0.13u w=0.67u m=1
M50 Y N_2 VDD VDD mp15  l=0.13u w=0.58u m=1
.ends buftd12
* SPICE INPUT		Tue Jul 31 18:56:22 2018	buftd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd16
.subckt buftd16 GND Y VDD E A
M1 GND A N_2 GND mn15  l=0.13u w=0.43u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M3 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M4 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M5 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M6 N_2 A GND GND mn15  l=0.13u w=0.4u m=1
M7 N_2 A GND GND mn15  l=0.13u w=0.37u m=1
M8 N_2 N_14 GND GND mn15  l=0.13u w=0.37u m=1
M9 N_2 N_14 GND GND mn15  l=0.13u w=0.37u m=1
M10 GND N_14 N_2 GND mn15  l=0.13u w=0.37u m=1
M11 GND N_14 N_2 GND mn15  l=0.13u w=0.35u m=1
M12 GND E N_14 GND mn15  l=0.13u w=0.44u m=1
M13 N_17 E N_2 GND mn15  l=0.13u w=0.55u m=1
M14 N_2 E N_17 GND mn15  l=0.13u w=0.55u m=1
M15 N_2 E N_17 GND mn15  l=0.13u w=0.48u m=1
M16 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M17 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M18 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M19 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M20 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M21 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M22 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M23 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M24 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M25 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M26 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M27 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M28 Y N_2 GND GND mn15  l=0.13u w=0.4u m=1
M29 Y N_2 GND GND mn15  l=0.13u w=0.4u m=1
M30 GND N_2 Y GND mn15  l=0.13u w=0.4u m=1
M31 Y N_2 GND GND mn15  l=0.13u w=0.4u m=1
M32 Y N_2 GND GND mn15  l=0.13u w=0.36u m=1
M33 N_17 A VDD VDD mp15  l=0.13u w=0.65u m=1
M34 VDD A N_17 VDD mp15  l=0.13u w=0.65u m=1
M35 N_17 A VDD VDD mp15  l=0.13u w=0.65u m=1
M36 VDD A N_17 VDD mp15  l=0.13u w=0.65u m=1
M37 N_17 A VDD VDD mp15  l=0.13u w=0.65u m=1
M38 VDD A N_17 VDD mp15  l=0.13u w=0.65u m=1
M39 N_17 A VDD VDD mp15  l=0.13u w=0.64u m=1
M40 N_17 E VDD VDD mp15  l=0.13u w=0.76u m=1
M41 N_17 E VDD VDD mp15  l=0.13u w=0.76u m=1
M42 VDD E N_17 VDD mp15  l=0.13u w=0.73u m=1
M43 N_14 E VDD VDD mp15  l=0.13u w=0.67u m=1
M44 N_2 N_14 N_17 VDD mp15  l=0.13u w=0.56u m=1
M45 N_17 N_14 N_2 VDD mp15  l=0.13u w=0.56u m=1
M46 N_17 N_14 N_2 VDD mp15  l=0.13u w=0.56u m=1
M47 N_2 N_14 N_17 VDD mp15  l=0.13u w=0.56u m=1
M48 N_17 N_14 N_2 VDD mp15  l=0.13u w=0.56u m=1
M49 N_2 N_14 N_17 VDD mp15  l=0.13u w=0.28u m=1
M50 Y N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M51 Y N_17 VDD VDD mp15  l=0.13u w=0.67u m=1
M52 Y N_17 VDD VDD mp15  l=0.13u w=0.67u m=1
M53 VDD N_17 Y VDD mp15  l=0.13u w=0.67u m=1
M54 Y N_17 VDD VDD mp15  l=0.13u w=0.67u m=1
M55 VDD N_17 Y VDD mp15  l=0.13u w=0.69u m=1
M56 VDD N_17 Y VDD mp15  l=0.13u w=0.69u m=1
M57 Y N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M58 VDD N_17 Y VDD mp15  l=0.13u w=0.69u m=1
M59 Y N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M60 VDD N_17 Y VDD mp15  l=0.13u w=0.69u m=1
M61 Y N_17 VDD VDD mp15  l=0.13u w=0.65u m=1
M62 Y N_17 VDD VDD mp15  l=0.13u w=0.62u m=1
M63 VDD N_17 Y VDD mp15  l=0.13u w=0.57u m=1
M64 Y N_17 VDD VDD mp15  l=0.13u w=0.57u m=1
M65 VDD N_17 Y VDD mp15  l=0.13u w=0.57u m=1
M66 Y N_17 VDD VDD mp15  l=0.13u w=0.57u m=1
.ends buftd16
* SPICE INPUT		Tue Jul 31 18:56:36 2018	buftd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd2
.subckt buftd2 GND Y VDD E A
M1 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 E GND GND mn15  l=0.13u w=0.46u m=1
M3 N_6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_6 E Y GND mn15  l=0.13u w=0.565u m=1
M8 N_6 E Y GND mn15  l=0.13u w=0.565u m=1
M9 N_6 E Y GND mn15  l=0.13u w=0.43u m=1
M10 Y E N_6 GND mn15  l=0.13u w=0.29u m=1
M11 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD E N_3 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_4 N_15 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_4 N_15 VDD mp15  l=0.13u w=0.69u m=1
M15 N_15 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_4 N_15 VDD mp15  l=0.13u w=0.69u m=1
M17 Y N_3 N_15 VDD mp15  l=0.13u w=0.595u m=1
M18 Y N_3 N_15 VDD mp15  l=0.13u w=0.595u m=1
M19 Y N_3 N_15 VDD mp15  l=0.13u w=0.595u m=1
M20 N_15 N_3 Y VDD mp15  l=0.13u w=0.595u m=1
M21 Y N_3 N_15 VDD mp15  l=0.13u w=0.46u m=1
.ends buftd2
* SPICE INPUT		Tue Jul 31 18:56:52 2018	buftd20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd20
.subckt buftd20 GND Y VDD E A
M1 N_5 N_2 GND GND mn15  l=0.13u w=0.47u m=1
M2 N_5 N_2 GND GND mn15  l=0.13u w=0.47u m=1
M3 GND N_2 N_5 GND mn15  l=0.13u w=0.47u m=1
M4 N_5 N_2 GND GND mn15  l=0.13u w=0.47u m=1
M5 GND E N_2 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M8 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M9 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M10 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M11 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M12 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M13 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M14 N_5 E N_16 GND mn15  l=0.13u w=0.56u m=1
M15 N_5 E N_16 GND mn15  l=0.13u w=0.56u m=1
M16 N_5 E N_16 GND mn15  l=0.13u w=0.56u m=1
M17 N_16 E N_5 GND mn15  l=0.13u w=0.32u m=1
M18 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M19 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M20 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M21 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M22 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M23 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M24 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M25 Y N_5 GND GND mn15  l=0.13u w=0.39u m=1
M26 Y N_5 GND GND mn15  l=0.13u w=0.39u m=1
M27 Y N_5 GND GND mn15  l=0.13u w=0.27u m=1
M28 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M29 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M30 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M31 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M32 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M33 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M34 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M35 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M36 Y N_5 GND GND mn15  l=0.13u w=0.39u m=1
M37 Y N_5 GND GND mn15  l=0.13u w=0.39u m=1
M38 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M39 N_2 E VDD VDD mp15  l=0.13u w=0.69u m=1
M40 N_16 E VDD VDD mp15  l=0.13u w=0.69u m=1
M41 N_16 E VDD VDD mp15  l=0.13u w=0.69u m=1
M42 VDD E N_16 VDD mp15  l=0.13u w=0.69u m=1
M43 N_16 E VDD VDD mp15  l=0.13u w=0.69u m=1
M44 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M45 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M46 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M47 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M48 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M49 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M50 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M51 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M52 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.575u m=1
M53 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.575u m=1
M54 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.575u m=1
M55 N_16 N_2 N_5 VDD mp15  l=0.13u w=0.575u m=1
M56 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.57u m=1
M57 N_16 N_2 N_5 VDD mp15  l=0.13u w=0.57u m=1
M58 N_5 N_2 N_16 VDD mp15  l=0.13u w=0.42u m=1
M59 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M60 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M61 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M62 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M63 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M64 Y N_16 VDD VDD mp15  l=0.13u w=0.64u m=1
M65 Y N_16 VDD VDD mp15  l=0.13u w=0.64u m=1
M66 VDD N_16 Y VDD mp15  l=0.13u w=0.64u m=1
M67 Y N_16 VDD VDD mp15  l=0.13u w=0.64u m=1
M68 VDD N_16 Y VDD mp15  l=0.13u w=0.62u m=1
M69 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M70 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M71 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M72 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M73 Y N_16 VDD VDD mp15  l=0.13u w=0.7u m=1
M74 VDD N_16 Y VDD mp15  l=0.13u w=0.7u m=1
M75 Y N_16 VDD VDD mp15  l=0.13u w=0.6u m=1
M76 VDD N_16 Y VDD mp15  l=0.13u w=0.57u m=1
M77 Y N_16 VDD VDD mp15  l=0.13u w=0.57u m=1
M78 VDD N_16 Y VDD mp15  l=0.13u w=0.57u m=1
M79 Y N_16 VDD VDD mp15  l=0.13u w=0.57u m=1
.ends buftd20
* SPICE INPUT		Tue Jul 31 18:57:04 2018	buftd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd3
.subckt buftd3 GND Y VDD E A
M1 N_5 E GND GND mn15  l=0.13u w=0.3u m=1
M2 N_2 A GND GND mn15  l=0.13u w=0.28u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.27u m=1
M4 GND N_5 N_2 GND mn15  l=0.13u w=0.28u m=1
M5 N_3 E N_2 GND mn15  l=0.13u w=0.3u m=1
M6 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M8 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M9 N_5 E VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_3 A VDD VDD mp15  l=0.13u w=0.83u m=1
M11 N_3 N_5 N_2 VDD mp15  l=0.13u w=0.6u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD E N_3 VDD mp15  l=0.13u w=0.41u m=1
.ends buftd3
* SPICE INPUT		Tue Jul 31 18:57:15 2018	buftd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd4
.subckt buftd4 GND Y VDD E A
M1 N_4 E GND GND mn15  l=0.13u w=0.3u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.37u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.37u m=1
M4 N_6 N_4 GND GND mn15  l=0.13u w=0.37u m=1
M5 N_6 E N_2 GND mn15  l=0.13u w=0.39u m=1
M6 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_4 E VDD VDD mp15  l=0.13u w=0.4u m=1
M11 VDD A N_2 VDD mp15  l=0.13u w=0.55u m=1
M12 N_2 A VDD VDD mp15  l=0.13u w=0.55u m=1
M13 VDD E N_2 VDD mp15  l=0.13u w=0.55u m=1
M14 N_6 N_4 N_2 VDD mp15  l=0.13u w=0.64u m=1
M15 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buftd4
* SPICE INPUT		Tue Jul 31 18:57:27 2018	buftd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd6
.subckt buftd6 GND Y VDD A E
M1 GND E N_4 GND mn15  l=0.13u w=0.3u m=1
M2 GND A N_3 GND mn15  l=0.13u w=0.37u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.37u m=1
M4 N_3 A GND GND mn15  l=0.13u w=0.37u m=1
M5 N_3 E N_2 GND mn15  l=0.13u w=0.59u m=1
M6 N_3 N_4 GND GND mn15  l=0.13u w=0.55u m=1
M7 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M13 VDD E N_4 VDD mp15  l=0.13u w=0.42u m=1
M14 N_2 A VDD VDD mp15  l=0.13u w=0.66u m=1
M15 N_2 A VDD VDD mp15  l=0.13u w=0.57u m=1
M16 N_2 A VDD VDD mp15  l=0.13u w=0.45u m=1
M17 N_2 E VDD VDD mp15  l=0.13u w=0.41u m=1
M18 VDD E N_2 VDD mp15  l=0.13u w=0.41u m=1
M19 N_2 N_4 N_3 VDD mp15  l=0.13u w=0.59u m=1
M20 N_3 N_4 N_2 VDD mp15  l=0.13u w=0.57u m=1
M21 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buftd6
* SPICE INPUT		Tue Jul 31 18:57:39 2018	buftd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftd8
.subckt buftd8 GND Y VDD E A
M1 N_4 E GND GND mn15  l=0.13u w=0.4u m=1
M2 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_8 E N_2 GND mn15  l=0.13u w=0.42u m=1
M6 N_2 E N_8 GND mn15  l=0.13u w=0.38u m=1
M7 GND N_4 N_2 GND mn15  l=0.13u w=0.35u m=1
M8 GND N_4 N_2 GND mn15  l=0.13u w=0.35u m=1
M9 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M10 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M16 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD E N_4 VDD mp15  l=0.13u w=0.3u m=1
M18 N_4 E VDD VDD mp15  l=0.13u w=0.3u m=1
M19 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_8 E VDD VDD mp15  l=0.13u w=0.595u m=1
M23 VDD E N_8 VDD mp15  l=0.13u w=0.445u m=1
M24 N_2 N_4 N_8 VDD mp15  l=0.13u w=0.81u m=1
M25 N_2 N_4 N_8 VDD mp15  l=0.13u w=0.75u m=1
M26 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M27 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M29 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M31 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M33 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends buftd8
* SPICE INPUT		Tue Jul 31 18:57:51 2018	buftdm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=buftdm
.subckt buftdm VDD Y GND E A
M1 GND A N_5 GND mn15  l=0.13u w=0.26u m=1
M2 N_31 N_5 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_32 N_5 GND GND mn15  l=0.13u w=0.24u m=1
M4 N_31 E Y GND mn15  l=0.13u w=0.46u m=1
M5 N_32 E Y GND mn15  l=0.13u w=0.24u m=1
M6 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M7 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_7 N_5 VDD VDD mp15  l=0.13u w=0.53u m=1
M9 N_8 N_3 Y VDD mp15  l=0.13u w=0.53u m=1
M10 Y N_3 N_7 VDD mp15  l=0.13u w=0.53u m=1
M11 N_8 N_5 VDD VDD mp15  l=0.13u w=0.53u m=1
M12 N_3 E VDD VDD mp15  l=0.13u w=0.4u m=1
.ends buftdm
* SPICE INPUT		Tue Jul 31 18:58:03 2018	ckandd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckandd0
.subckt ckandd0 Y GND VDD A B
M1 GND N_4 Y GND mn15  l=0.13u w=0.2u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.2u m=1
M3 N_5 B N_4 GND mn15  l=0.13u w=0.2u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.5u m=1
M6 N_4 B VDD VDD mp15  l=0.13u w=0.5u m=1
.ends ckandd0
* SPICE INPUT		Tue Jul 31 18:58:15 2018	ckandd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckandd1
.subckt ckandd1 GND Y VDD A B
M1 Y N_4 GND GND mn15  l=0.13u w=0.39u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M3 N_5 B N_4 GND mn15  l=0.13u w=0.26u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.59u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.59u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.6u m=1
M7 N_4 B VDD VDD mp15  l=0.13u w=0.6u m=1
.ends ckandd1
* SPICE INPUT		Tue Jul 31 18:58:27 2018	ckandd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckandd2
.subckt ckandd2 GND Y VDD A B
M1 N_5 A GND GND mn15  l=0.13u w=0.3u m=1
M2 N_5 B N_4 GND mn15  l=0.13u w=0.3u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M5 N_4 B VDD VDD mp15  l=0.13u w=0.69u m=1
M6 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckandd2
* SPICE INPUT		Tue Jul 31 18:58:39 2018	ckandd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckandd4
.subckt ckandd4 Y GND VDD A B
M1 GND A N_9 GND mn15  l=0.13u w=0.33u m=1
M2 Y N_5 GND GND mn15  l=0.13u w=0.265u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.265u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.265u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.265u m=1
M6 GND A N_10 GND mn15  l=0.13u w=0.27u m=1
M7 N_5 B N_10 GND mn15  l=0.13u w=0.3u m=1
M8 N_5 B N_9 GND mn15  l=0.13u w=0.3u m=1
M9 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.865u m=1
M11 Y N_5 VDD VDD mp15  l=0.13u w=0.865u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.79u m=1
M13 Y N_5 VDD VDD mp15  l=0.13u w=0.24u m=1
M14 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M15 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M16 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends ckandd4
* SPICE INPUT		Tue Jul 31 18:58:51 2018	ckbufd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd0
.subckt ckbufd0 VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.2u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd0
* SPICE INPUT		Tue Jul 31 18:59:05 2018	ckbufd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd1
.subckt ckbufd1 GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.4u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
.ends ckbufd1
* SPICE INPUT		Tue Jul 31 18:59:19 2018	ckbufd10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd10
.subckt ckbufd10 GND Y VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M2 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.35u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_4 A VDD VDD mp15  l=0.13u w=0.735u m=1
M11 VDD A N_4 VDD mp15  l=0.13u w=0.72u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.72u m=1
M13 N_4 A VDD VDD mp15  l=0.13u w=0.705u m=1
M14 Y N_4 VDD VDD mp15  l=0.13u w=1.38u m=1
M15 Y N_4 VDD VDD mp15  l=0.13u w=0.795u m=1
M16 VDD N_4 Y VDD mp15  l=0.13u w=0.72u m=1
M17 Y N_4 VDD VDD mp15  l=0.13u w=0.72u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.72u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.72u m=1
M20 VDD N_4 Y VDD mp15  l=0.13u w=0.72u m=1
M21 Y N_4 VDD VDD mp15  l=0.13u w=0.72u m=1
M22 Y N_4 VDD VDD mp15  l=0.13u w=0.71u m=1
.ends ckbufd10
* SPICE INPUT		Tue Jul 31 18:59:34 2018	ckbufd12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd12
.subckt ckbufd12 Y GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M2 GND A N_4 GND mn15  l=0.13u w=0.36u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.35u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M6 Y N_4 GND GND mn15  l=0.13u w=0.41u m=1
M7 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.41u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.41u m=1
M11 Y N_4 GND GND mn15  l=0.13u w=0.41u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.73u m=1
M13 N_4 A VDD VDD mp15  l=0.13u w=0.72u m=1
M14 N_4 A VDD VDD mp15  l=0.13u w=0.72u m=1
M15 N_4 A VDD VDD mp15  l=0.13u w=0.67u m=1
M16 Y N_4 VDD VDD mp15  l=0.13u w=1.23u m=1
M17 Y N_4 VDD VDD mp15  l=0.13u w=0.91u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.71u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
M21 VDD N_4 Y VDD mp15  l=0.13u w=0.695u m=1
M22 Y N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
M23 VDD N_4 Y VDD mp15  l=0.13u w=0.695u m=1
M24 Y N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
M25 VDD N_4 Y VDD mp15  l=0.13u w=0.695u m=1
M26 Y N_4 VDD VDD mp15  l=0.13u w=0.695u m=1
.ends ckbufd12
* SPICE INPUT		Tue Jul 31 18:59:47 2018	ckbufd14
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd14
.subckt ckbufd14 GND Y VDD A
M1 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.44u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M5 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.44u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.43u m=1
M8 Y N_4 GND GND mn15  l=0.13u w=0.43u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.43u m=1
M10 GND A N_4 GND mn15  l=0.13u w=0.44u m=1
M11 N_4 A GND GND mn15  l=0.13u w=0.435u m=1
M12 GND A N_4 GND mn15  l=0.13u w=0.435u m=1
M13 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M14 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M15 Y N_4 VDD VDD mp15  l=0.13u w=0.8u m=1
M16 VDD N_4 Y VDD mp15  l=0.13u w=0.735u m=1
M17 Y N_4 VDD VDD mp15  l=0.13u w=0.735u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.735u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.725u m=1
M20 VDD N_4 Y VDD mp15  l=0.13u w=0.725u m=1
M21 Y N_4 VDD VDD mp15  l=0.13u w=0.725u m=1
M22 VDD N_4 Y VDD mp15  l=0.13u w=0.725u m=1
M23 Y N_4 VDD VDD mp15  l=0.13u w=0.725u m=1
M24 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M25 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M26 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M27 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M28 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M29 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd14
* SPICE INPUT		Tue Jul 31 19:00:03 2018	ckbufd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd16
.subckt ckbufd16 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.405u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.405u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.405u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.405u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 VDD A N_5 VDD mp15  l=0.13u w=0.72u m=1
M15 VDD A N_5 VDD mp15  l=0.13u w=0.72u m=1
M16 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M18 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M21 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M22 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M23 Y N_5 VDD VDD mp15  l=0.13u w=0.785u m=1
M24 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M25 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M26 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M27 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M28 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M29 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M30 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M31 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M32 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
.ends ckbufd16
* SPICE INPUT		Tue Jul 31 19:00:16 2018	ckbufd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd2
.subckt ckbufd2 GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd2
* SPICE INPUT		Tue Jul 31 19:00:27 2018	ckbufd20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd20
.subckt ckbufd20 GND Y VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M10 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M16 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M18 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M21 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M23 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M25 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M26 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M27 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M28 Y N_5 VDD VDD mp15  l=0.13u w=0.83u m=1
M29 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M30 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M31 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
M32 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M33 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
M34 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M35 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
M36 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M37 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
M38 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
M39 Y N_5 VDD VDD mp15  l=0.13u w=0.705u m=1
.ends ckbufd20
* SPICE INPUT		Tue Jul 31 19:00:39 2018	ckbufd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd3
.subckt ckbufd3 GND Y VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.2u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M5 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd3
* SPICE INPUT		Tue Jul 31 19:00:51 2018	ckbufd30
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd30
.subckt ckbufd30 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.41u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.41u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.41u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.41u m=1
M5 GND A N_5 GND mn15  l=0.13u w=0.41u m=1
M6 N_5 A GND GND mn15  l=0.13u w=0.41u m=1
M7 GND A N_5 GND mn15  l=0.13u w=0.41u m=1
M8 N_5 A GND GND mn15  l=0.13u w=0.41u m=1
M9 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M10 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M11 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M12 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M13 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M14 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M15 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M16 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M17 Y N_5 GND GND mn15  l=0.13u w=0.44u m=1
M18 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M19 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M20 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M21 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M22 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M23 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M24 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M25 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M26 Y N_5 GND GND mn15  l=0.13u w=0.445u m=1
M27 GND N_5 Y GND mn15  l=0.13u w=0.445u m=1
M28 N_5 A VDD VDD mp15  l=0.13u w=0.71u m=1
M29 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M30 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M31 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M32 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M33 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M34 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M35 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M36 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M37 VDD A N_5 VDD mp15  l=0.13u w=0.7u m=1
M38 N_5 A VDD VDD mp15  l=0.13u w=0.7u m=1
M39 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M40 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M41 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M42 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M43 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M44 Y N_5 VDD VDD mp15  l=0.13u w=1.38u m=1
M45 VDD N_5 Y VDD mp15  l=0.13u w=1.38u m=1
M46 Y N_5 VDD VDD mp15  l=0.13u w=0.875u m=1
M47 VDD N_5 Y VDD mp15  l=0.13u w=0.725u m=1
M48 Y N_5 VDD VDD mp15  l=0.13u w=0.725u m=1
M49 VDD N_5 Y VDD mp15  l=0.13u w=0.725u m=1
M50 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M51 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M52 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M53 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M54 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M55 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M56 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M57 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M58 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M59 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M60 VDD N_5 Y VDD mp15  l=0.13u w=0.71u m=1
M61 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M62 Y N_5 VDD VDD mp15  l=0.13u w=0.71u m=1
M63 VDD N_5 Y VDD mp15  l=0.13u w=0.705u m=1
.ends ckbufd30
* SPICE INPUT		Tue Jul 31 19:01:03 2018	ckbufd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd4
.subckt ckbufd4 Y GND VDD A
M1 GND A N_5 GND mn15  l=0.13u w=0.26u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.23u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.27u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.27u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.27u m=1
M6 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_5 A VDD VDD mp15  l=0.13u w=0.71u m=1
M8 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_5 Y VDD mp15  l=0.13u w=0.7u m=1
M10 VDD N_5 Y VDD mp15  l=0.13u w=0.7u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.7u m=1
M12 Y N_5 VDD VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd4
* SPICE INPUT		Tue Jul 31 19:01:15 2018	ckbufd40
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd40
.subckt ckbufd40 GND Y VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M2 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M3 N_4 A GND GND mn15  l=0.13u w=0.43u m=1
M4 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M5 N_4 A GND GND mn15  l=0.13u w=0.43u m=1
M6 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M7 N_4 A GND GND mn15  l=0.13u w=0.43u m=1
M8 GND A N_4 GND mn15  l=0.13u w=0.43u m=1
M9 GND A N_4 GND mn15  l=0.13u w=0.4u m=1
M10 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M11 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M12 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M13 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M14 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M15 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M16 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M17 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M18 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M19 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M20 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M21 Y N_4 GND GND mn15  l=0.13u w=0.44u m=1
M22 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M23 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M24 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M25 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M26 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M27 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M28 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M29 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M30 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M31 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M32 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M33 GND N_4 Y GND mn15  l=0.13u w=0.45u m=1
M34 Y N_4 GND GND mn15  l=0.13u w=0.45u m=1
M35 N_4 A VDD VDD mp15  l=0.13u w=0.71u m=1
M36 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M37 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M38 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M39 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M40 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M41 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M42 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M43 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M44 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M45 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M46 VDD A N_4 VDD mp15  l=0.13u w=0.7u m=1
M47 N_4 A VDD VDD mp15  l=0.13u w=0.7u m=1
M48 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M49 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M50 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M51 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M52 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M53 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M54 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M55 VDD N_4 Y VDD mp15  l=0.13u w=1.37u m=1
M56 Y N_4 VDD VDD mp15  l=0.13u w=1.37u m=1
M57 VDD N_4 Y VDD mp15  l=0.13u w=1.28u m=1
M58 VDD N_4 Y VDD mp15  l=0.13u w=0.705u m=1
M59 Y N_4 VDD VDD mp15  l=0.13u w=0.705u m=1
M60 VDD N_4 Y VDD mp15  l=0.13u w=0.705u m=1
M61 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M62 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M63 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M64 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M65 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M66 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M67 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M68 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M69 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M70 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M71 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M72 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M73 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M74 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M75 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M76 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M77 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M78 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
M79 VDD N_4 Y VDD mp15  l=0.13u w=0.7u m=1
M80 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd40
* SPICE INPUT		Tue Jul 31 19:01:27 2018	ckbufd5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd5
.subckt ckbufd5 GND Y VDD A
M1 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.26u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.27u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.27u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.27u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.27u m=1
M7 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M8 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
M9 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd5
* SPICE INPUT		Tue Jul 31 19:01:39 2018	ckbufd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd6
.subckt ckbufd6 Y GND VDD A
M1 GND A N_4 GND mn15  l=0.13u w=0.44u m=1
M2 GND A N_4 GND mn15  l=0.13u w=0.32u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.27u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.27u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.27u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.27u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.27u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.27u m=1
M9 VDD A N_4 VDD mp15  l=0.13u w=0.72u m=1
M10 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_4 VDD VDD mp15  l=0.13u w=0.88u m=1
M13 Y N_4 VDD VDD mp15  l=0.13u w=0.88u m=1
M14 VDD N_4 Y VDD mp15  l=0.13u w=0.88u m=1
M15 Y N_4 VDD VDD mp15  l=0.13u w=0.88u m=1
M16 Y N_4 VDD VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd6
* SPICE INPUT		Tue Jul 31 19:01:51 2018	ckbufd7
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd7
.subckt ckbufd7 GND Y VDD A
M1 N_6 A GND GND mn15  l=0.13u w=0.39u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.39u m=1
M3 Y N_6 GND GND mn15  l=0.13u w=0.27u m=1
M4 GND N_6 Y GND mn15  l=0.13u w=0.26u m=1
M5 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M6 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M7 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M8 GND N_6 Y GND mn15  l=0.13u w=0.26u m=1
M9 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M10 VDD A N_6 VDD mp15  l=0.13u w=0.705u m=1
M11 N_6 A VDD VDD mp15  l=0.13u w=0.705u m=1
M12 VDD A N_6 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.89u m=1
M14 VDD N_6 Y VDD mp15  l=0.13u w=0.89u m=1
M15 Y N_6 VDD VDD mp15  l=0.13u w=0.89u m=1
M16 VDD N_6 Y VDD mp15  l=0.13u w=0.775u m=1
M17 Y N_6 VDD VDD mp15  l=0.13u w=0.775u m=1
M18 VDD N_6 Y VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd7
* SPICE INPUT		Tue Jul 31 19:02:03 2018	ckbufd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd8
.subckt ckbufd8 Y GND VDD A
M1 N_6 A GND GND mn15  l=0.13u w=0.39u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.39u m=1
M3 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M4 Y N_6 GND GND mn15  l=0.13u w=0.27u m=1
M5 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M6 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M7 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M8 Y N_6 GND GND mn15  l=0.13u w=0.27u m=1
M9 GND N_6 Y GND mn15  l=0.13u w=0.27u m=1
M10 Y N_6 GND GND mn15  l=0.13u w=0.27u m=1
M11 VDD A N_6 VDD mp15  l=0.13u w=0.755u m=1
M12 N_6 A VDD VDD mp15  l=0.13u w=0.7u m=1
M13 VDD A N_6 VDD mp15  l=0.13u w=0.7u m=1
M14 Y N_6 VDD VDD mp15  l=0.13u w=0.825u m=1
M15 VDD N_6 Y VDD mp15  l=0.13u w=0.895u m=1
M16 VDD N_6 Y VDD mp15  l=0.13u w=0.895u m=1
M17 Y N_6 VDD VDD mp15  l=0.13u w=0.895u m=1
M18 VDD N_6 Y VDD mp15  l=0.13u w=0.775u m=1
M19 Y N_6 VDD VDD mp15  l=0.13u w=0.775u m=1
M20 Y N_6 VDD VDD mp15  l=0.13u w=0.7u m=1
.ends ckbufd8
* SPICE INPUT		Tue Jul 31 19:02:16 2018	ckbufd80
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufd80
.subckt ckbufd80 GND Y VDD A
M1 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M2 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M3 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M4 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M5 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M6 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M7 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M8 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M9 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M10 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M12 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M13 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M14 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M15 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M16 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M17 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M18 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M19 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M20 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M21 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M22 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M23 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M24 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M25 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M26 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M27 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M28 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M29 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M30 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M31 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M32 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M33 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M34 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M35 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M36 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M37 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M38 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M39 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M40 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M41 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M42 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M43 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M44 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M45 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M46 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M47 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M48 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M49 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M50 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M51 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M52 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M53 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M54 Y N_2 GND GND mn15  l=0.13u w=0.45u m=1
M55 GND N_2 Y GND mn15  l=0.13u w=0.45u m=1
M56 Y N_2 GND GND mn15  l=0.13u w=0.44u m=1
M57 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M58 N_2 A GND GND mn15  l=0.13u w=0.45u m=1
M59 GND A N_2 GND mn15  l=0.13u w=0.45u m=1
M60 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M61 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M62 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M63 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M64 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M65 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M66 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M67 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M68 N_2 A GND GND mn15  l=0.13u w=0.44u m=1
M69 GND A N_2 GND mn15  l=0.13u w=0.44u m=1
M70 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M71 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M72 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M73 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M74 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M75 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M76 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M77 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M78 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M79 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M80 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M81 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M82 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M83 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M84 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M85 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M86 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M87 VDD N_2 Y VDD mp15  l=0.13u w=1.28u m=1
M88 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M89 Y N_2 VDD VDD mp15  l=0.13u w=1.37u m=1
M90 VDD N_2 Y VDD mp15  l=0.13u w=1.37u m=1
M91 Y N_2 VDD VDD mp15  l=0.13u w=0.715u m=1
M92 VDD N_2 Y VDD mp15  l=0.13u w=0.715u m=1
M93 VDD N_2 Y VDD mp15  l=0.13u w=0.715u m=1
M94 VDD N_2 Y VDD mp15  l=0.13u w=0.71u m=1
M95 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M96 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M97 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M98 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M99 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M100 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M101 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M102 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M103 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M104 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M105 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M106 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M107 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M108 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M109 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M110 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M111 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M112 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M113 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M114 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M115 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M116 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M117 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M118 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M119 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M120 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M121 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M122 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M123 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M124 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M125 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M126 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M127 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M128 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M129 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M130 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M131 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M132 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M133 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M134 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M135 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M136 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M137 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M138 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M139 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M140 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M141 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M142 VDD N_2 Y VDD mp15  l=0.13u w=0.7u m=1
M143 Y N_2 VDD VDD mp15  l=0.13u w=0.7u m=1
M144 VDD A N_2 VDD mp15  l=0.13u w=0.71u m=1
M145 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M146 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M147 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M148 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M149 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M150 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M151 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M152 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M153 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M154 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M155 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M156 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M157 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M158 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M159 VDD A N_2 VDD mp15  l=0.13u w=0.7u m=1
M160 N_2 A VDD VDD mp15  l=0.13u w=0.7u m=1
M161 N_2 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckbufd80
* SPICE INPUT		Tue Jul 31 19:02:31 2018	ckbufdm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckbufdm
.subckt ckbufdm GND Y VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.3u m=1
M3 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
M5 VDD N_4 Y VDD mp15  l=0.13u w=0.37u m=1
.ends ckbufdm
* SPICE INPUT		Tue Jul 31 19:02:46 2018	ckinvd0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd0
.subckt ckinvd0 GND VDD Y A
M1 GND A Y GND mn15  l=0.13u w=0.2u m=1
M2 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd0
* SPICE INPUT		Tue Jul 31 19:03:00 2018	ckinvd1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd1
.subckt ckinvd1 Y VDD GND A
M1 Y A GND GND mn15  l=0.13u w=0.4u m=1
M2 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
.ends ckinvd1
* SPICE INPUT		Tue Jul 31 19:03:15 2018	ckinvd10
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd10
.subckt ckinvd10 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.3u m=1
M2 Y A GND GND mn15  l=0.13u w=0.3u m=1
M3 Y A GND GND mn15  l=0.13u w=0.3u m=1
M4 Y A GND GND mn15  l=0.13u w=0.295u m=1
M5 Y A GND GND mn15  l=0.13u w=0.295u m=1
M6 Y A GND GND mn15  l=0.13u w=0.295u m=1
M7 Y A GND GND mn15  l=0.13u w=0.295u m=1
M8 Y A GND GND mn15  l=0.13u w=0.295u m=1
M9 GND A Y GND mn15  l=0.13u w=0.295u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.805u m=1
M11 Y A VDD VDD mp15  l=0.13u w=0.805u m=1
M12 VDD A Y VDD mp15  l=0.13u w=0.805u m=1
M13 Y A VDD VDD mp15  l=0.13u w=0.805u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.805u m=1
M15 Y A VDD VDD mp15  l=0.13u w=0.805u m=1
M16 VDD A Y VDD mp15  l=0.13u w=0.805u m=1
M17 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 Y A VDD VDD mp15  l=0.13u w=0.685u m=1
.ends ckinvd10
* SPICE INPUT		Tue Jul 31 19:03:31 2018	ckinvd12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd12
.subckt ckinvd12 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.3u m=1
M2 Y A GND GND mn15  l=0.13u w=0.295u m=1
M3 Y A GND GND mn15  l=0.13u w=0.295u m=1
M4 Y A GND GND mn15  l=0.13u w=0.295u m=1
M5 GND A Y GND mn15  l=0.13u w=0.295u m=1
M6 Y A GND GND mn15  l=0.13u w=0.295u m=1
M7 GND A Y GND mn15  l=0.13u w=0.295u m=1
M8 Y A GND GND mn15  l=0.13u w=0.295u m=1
M9 GND A Y GND mn15  l=0.13u w=0.295u m=1
M10 Y A GND GND mn15  l=0.13u w=0.295u m=1
M11 GND A Y GND mn15  l=0.13u w=0.295u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.79u m=1
M13 Y A VDD VDD mp15  l=0.13u w=0.79u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M15 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M16 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M17 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M18 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M19 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M20 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M21 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd12
* SPICE INPUT		Tue Jul 31 19:03:43 2018	ckinvd14
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd14
.subckt ckinvd14 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.345u m=1
M2 GND A Y GND mn15  l=0.13u w=0.315u m=1
M3 Y A GND GND mn15  l=0.13u w=0.315u m=1
M4 Y A GND GND mn15  l=0.13u w=0.315u m=1
M5 Y A GND GND mn15  l=0.13u w=0.315u m=1
M6 Y A GND GND mn15  l=0.13u w=0.315u m=1
M7 Y A GND GND mn15  l=0.13u w=0.315u m=1
M8 Y A GND GND mn15  l=0.13u w=0.315u m=1
M9 Y A GND GND mn15  l=0.13u w=0.315u m=1
M10 Y A GND GND mn15  l=0.13u w=0.315u m=1
M11 Y A GND GND mn15  l=0.13u w=0.315u m=1
M12 Y A GND GND mn15  l=0.13u w=0.315u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M15 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M16 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M17 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M18 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M19 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M20 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M21 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M22 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M23 Y A VDD VDD mp15  l=0.13u w=0.782u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd14
* SPICE INPUT		Tue Jul 31 19:03:55 2018	ckinvd16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd16
.subckt ckinvd16 Y GND VDD A
M1 Y A GND GND mn15  l=0.13u w=0.315u m=1
M2 Y A GND GND mn15  l=0.13u w=0.315u m=1
M3 Y A GND GND mn15  l=0.13u w=0.315u m=1
M4 Y A GND GND mn15  l=0.13u w=0.315u m=1
M5 GND A Y GND mn15  l=0.13u w=0.31u m=1
M6 GND A Y GND mn15  l=0.13u w=0.31u m=1
M7 GND A Y GND mn15  l=0.13u w=0.31u m=1
M8 Y A GND GND mn15  l=0.13u w=0.31u m=1
M9 GND A Y GND mn15  l=0.13u w=0.31u m=1
M10 Y A GND GND mn15  l=0.13u w=0.31u m=1
M11 GND A Y GND mn15  l=0.13u w=0.31u m=1
M12 Y A GND GND mn15  l=0.13u w=0.31u m=1
M13 GND A Y GND mn15  l=0.13u w=0.31u m=1
M14 Y A GND GND mn15  l=0.13u w=0.31u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M16 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M17 Y A VDD VDD mp15  l=0.13u w=0.825u m=1
M18 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M19 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M20 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M21 Y A VDD VDD mp15  l=0.13u w=0.82u m=1
M22 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M23 Y A VDD VDD mp15  l=0.13u w=0.82u m=1
M24 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M25 Y A VDD VDD mp15  l=0.13u w=0.82u m=1
M26 VDD A Y VDD mp15  l=0.13u w=0.82u m=1
M27 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd16
* SPICE INPUT		Tue Jul 31 19:04:07 2018	ckinvd2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd2
.subckt ckinvd2 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.26u m=1
M2 Y A GND GND mn15  l=0.13u w=0.23u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M4 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd2
* SPICE INPUT		Tue Jul 31 19:04:18 2018	ckinvd20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd20
.subckt ckinvd20 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.31u m=1
M2 GND A Y GND mn15  l=0.13u w=0.31u m=1
M3 GND A Y GND mn15  l=0.13u w=0.31u m=1
M4 Y A GND GND mn15  l=0.13u w=0.31u m=1
M5 GND A Y GND mn15  l=0.13u w=0.31u m=1
M6 Y A GND GND mn15  l=0.13u w=0.31u m=1
M7 GND A Y GND mn15  l=0.13u w=0.31u m=1
M8 Y A GND GND mn15  l=0.13u w=0.31u m=1
M9 GND A Y GND mn15  l=0.13u w=0.31u m=1
M10 Y A GND GND mn15  l=0.13u w=0.31u m=1
M11 GND A Y GND mn15  l=0.13u w=0.31u m=1
M12 Y A GND GND mn15  l=0.13u w=0.31u m=1
M13 GND A Y GND mn15  l=0.13u w=0.31u m=1
M14 Y A GND GND mn15  l=0.13u w=0.31u m=1
M15 GND A Y GND mn15  l=0.13u w=0.31u m=1
M16 Y A GND GND mn15  l=0.13u w=0.31u m=1
M17 GND A Y GND mn15  l=0.13u w=0.31u m=1
M18 Y A GND GND mn15  l=0.13u w=0.31u m=1
M19 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M20 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M21 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M23 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M25 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M26 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M27 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M29 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M30 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M31 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M32 Y A VDD VDD mp15  l=0.13u w=0.75u m=1
M33 VDD A Y VDD mp15  l=0.13u w=0.75u m=1
M34 Y A VDD VDD mp15  l=0.13u w=0.7u m=1
M35 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M36 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M37 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd20
* SPICE INPUT		Tue Jul 31 19:04:30 2018	ckinvd3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd3
.subckt ckinvd3 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M5 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd3
* SPICE INPUT		Tue Jul 31 19:04:42 2018	ckinvd30
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd30
.subckt ckinvd30 Y GND VDD A
M1 Y A GND GND mn15  l=0.13u w=0.325u m=1
M2 Y A GND GND mn15  l=0.13u w=0.325u m=1
M3 GND A Y GND mn15  l=0.13u w=0.325u m=1
M4 Y A GND GND mn15  l=0.13u w=0.325u m=1
M5 GND A Y GND mn15  l=0.13u w=0.325u m=1
M6 Y A GND GND mn15  l=0.13u w=0.325u m=1
M7 GND A Y GND mn15  l=0.13u w=0.325u m=1
M8 Y A GND GND mn15  l=0.13u w=0.325u m=1
M9 GND A Y GND mn15  l=0.13u w=0.325u m=1
M10 Y A GND GND mn15  l=0.13u w=0.325u m=1
M11 GND A Y GND mn15  l=0.13u w=0.325u m=1
M12 Y A GND GND mn15  l=0.13u w=0.325u m=1
M13 GND A Y GND mn15  l=0.13u w=0.32u m=1
M14 Y A GND GND mn15  l=0.13u w=0.32u m=1
M15 GND A Y GND mn15  l=0.13u w=0.32u m=1
M16 GND A Y GND mn15  l=0.13u w=0.32u m=1
M17 GND A Y GND mn15  l=0.13u w=0.32u m=1
M18 Y A GND GND mn15  l=0.13u w=0.32u m=1
M19 GND A Y GND mn15  l=0.13u w=0.32u m=1
M20 Y A GND GND mn15  l=0.13u w=0.32u m=1
M21 GND A Y GND mn15  l=0.13u w=0.32u m=1
M22 Y A GND GND mn15  l=0.13u w=0.32u m=1
M23 GND A Y GND mn15  l=0.13u w=0.32u m=1
M24 Y A GND GND mn15  l=0.13u w=0.32u m=1
M25 GND A Y GND mn15  l=0.13u w=0.32u m=1
M26 Y A GND GND mn15  l=0.13u w=0.32u m=1
M27 Y A VDD VDD mp15  l=0.13u w=0.83u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.83u m=1
M29 VDD A Y VDD mp15  l=0.13u w=0.83u m=1
M30 Y A VDD VDD mp15  l=0.13u w=0.83u m=1
M31 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M32 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M33 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M34 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M35 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M36 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M37 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M38 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M39 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M40 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M41 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M42 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M43 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M44 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M45 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M46 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M47 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M48 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M49 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M50 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M51 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M52 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M53 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd30
* SPICE INPUT		Tue Jul 31 19:04:55 2018	ckinvd4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd4
.subckt ckinvd4 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.29u m=1
M2 GND A Y GND mn15  l=0.13u w=0.26u m=1
M3 GND A Y GND mn15  l=0.13u w=0.26u m=1
M4 GND A Y GND mn15  l=0.13u w=0.26u m=1
M5 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M6 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd4
* SPICE INPUT		Tue Jul 31 19:05:07 2018	ckinvd40
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd40
.subckt ckinvd40 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.32u m=1
M2 GND A Y GND mn15  l=0.13u w=0.32u m=1
M3 Y A GND GND mn15  l=0.13u w=0.32u m=1
M4 GND A Y GND mn15  l=0.13u w=0.32u m=1
M5 Y A GND GND mn15  l=0.13u w=0.32u m=1
M6 GND A Y GND mn15  l=0.13u w=0.32u m=1
M7 Y A GND GND mn15  l=0.13u w=0.32u m=1
M8 GND A Y GND mn15  l=0.13u w=0.32u m=1
M9 Y A GND GND mn15  l=0.13u w=0.32u m=1
M10 Y A GND GND mn15  l=0.13u w=0.32u m=1
M11 GND A Y GND mn15  l=0.13u w=0.32u m=1
M12 Y A GND GND mn15  l=0.13u w=0.32u m=1
M13 GND A Y GND mn15  l=0.13u w=0.32u m=1
M14 Y A GND GND mn15  l=0.13u w=0.32u m=1
M15 GND A Y GND mn15  l=0.13u w=0.32u m=1
M16 Y A GND GND mn15  l=0.13u w=0.32u m=1
M17 GND A Y GND mn15  l=0.13u w=0.32u m=1
M18 GND A Y GND mn15  l=0.13u w=0.32u m=1
M19 Y A GND GND mn15  l=0.13u w=0.32u m=1
M20 GND A Y GND mn15  l=0.13u w=0.32u m=1
M21 Y A GND GND mn15  l=0.13u w=0.32u m=1
M22 GND A Y GND mn15  l=0.13u w=0.32u m=1
M23 Y A GND GND mn15  l=0.13u w=0.32u m=1
M24 GND A Y GND mn15  l=0.13u w=0.32u m=1
M25 Y A GND GND mn15  l=0.13u w=0.32u m=1
M26 Y A GND GND mn15  l=0.13u w=0.315u m=1
M27 Y A GND GND mn15  l=0.13u w=0.315u m=1
M28 Y A GND GND mn15  l=0.13u w=0.315u m=1
M29 GND A Y GND mn15  l=0.13u w=0.315u m=1
M30 Y A GND GND mn15  l=0.13u w=0.315u m=1
M31 GND A Y GND mn15  l=0.13u w=0.315u m=1
M32 GND A Y GND mn15  l=0.13u w=0.32u m=1
M33 GND A Y GND mn15  l=0.13u w=0.32u m=1
M34 Y A GND GND mn15  l=0.13u w=0.32u m=1
M35 GND A Y GND mn15  l=0.13u w=0.32u m=1
M36 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M37 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M38 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M39 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M40 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M41 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M42 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M43 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M44 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M45 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M46 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M47 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M48 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M49 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M50 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M51 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M52 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M53 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M54 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M55 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M56 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M57 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M58 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M59 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M60 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M61 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M62 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M63 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M64 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M65 Y A VDD VDD mp15  l=0.13u w=0.825u m=1
M66 VDD A Y VDD mp15  l=0.13u w=0.825u m=1
M67 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M68 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M69 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M70 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M71 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd40
* SPICE INPUT		Tue Jul 31 19:05:20 2018	ckinvd5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd5
.subckt ckinvd5 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.3u m=1
M2 Y A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y A GND GND mn15  l=0.13u w=0.26u m=1
M5 GND A Y GND mn15  l=0.13u w=0.26u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd5
* SPICE INPUT		Tue Jul 31 19:05:35 2018	ckinvd6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd6
.subckt ckinvd6 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.27u m=1
M2 GND A Y GND mn15  l=0.13u w=0.27u m=1
M3 GND A Y GND mn15  l=0.13u w=0.27u m=1
M4 Y A GND GND mn15  l=0.13u w=0.27u m=1
M5 GND A Y GND mn15  l=0.13u w=0.27u m=1
M6 Y A GND GND mn15  l=0.13u w=0.27u m=1
M7 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd6
* SPICE INPUT		Tue Jul 31 19:05:49 2018	ckinvd7
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd7
.subckt ckinvd7 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.28u m=1
M2 Y A GND GND mn15  l=0.13u w=0.27u m=1
M3 Y A GND GND mn15  l=0.13u w=0.27u m=1
M4 Y A GND GND mn15  l=0.13u w=0.27u m=1
M5 GND A Y GND mn15  l=0.13u w=0.27u m=1
M6 Y A GND GND mn15  l=0.13u w=0.27u m=1
M7 GND A Y GND mn15  l=0.13u w=0.27u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd7
* SPICE INPUT		Tue Jul 31 19:06:02 2018	ckinvd8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd8
.subckt ckinvd8 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.3u m=1
M2 GND A Y GND mn15  l=0.13u w=0.3u m=1
M3 Y A GND GND mn15  l=0.13u w=0.3u m=1
M4 GND A Y GND mn15  l=0.13u w=0.3u m=1
M5 Y A GND GND mn15  l=0.13u w=0.3u m=1
M6 Y A GND GND mn15  l=0.13u w=0.295u m=1
M7 Y A GND GND mn15  l=0.13u w=0.295u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.85u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.85u m=1
M10 VDD A Y VDD mp15  l=0.13u w=0.85u m=1
M11 Y A VDD VDD mp15  l=0.13u w=0.845u m=1
M12 VDD A Y VDD mp15  l=0.13u w=0.845u m=1
M13 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckinvd8
* SPICE INPUT		Tue Jul 31 19:06:17 2018	ckinvd80
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvd80
.subckt ckinvd80 GND Y VDD A
M1 GND A Y GND mn15  l=0.13u w=0.315u m=1
M2 Y A GND GND mn15  l=0.13u w=0.315u m=1
M3 GND A Y GND mn15  l=0.13u w=0.315u m=1
M4 Y A GND GND mn15  l=0.13u w=0.315u m=1
M5 GND A Y GND mn15  l=0.13u w=0.315u m=1
M6 Y A GND GND mn15  l=0.13u w=0.315u m=1
M7 GND A Y GND mn15  l=0.13u w=0.315u m=1
M8 Y A GND GND mn15  l=0.13u w=0.315u m=1
M9 GND A Y GND mn15  l=0.13u w=0.315u m=1
M10 GND A Y GND mn15  l=0.13u w=0.315u m=1
M11 GND A Y GND mn15  l=0.13u w=0.27u m=1
M12 Y A GND GND mn15  l=0.13u w=0.27u m=1
M13 GND A Y GND mn15  l=0.13u w=0.27u m=1
M14 Y A GND GND mn15  l=0.13u w=0.27u m=1
M15 GND A Y GND mn15  l=0.13u w=0.275u m=1
M16 Y A GND GND mn15  l=0.13u w=0.315u m=1
M17 GND A Y GND mn15  l=0.13u w=0.315u m=1
M18 Y A GND GND mn15  l=0.13u w=0.315u m=1
M19 Y A GND GND mn15  l=0.13u w=0.315u m=1
M20 GND A Y GND mn15  l=0.13u w=0.325u m=1
M21 GND A Y GND mn15  l=0.13u w=0.325u m=1
M22 Y A GND GND mn15  l=0.13u w=0.325u m=1
M23 Y A GND GND mn15  l=0.13u w=0.325u m=1
M24 GND A Y GND mn15  l=0.13u w=0.325u m=1
M25 Y A GND GND mn15  l=0.13u w=0.325u m=1
M26 GND A Y GND mn15  l=0.13u w=0.325u m=1
M27 Y A GND GND mn15  l=0.13u w=0.325u m=1
M28 GND A Y GND mn15  l=0.13u w=0.325u m=1
M29 Y A GND GND mn15  l=0.13u w=0.325u m=1
M30 GND A Y GND mn15  l=0.13u w=0.325u m=1
M31 GND A Y GND mn15  l=0.13u w=0.325u m=1
M32 GND A Y GND mn15  l=0.13u w=0.325u m=1
M33 Y A GND GND mn15  l=0.13u w=0.325u m=1
M34 GND A Y GND mn15  l=0.13u w=0.325u m=1
M35 Y A GND GND mn15  l=0.13u w=0.325u m=1
M36 GND A Y GND mn15  l=0.13u w=0.325u m=1
M37 Y A GND GND mn15  l=0.13u w=0.325u m=1
M38 Y A GND GND mn15  l=0.13u w=0.325u m=1
M39 Y A GND GND mn15  l=0.13u w=0.325u m=1
M40 GND A Y GND mn15  l=0.13u w=0.325u m=1
M41 Y A GND GND mn15  l=0.13u w=0.325u m=1
M42 Y A GND GND mn15  l=0.13u w=0.325u m=1
M43 Y A GND GND mn15  l=0.13u w=0.325u m=1
M44 GND A Y GND mn15  l=0.13u w=0.325u m=1
M45 Y A GND GND mn15  l=0.13u w=0.325u m=1
M46 GND A Y GND mn15  l=0.13u w=0.325u m=1
M47 Y A GND GND mn15  l=0.13u w=0.325u m=1
M48 GND A Y GND mn15  l=0.13u w=0.325u m=1
M49 Y A GND GND mn15  l=0.13u w=0.325u m=1
M50 Y A GND GND mn15  l=0.13u w=0.325u m=1
M51 GND A Y GND mn15  l=0.13u w=0.325u m=1
M52 Y A GND GND mn15  l=0.13u w=0.325u m=1
M53 GND A Y GND mn15  l=0.13u w=0.325u m=1
M54 Y A GND GND mn15  l=0.13u w=0.325u m=1
M55 GND A Y GND mn15  l=0.13u w=0.325u m=1
M56 Y A GND GND mn15  l=0.13u w=0.325u m=1
M57 Y A GND GND mn15  l=0.13u w=0.325u m=1
M58 GND A Y GND mn15  l=0.13u w=0.325u m=1
M59 Y A GND GND mn15  l=0.13u w=0.325u m=1
M60 GND A Y GND mn15  l=0.13u w=0.325u m=1
M61 Y A GND GND mn15  l=0.13u w=0.325u m=1
M62 GND A Y GND mn15  l=0.13u w=0.325u m=1
M63 Y A GND GND mn15  l=0.13u w=0.325u m=1
M64 GND A Y GND mn15  l=0.13u w=0.325u m=1
M65 Y A GND GND mn15  l=0.13u w=0.325u m=1
M66 GND A Y GND mn15  l=0.13u w=0.325u m=1
M67 Y A GND GND mn15  l=0.13u w=0.325u m=1
M68 GND A Y GND mn15  l=0.13u w=0.325u m=1
M69 Y A GND GND mn15  l=0.13u w=0.325u m=1
M70 GND A Y GND mn15  l=0.13u w=0.325u m=1
M71 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M72 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M73 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M74 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M75 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M76 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M77 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M78 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M79 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M80 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M81 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M82 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M83 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M84 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M85 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M86 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M87 VDD A Y VDD mp15  l=0.13u w=0.835u m=1
M88 Y A VDD VDD mp15  l=0.13u w=0.835u m=1
M89 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M90 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M91 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M92 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M93 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M94 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M95 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M96 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M97 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M98 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M99 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M100 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M101 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M102 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M103 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M104 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M105 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M106 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M107 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M108 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M109 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M110 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M111 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M112 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M113 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M114 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M115 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M116 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M117 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M118 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M119 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M120 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M121 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M122 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M123 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M124 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M125 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M126 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M127 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M128 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M129 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M130 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M131 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M132 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M133 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M134 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M135 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M136 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M137 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M138 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M139 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
M140 Y A VDD VDD mp15  l=0.13u w=0.78u m=1
M141 VDD A Y VDD mp15  l=0.13u w=0.78u m=1
.ends ckinvd80
* SPICE INPUT		Tue Jul 31 19:06:32 2018	ckinvdm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckinvdm
.subckt ckinvdm Y VDD GND A
M1 Y A GND GND mn15  l=0.13u w=0.3u m=1
M2 VDD A Y VDD mp15  l=0.13u w=0.49u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.49u m=1
.ends ckinvdm
* SPICE INPUT		Tue Jul 31 19:06:44 2018	ckmx02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckmx02d0
.subckt ckmx02d0 VDD Y GND S0 B A
M1 N_16 B GND GND mn15  l=0.13u w=0.19u m=1
M2 GND S0 N_3 GND mn15  l=0.13u w=0.18u m=1
M3 N_15 N_3 N_6 GND mn15  l=0.13u w=0.19u m=1
M4 N_15 A GND GND mn15  l=0.13u w=0.19u m=1
M5 GND N_6 Y GND mn15  l=0.13u w=0.19u m=1
M6 N_16 S0 N_6 GND mn15  l=0.13u w=0.19u m=1
M7 N_8 B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_8 N_3 N_6 VDD mp15  l=0.13u w=0.69u m=1
M9 N_3 S0 VDD VDD mp15  l=0.13u w=0.26u m=1
M10 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M12 N_6 S0 N_7 VDD mp15  l=0.13u w=0.69u m=1
.ends ckmx02d0
* SPICE INPUT		Tue Jul 31 19:06:55 2018	ckmx02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckmx02d1
.subckt ckmx02d1 VDD Y GND S0 B A
M1 N_16 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_7 GND GND mn15  l=0.13u w=0.39u m=1
M3 GND S0 N_2 GND mn15  l=0.13u w=0.18u m=1
M4 N_17 B GND GND mn15  l=0.13u w=0.2u m=1
M5 N_7 N_2 N_16 GND mn15  l=0.13u w=0.2u m=1
M6 N_17 S0 N_7 GND mn15  l=0.13u w=0.2u m=1
M7 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_7 Y VDD mp15  l=0.13u w=0.59u m=1
M9 Y N_7 VDD VDD mp15  l=0.13u w=0.59u m=1
M10 VDD S0 N_2 VDD mp15  l=0.13u w=0.24u m=1
M11 N_9 B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_9 N_2 N_7 VDD mp15  l=0.13u w=0.69u m=1
M13 N_7 S0 N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends ckmx02d1
* SPICE INPUT		Tue Jul 31 19:07:07 2018	ckmx02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckmx02d2
.subckt ckmx02d2 GND Y VDD S0 B A
M1 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.19u m=1
M3 N_3 S0 GND GND mn15  l=0.13u w=0.32u m=1
M4 N_8 S0 N_6 GND mn15  l=0.13u w=0.32u m=1
M5 N_8 B GND GND mn15  l=0.13u w=0.18u m=1
M6 N_7 N_3 N_6 GND mn15  l=0.13u w=0.32u m=1
M7 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_3 S0 VDD VDD mp15  l=0.13u w=0.46u m=1
M11 N_6 S0 N_7 VDD mp15  l=0.13u w=0.5u m=1
M12 N_8 B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_8 N_3 N_6 VDD mp15  l=0.13u w=0.5u m=1
.ends ckmx02d2
* SPICE INPUT		Tue Jul 31 19:07:19 2018	ckmx02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckmx02d4
.subckt ckmx02d4 GND Y A B S0 VDD
M1 N_5 S0 N_4 GND mn15  l=0.13u w=0.45u m=1
M2 N_3 S0 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_5 B GND GND mn15  l=0.13u w=0.155u m=1
M4 GND B N_5 GND mn15  l=0.13u w=0.155u m=1
M5 N_5 B GND GND mn15  l=0.13u w=0.15u m=1
M6 N_9 N_3 N_4 GND mn15  l=0.13u w=0.45u m=1
M7 GND A N_9 GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.3u m=1
M10 Y N_4 GND GND mn15  l=0.13u w=0.29u m=1
M11 VDD S0 N_3 VDD mp15  l=0.13u w=0.42u m=1
M12 N_9 S0 N_4 VDD mp15  l=0.13u w=0.67u m=1
M13 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_5 B VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_5 N_3 N_4 VDD mp15  l=0.13u w=0.64u m=1
M16 N_9 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_9 VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckmx02d4
* SPICE INPUT		Tue Jul 31 19:07:31 2018	cknd02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknd02d0
.subckt cknd02d0 Y VDD A GND B
M1 GND A N_14 GND mn15  l=0.13u w=0.27u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.27u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.6u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.6u m=1
.ends cknd02d0
* SPICE INPUT		Tue Jul 31 19:07:43 2018	cknd02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknd02d1
.subckt cknd02d1 Y VDD A B GND
M1 GND A N_9 GND mn15  l=0.13u w=0.36u m=1
M2 Y B N_9 GND mn15  l=0.13u w=0.36u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
.ends cknd02d1
* SPICE INPUT		Tue Jul 31 19:07:56 2018	cknd02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknd02d2
.subckt cknd02d2 GND Y VDD A B
M1 N_6 A GND GND mn15  l=0.13u w=0.43u m=1
M2 N_6 B Y GND mn15  l=0.13u w=0.43u m=1
M3 Y B N_5 GND mn15  l=0.13u w=0.42u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.42u m=1
M5 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends cknd02d2
* SPICE INPUT		Tue Jul 31 19:08:08 2018	cknd02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknd02d4
.subckt cknd02d4 Y GND A B VDD
M1 Y B N_7 GND mn15  l=0.13u w=0.4u m=1
M2 GND A N_7 GND mn15  l=0.13u w=0.4u m=1
M3 N_10 A GND GND mn15  l=0.13u w=0.4u m=1
M4 N_10 B Y GND mn15  l=0.13u w=0.4u m=1
M5 Y B N_9 GND mn15  l=0.13u w=0.4u m=1
M6 N_8 A GND GND mn15  l=0.13u w=0.4u m=1
M7 N_9 A GND GND mn15  l=0.13u w=0.4u m=1
M8 N_8 B Y GND mn15  l=0.13u w=0.4u m=1
M9 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
.ends cknd02d4
* SPICE INPUT		Tue Jul 31 19:08:21 2018	cknr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknr02d0
.subckt cknr02d0 GND Y VDD B A
M1 GND A Y GND mn15  l=0.13u w=0.18u m=1
M2 Y B GND GND mn15  l=0.13u w=0.18u m=1
M3 N_10 A VDD VDD mp15  l=0.13u w=0.6u m=1
M4 N_11 A VDD VDD mp15  l=0.13u w=0.6u m=1
M5 Y B N_10 VDD mp15  l=0.13u w=0.6u m=1
M6 Y B N_11 VDD mp15  l=0.13u w=0.6u m=1
.ends cknr02d0
* SPICE INPUT		Tue Jul 31 19:08:36 2018	cknr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknr02d1
.subckt cknr02d1 GND Y VDD B A
M1 Y B GND GND mn15  l=0.13u w=0.23u m=1
M2 GND A Y GND mn15  l=0.13u w=0.23u m=1
M3 N_10 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 Y B N_10 VDD mp15  l=0.13u w=0.69u m=1
M5 Y B N_11 VDD mp15  l=0.13u w=0.69u m=1
M6 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends cknr02d1
* SPICE INPUT		Tue Jul 31 19:08:51 2018	cknr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknr02d2
.subckt cknr02d2 Y GND VDD B A
M1 GND B Y GND mn15  l=0.13u w=0.4u m=1
M2 GND A Y GND mn15  l=0.13u w=0.4u m=1
M3 N_9 A VDD VDD mp15  l=0.13u w=0.69u m=1
M4 N_10 B Y VDD mp15  l=0.13u w=0.69u m=1
M5 Y B N_9 VDD mp15  l=0.13u w=0.69u m=1
M6 VDD A N_8 VDD mp15  l=0.13u w=0.69u m=1
M7 N_10 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y B N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends cknr02d2
* SPICE INPUT		Tue Jul 31 19:09:04 2018	cknr02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=cknr02d4
.subckt cknr02d4 Y GND VDD A B
M1 GND A Y GND mn15  l=0.13u w=0.3u m=1
M2 GND A Y GND mn15  l=0.13u w=0.3u m=1
M3 GND B Y GND mn15  l=0.13u w=0.3u m=1
M4 GND B Y GND mn15  l=0.13u w=0.3u m=1
M5 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 N_17 B Y VDD mp15  l=0.13u w=0.69u m=1
M7 Y B N_16 VDD mp15  l=0.13u w=0.69u m=1
M8 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y B N_15 VDD mp15  l=0.13u w=0.69u m=1
M11 Y B N_18 VDD mp15  l=0.13u w=0.69u m=1
M12 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends cknr02d4
* SPICE INPUT		Tue Jul 31 19:09:21 2018	ckor02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckor02d0
.subckt ckor02d0 GND Y B VDD A
M1 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.26u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M5 N_19 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M6 N_19 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckor02d0
* SPICE INPUT		Tue Jul 31 19:09:34 2018	ckor02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckor02d1
.subckt ckor02d1 GND Y VDD A B
M1 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M3 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_13 A VDD VDD mp15  l=0.13u w=0.68u m=1
M5 N_13 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M6 N_3 B N_12 VDD mp15  l=0.13u w=0.68u m=1
M7 N_12 A VDD VDD mp15  l=0.13u w=0.68u m=1
M8 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckor02d1
* SPICE INPUT		Tue Jul 31 19:09:45 2018	ckor02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckor02d2
.subckt ckor02d2 GND Y VDD A B
M1 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M7 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_43 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M10 N_3 B N_42 VDD mp15  l=0.13u w=0.68u m=1
M11 N_43 A VDD VDD mp15  l=0.13u w=0.68u m=1
M12 N_40 A VDD VDD mp15  l=0.13u w=0.68u m=1
M13 N_41 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M14 N_3 B N_40 VDD mp15  l=0.13u w=0.68u m=1
M15 N_42 A VDD VDD mp15  l=0.13u w=0.68u m=1
M16 VDD A N_41 VDD mp15  l=0.13u w=0.68u m=1
.ends ckor02d2
* SPICE INPUT		Tue Jul 31 19:09:57 2018	ckor02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckor02d4
.subckt ckor02d4 GND Y A B VDD
M1 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND B N_3 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_60 A VDD VDD mp15  l=0.13u w=0.68u m=1
M12 N_61 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M13 N_3 B N_60 VDD mp15  l=0.13u w=0.68u m=1
M14 N_62 A VDD VDD mp15  l=0.13u w=0.68u m=1
M15 VDD A N_61 VDD mp15  l=0.13u w=0.68u m=1
M16 N_63 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M17 N_3 B N_62 VDD mp15  l=0.13u w=0.68u m=1
M18 N_64 A VDD VDD mp15  l=0.13u w=0.68u m=1
M19 VDD A N_63 VDD mp15  l=0.13u w=0.68u m=1
M20 N_65 B N_3 VDD mp15  l=0.13u w=0.68u m=1
M21 N_3 B N_64 VDD mp15  l=0.13u w=0.68u m=1
M22 N_65 A VDD VDD mp15  l=0.13u w=0.68u m=1
M23 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckor02d4
* SPICE INPUT		Tue Jul 31 19:10:09 2018	ckxn02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxn02d0
.subckt ckxn02d0 GND Y VDD A B
M1 GND B N_2 GND mn15  l=0.13u w=0.2u m=1
M2 N_9 N_2 GND GND mn15  l=0.13u w=0.2u m=1
M3 N_9 N_8 N_3 GND mn15  l=0.13u w=0.2u m=1
M4 N_3 A N_2 GND mn15  l=0.13u w=0.2u m=1
M5 GND N_3 Y GND mn15  l=0.13u w=0.2u m=1
M6 N_8 A GND GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M8 N_16 N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_16 A N_3 VDD mp15  l=0.13u w=0.69u m=1
M10 N_2 N_8 N_3 VDD mp15  l=0.13u w=0.345u m=1
M11 N_2 N_8 N_3 VDD mp15  l=0.13u w=0.345u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckxn02d0
* SPICE INPUT		Tue Jul 31 19:10:20 2018	ckxn02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxn02d1
.subckt ckxn02d1 GND Y VDD A B
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_6 GND GND mn15  l=0.13u w=0.4u m=1
M3 N_6 A N_5 GND mn15  l=0.13u w=0.2u m=1
M4 GND B N_5 GND mn15  l=0.13u w=0.2u m=1
M5 N_9 N_5 GND GND mn15  l=0.13u w=0.2u m=1
M6 N_9 N_4 N_6 GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_38 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_38 A N_6 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.35u m=1
M11 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.34u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.59u m=1
M14 VDD N_6 Y VDD mp15  l=0.13u w=0.59u m=1
.ends ckxn02d1
* SPICE INPUT		Tue Jul 31 19:10:32 2018	ckxn02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxn02d2
.subckt ckxn02d2 GND Y VDD A B
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_6 A N_5 GND mn15  l=0.13u w=0.2u m=1
M4 GND B N_5 GND mn15  l=0.13u w=0.2u m=1
M5 N_9 N_5 GND GND mn15  l=0.13u w=0.2u m=1
M6 N_9 N_4 N_6 GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_38 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_38 A N_6 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.35u m=1
M11 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.34u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckxn02d2
* SPICE INPUT		Tue Jul 31 19:10:44 2018	ckxn02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxn02d4
.subckt ckxn02d4 GND Y VDD B A
M1 N_3 N_6 N_2 GND mn15  l=0.13u w=0.39u m=1
M2 N_6 A GND GND mn15  l=0.13u w=0.18u m=1
M3 N_2 N_8 GND GND mn15  l=0.13u w=0.39u m=1
M4 N_8 A N_3 GND mn15  l=0.13u w=0.39u m=1
M5 N_8 B GND GND mn15  l=0.13u w=0.39u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.355u m=1
M7 Y N_3 GND GND mn15  l=0.13u w=0.355u m=1
M8 Y N_3 GND GND mn15  l=0.13u w=0.35u m=1
M9 N_8 N_6 N_3 VDD mp15  l=0.13u w=0.59u m=1
M10 N_3 N_6 N_8 VDD mp15  l=0.13u w=0.59u m=1
M11 N_20 A N_3 VDD mp15  l=0.13u w=0.59u m=1
M12 N_3 A N_19 VDD mp15  l=0.13u w=0.59u m=1
M13 N_6 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_8 B VDD VDD mp15  l=0.13u w=0.59u m=1
M15 N_8 B VDD VDD mp15  l=0.13u w=0.59u m=1
M16 N_19 N_8 VDD VDD mp15  l=0.13u w=0.59u m=1
M17 N_20 N_8 VDD VDD mp15  l=0.13u w=0.59u m=1
M18 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M21 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckxn02d4
* SPICE INPUT		Tue Jul 31 19:10:57 2018	ckxr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxr02d0
.subckt ckxr02d0 GND Y A VDD B
M1 GND B N_2 GND mn15  l=0.13u w=0.2u m=1
M2 N_9 N_2 GND GND mn15  l=0.13u w=0.2u m=1
M3 N_3 N_8 N_2 GND mn15  l=0.13u w=0.2u m=1
M4 N_9 A N_3 GND mn15  l=0.13u w=0.2u m=1
M5 N_8 A GND GND mn15  l=0.13u w=0.2u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M8 N_37 N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_37 N_8 N_3 VDD mp15  l=0.13u w=0.69u m=1
M10 N_2 A N_3 VDD mp15  l=0.13u w=0.345u m=1
M11 N_3 A N_2 VDD mp15  l=0.13u w=0.345u m=1
M12 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckxr02d0
* SPICE INPUT		Tue Jul 31 19:11:08 2018	ckxr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxr02d1
.subckt ckxr02d1 GND Y A VDD B
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_8 GND GND mn15  l=0.13u w=0.4u m=1
M3 GND B N_5 GND mn15  l=0.13u w=0.2u m=1
M4 N_9 N_5 GND GND mn15  l=0.13u w=0.2u m=1
M5 N_8 N_4 N_5 GND mn15  l=0.13u w=0.2u m=1
M6 N_8 A N_9 GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_16 N_4 N_8 VDD mp15  l=0.13u w=0.69u m=1
M9 N_16 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_8 A N_5 VDD mp15  l=0.13u w=0.345u m=1
M11 N_5 A N_8 VDD mp15  l=0.13u w=0.345u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_8 Y VDD mp15  l=0.13u w=0.61u m=1
M14 VDD N_8 Y VDD mp15  l=0.13u w=0.61u m=1
.ends ckxr02d1
* SPICE INPUT		Tue Jul 31 19:11:22 2018	ckxr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxr02d2
.subckt ckxr02d2 GND Y A VDD B
M1 N_4 A GND GND mn15  l=0.13u w=0.2u m=1
M2 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_5 GND mn15  l=0.13u w=0.2u m=1
M4 N_9 N_5 GND GND mn15  l=0.13u w=0.2u m=1
M5 N_8 N_4 N_5 GND mn15  l=0.13u w=0.2u m=1
M6 N_8 A N_9 GND mn15  l=0.13u w=0.2u m=1
M7 VDD B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_16 N_4 N_8 VDD mp15  l=0.13u w=0.69u m=1
M9 N_16 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_8 A N_5 VDD mp15  l=0.13u w=0.345u m=1
M11 N_5 A N_8 VDD mp15  l=0.13u w=0.345u m=1
M12 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ckxr02d2
* SPICE INPUT		Tue Jul 31 19:11:37 2018	ckxr02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ckxr02d4
.subckt ckxr02d4 GND Y VDD A B
M1 N_3 B GND GND mn15  l=0.13u w=0.39u m=1
M2 N_11 N_3 GND GND mn15  l=0.13u w=0.39u m=1
M3 N_11 A N_2 GND mn15  l=0.13u w=0.39u m=1
M4 N_3 N_8 N_2 GND mn15  l=0.13u w=0.39u m=1
M5 GND A N_8 GND mn15  l=0.13u w=0.19u m=1
M6 Y N_2 GND GND mn15  l=0.13u w=0.355u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.355u m=1
M8 Y N_2 GND GND mn15  l=0.13u w=0.35u m=1
M9 VDD B N_3 VDD mp15  l=0.13u w=0.59u m=1
M10 N_3 B VDD VDD mp15  l=0.13u w=0.59u m=1
M11 N_16 N_3 VDD VDD mp15  l=0.13u w=0.59u m=1
M12 VDD N_3 N_16 VDD mp15  l=0.13u w=0.59u m=1
M13 N_16 N_8 N_2 VDD mp15  l=0.13u w=0.59u m=1
M14 N_16 N_8 N_2 VDD mp15  l=0.13u w=0.59u m=1
M15 N_2 A N_3 VDD mp15  l=0.13u w=1.18u m=1
M16 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ckxr02d4
* SPICE INPUT		Tue Jul 31 19:11:52 2018	denrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=denrq0
.subckt denrq0 VDD Q GND CK D E
M1 N_33 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_6 E N_33 GND mn15  l=0.13u w=0.18u m=1
M3 GND E N_5 GND mn15  l=0.13u w=0.18u m=1
M4 N_34 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M5 N_34 N_17 GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.17u m=1
M7 N_12 N_2 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_35 N_12 N_9 GND mn15  l=0.13u w=0.17u m=1
M9 GND N_8 N_35 GND mn15  l=0.13u w=0.17u m=1
M10 N_8 N_9 GND GND mn15  l=0.13u w=0.18u m=1
M11 Q N_16 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_17 N_16 GND GND mn15  l=0.13u w=0.18u m=1
M13 N_9 N_2 N_6 GND mn15  l=0.13u w=0.28u m=1
M14 N_37 N_2 N_16 GND mn15  l=0.13u w=0.17u m=1
M15 N_36 N_8 GND GND mn15  l=0.13u w=0.17u m=1
M16 N_16 N_12 N_36 GND mn15  l=0.13u w=0.17u m=1
M17 N_37 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M18 N_18 D VDD VDD mp15  l=0.13u w=0.28u m=1
M19 N_5 E VDD VDD mp15  l=0.13u w=0.26u m=1
M20 N_6 E N_19 VDD mp15  l=0.13u w=0.28u m=1
M21 N_6 N_5 N_18 VDD mp15  l=0.13u w=0.28u m=1
M22 N_19 N_17 VDD VDD mp15  l=0.13u w=0.28u m=1
M23 VDD CK N_2 VDD mp15  l=0.13u w=0.42u m=1
M24 N_6 N_12 N_9 VDD mp15  l=0.13u w=0.42u m=1
M25 N_20 N_8 VDD VDD mp15  l=0.13u w=0.17u m=1
M26 N_8 N_9 VDD VDD mp15  l=0.13u w=0.26u m=1
M27 N_20 N_2 N_9 VDD mp15  l=0.13u w=0.17u m=1
M28 N_12 N_2 VDD VDD mp15  l=0.13u w=0.42u m=1
M29 Q N_16 VDD VDD mp15  l=0.13u w=0.4u m=1
M30 N_17 N_16 VDD VDD mp15  l=0.13u w=0.26u m=1
M31 N_21 N_2 N_16 VDD mp15  l=0.13u w=0.27u m=1
M32 N_21 N_8 VDD VDD mp15  l=0.13u w=0.27u m=1
M33 N_22 N_12 N_16 VDD mp15  l=0.13u w=0.17u m=1
M34 N_22 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
.ends denrq0
* SPICE INPUT		Tue Jul 31 19:12:05 2018	denrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=denrq1
.subckt denrq1 VDD Q GND CK E D
M1 N_35 D GND GND mn15  l=0.13u w=0.28u m=1
M2 N_6 E N_35 GND mn15  l=0.13u w=0.28u m=1
M3 GND E N_4 GND mn15  l=0.13u w=0.17u m=1
M4 N_36 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_36 N_18 GND GND mn15  l=0.13u w=0.28u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_37 N_15 N_9 GND mn15  l=0.13u w=0.17u m=1
M8 N_37 N_8 GND GND mn15  l=0.13u w=0.17u m=1
M9 GND N_9 N_8 GND mn15  l=0.13u w=0.28u m=1
M10 N_6 N_2 N_9 GND mn15  l=0.13u w=0.28u m=1
M11 N_12 N_15 N_38 GND mn15  l=0.13u w=0.36u m=1
M12 N_38 N_8 GND GND mn15  l=0.13u w=0.36u m=1
M13 GND N_18 N_39 GND mn15  l=0.13u w=0.17u m=1
M14 N_39 N_2 N_12 GND mn15  l=0.13u w=0.17u m=1
M15 GND N_2 N_15 GND mn15  l=0.13u w=0.2u m=1
M16 Q N_12 GND GND mn15  l=0.13u w=0.46u m=1
M17 N_18 N_12 GND GND mn15  l=0.13u w=0.28u m=1
M18 N_24 D VDD VDD mp15  l=0.13u w=0.42u m=1
M19 VDD E N_4 VDD mp15  l=0.13u w=0.24u m=1
M20 N_24 N_4 N_6 VDD mp15  l=0.13u w=0.42u m=1
M21 N_25 E N_6 VDD mp15  l=0.13u w=0.42u m=1
M22 N_25 N_18 VDD VDD mp15  l=0.13u w=0.42u m=1
M23 VDD CK N_2 VDD mp15  l=0.13u w=0.51u m=1
M24 N_6 N_15 N_9 VDD mp15  l=0.13u w=0.42u m=1
M25 N_26 N_8 VDD VDD mp15  l=0.13u w=0.17u m=1
M26 N_8 N_9 VDD VDD mp15  l=0.13u w=0.26u m=1
M27 VDD N_9 N_8 VDD mp15  l=0.13u w=0.16u m=1
M28 N_26 N_2 N_9 VDD mp15  l=0.13u w=0.17u m=1
M29 N_27 N_15 N_12 VDD mp15  l=0.13u w=0.17u m=1
M30 VDD N_18 N_27 VDD mp15  l=0.13u w=0.17u m=1
M31 N_28 N_2 N_12 VDD mp15  l=0.13u w=0.52u m=1
M32 VDD N_8 N_28 VDD mp15  l=0.13u w=0.52u m=1
M33 N_15 N_2 VDD VDD mp15  l=0.13u w=0.51u m=1
M34 Q N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 N_18 N_12 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends denrq1
* SPICE INPUT		Tue Jul 31 19:12:21 2018	denrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=denrq2
.subckt denrq2 Q GND D E CK VDD
M1 GND N_12 Q GND mn15  l=0.13u w=0.46u m=1
M2 GND N_12 Q GND mn15  l=0.13u w=0.46u m=1
M3 GND N_12 N_4 GND mn15  l=0.13u w=0.37u m=1
M4 GND CK N_6 GND mn15  l=0.13u w=0.27u m=1
M5 N_22 N_4 GND GND mn15  l=0.13u w=0.28u m=1
M6 N_22 N_8 N_10 GND mn15  l=0.13u w=0.28u m=1
M7 N_10 E N_21 GND mn15  l=0.13u w=0.28u m=1
M8 GND E N_8 GND mn15  l=0.13u w=0.24u m=1
M9 N_21 D GND GND mn15  l=0.13u w=0.28u m=1
M10 N_23 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_12 N_6 N_23 GND mn15  l=0.13u w=0.17u m=1
M12 N_14 N_6 GND GND mn15  l=0.13u w=0.22u m=1
M13 GND N_17 N_24 GND mn15  l=0.13u w=0.41u m=1
M14 N_12 N_14 N_24 GND mn15  l=0.13u w=0.41u m=1
M15 N_10 N_6 N_19 GND mn15  l=0.13u w=0.41u m=1
M16 GND N_19 N_17 GND mn15  l=0.13u w=0.41u m=1
M17 N_25 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M18 N_25 N_14 N_19 GND mn15  l=0.13u w=0.17u m=1
M19 VDD N_12 Q VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_12 Q VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_12 N_4 VDD mp15  l=0.13u w=0.55u m=1
M22 N_96 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M23 N_12 N_14 N_96 VDD mp15  l=0.13u w=0.17u m=1
M24 VDD N_6 N_14 VDD mp15  l=0.13u w=0.55u m=1
M25 N_97 N_17 VDD VDD mp15  l=0.13u w=0.62u m=1
M26 N_97 N_6 N_12 VDD mp15  l=0.13u w=0.62u m=1
M27 N_98 N_6 N_19 VDD mp15  l=0.13u w=0.17u m=1
M28 N_17 N_19 VDD VDD mp15  l=0.13u w=0.315u m=1
M29 VDD N_19 N_17 VDD mp15  l=0.13u w=0.315u m=1
M30 N_98 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M31 N_10 N_14 N_19 VDD mp15  l=0.13u w=0.615u m=1
M32 VDD CK N_6 VDD mp15  l=0.13u w=0.67u m=1
M33 N_100 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M34 N_100 E N_10 VDD mp15  l=0.13u w=0.42u m=1
M35 N_99 N_8 N_10 VDD mp15  l=0.13u w=0.42u m=1
M36 VDD E N_8 VDD mp15  l=0.13u w=0.37u m=1
M37 N_99 D VDD VDD mp15  l=0.13u w=0.42u m=1
.ends denrq2
* SPICE INPUT		Tue Jul 31 19:12:37 2018	dfanrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfanrq0
.subckt dfanrq0 VDD Q GND D1 D0 CK
M1 GND CK N_15 GND mn15  l=0.13u w=0.17u m=1
M2 N_26 D0 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_5 N_15 N_4 GND mn15  l=0.13u w=0.28u m=1
M4 N_27 N_8 N_5 GND mn15  l=0.13u w=0.17u m=1
M5 GND N_2 N_27 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_5 N_2 GND mn15  l=0.13u w=0.18u m=1
M7 N_4 D1 N_26 GND mn15  l=0.13u w=0.26u m=1
M8 GND N_15 N_8 GND mn15  l=0.13u w=0.17u m=1
M9 N_28 N_8 N_10 GND mn15  l=0.13u w=0.17u m=1
M10 N_29 N_11 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_28 N_2 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_29 N_15 N_10 GND mn15  l=0.13u w=0.17u m=1
M13 Q N_10 GND GND mn15  l=0.13u w=0.26u m=1
M14 N_11 N_10 GND GND mn15  l=0.13u w=0.18u m=1
M15 N_5 N_8 N_4 VDD mp15  l=0.13u w=0.42u m=1
M16 N_16 N_2 VDD VDD mp15  l=0.13u w=0.17u m=1
M17 N_16 N_15 N_5 VDD mp15  l=0.13u w=0.17u m=1
M18 VDD N_5 N_2 VDD mp15  l=0.13u w=0.26u m=1
M19 VDD N_15 N_8 VDD mp15  l=0.13u w=0.42u m=1
M20 N_18 N_11 VDD VDD mp15  l=0.13u w=0.17u m=1
M21 N_17 N_2 VDD VDD mp15  l=0.13u w=0.27u m=1
M22 N_10 N_15 N_17 VDD mp15  l=0.13u w=0.27u m=1
M23 N_18 N_8 N_10 VDD mp15  l=0.13u w=0.17u m=1
M24 Q N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M25 N_11 N_10 VDD VDD mp15  l=0.13u w=0.26u m=1
M26 N_15 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M27 VDD D0 N_4 VDD mp15  l=0.13u w=0.35u m=1
M28 N_4 D1 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends dfanrq0
* SPICE INPUT		Tue Jul 31 19:12:49 2018	dfanrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfanrq1
.subckt dfanrq1 GND Q VDD D1 D0 CK
M1 GND CK N_3 GND mn15  l=0.13u w=0.2u m=1
M2 N_15 D0 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_5 D1 N_15 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 N_3 N_5 GND mn15  l=0.13u w=0.28u m=1
M5 GND N_2 N_16 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_6 N_2 GND mn15  l=0.13u w=0.28u m=1
M7 N_16 N_9 N_6 GND mn15  l=0.13u w=0.17u m=1
M8 N_18 N_9 N_11 GND mn15  l=0.13u w=0.37u m=1
M9 N_11 N_3 N_17 GND mn15  l=0.13u w=0.17u m=1
M10 N_17 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_18 N_2 GND GND mn15  l=0.13u w=0.37u m=1
M12 GND N_3 N_9 GND mn15  l=0.13u w=0.2u m=1
M13 Q N_11 GND GND mn15  l=0.13u w=0.46u m=1
M14 N_14 N_11 GND GND mn15  l=0.13u w=0.28u m=1
M15 N_3 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M16 N_5 D0 VDD VDD mp15  l=0.13u w=0.35u m=1
M17 N_5 D1 VDD VDD mp15  l=0.13u w=0.35u m=1
M18 N_30 N_3 N_6 VDD mp15  l=0.13u w=0.17u m=1
M19 N_30 N_2 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 VDD N_6 N_2 VDD mp15  l=0.13u w=0.41u m=1
M21 N_5 N_9 N_6 VDD mp15  l=0.13u w=0.42u m=1
M22 Q N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_14 N_11 VDD VDD mp15  l=0.13u w=0.35u m=1
M24 N_11 N_9 N_31 VDD mp15  l=0.13u w=0.17u m=1
M25 N_32 N_3 N_11 VDD mp15  l=0.13u w=0.54u m=1
M26 N_31 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_32 N_2 VDD VDD mp15  l=0.13u w=0.54u m=1
M28 VDD N_3 N_9 VDD mp15  l=0.13u w=0.51u m=1
.ends dfanrq1
* SPICE INPUT		Tue Jul 31 19:13:02 2018	dfanrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfanrq2
.subckt dfanrq2 GND Q VDD D0 D1 CK
M1 N_5 CK GND GND mn15  l=0.13u w=0.28u m=1
M2 N_16 D1 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_16 D0 N_6 GND mn15  l=0.13u w=0.46u m=1
M4 N_7 N_5 N_6 GND mn15  l=0.13u w=0.41u m=1
M5 GND N_3 N_17 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_7 N_3 GND mn15  l=0.13u w=0.205u m=1
M7 N_3 N_7 GND GND mn15  l=0.13u w=0.205u m=1
M8 N_17 N_11 N_7 GND mn15  l=0.13u w=0.17u m=1
M9 GND N_5 N_11 GND mn15  l=0.13u w=0.22u m=1
M10 N_18 N_3 GND GND mn15  l=0.13u w=0.41u m=1
M11 N_18 N_11 N_13 GND mn15  l=0.13u w=0.41u m=1
M12 N_19 N_5 N_13 GND mn15  l=0.13u w=0.17u m=1
M13 GND N_10 N_19 GND mn15  l=0.13u w=0.17u m=1
M14 Q N_13 GND GND mn15  l=0.13u w=0.46u m=1
M15 Q N_13 GND GND mn15  l=0.13u w=0.46u m=1
M16 N_10 N_13 GND GND mn15  l=0.13u w=0.37u m=1
M17 N_5 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M18 VDD D1 N_6 VDD mp15  l=0.13u w=0.61u m=1
M19 N_6 D0 VDD VDD mp15  l=0.13u w=0.61u m=1
M20 N_31 N_5 N_7 VDD mp15  l=0.13u w=0.17u m=1
M21 N_31 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_3 N_7 VDD VDD mp15  l=0.13u w=0.3u m=1
M23 N_3 N_7 VDD VDD mp15  l=0.13u w=0.33u m=1
M24 N_7 N_11 N_6 VDD mp15  l=0.13u w=0.63u m=1
M25 N_11 N_5 VDD VDD mp15  l=0.13u w=0.55u m=1
M26 N_32 N_3 VDD VDD mp15  l=0.13u w=0.63u m=1
M27 N_33 N_11 N_13 VDD mp15  l=0.13u w=0.17u m=1
M28 N_32 N_5 N_13 VDD mp15  l=0.13u w=0.63u m=1
M29 VDD N_10 N_33 VDD mp15  l=0.13u w=0.17u m=1
M30 Q N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 Q N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 N_10 N_13 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends dfanrq2
* SPICE INPUT		Tue Jul 31 19:13:14 2018	dfbfb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb0
.subckt dfbfb0 GND Q QN VDD RN SN D CKN
M1 GND N_2 N_3 GND mn15  l=0.13u w=0.17u m=1
M2 GND CKN N_2 GND mn15  l=0.13u w=0.18u m=1
M3 N_22 D GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 N_2 N_21 GND mn15  l=0.13u w=0.17u m=1
M5 N_21 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M6 N_22 N_3 N_7 GND mn15  l=0.13u w=0.26u m=1
M7 N_11 N_2 N_9 GND mn15  l=0.13u w=0.28u m=1
M8 N_11 N_3 N_23 GND mn15  l=0.13u w=0.17u m=1
M9 N_23 N_20 N_8 GND mn15  l=0.13u w=0.17u m=1
M10 N_8 N_7 N_9 GND mn15  l=0.13u w=0.28u m=1
M11 N_11 N_17 N_8 GND mn15  l=0.13u w=0.2u m=1
M12 N_8 SN GND GND mn15  l=0.13u w=0.36u m=1
M13 N_17 RN GND GND mn15  l=0.13u w=0.18u m=1
M14 Q N_20 GND GND mn15  l=0.13u w=0.26u m=1
M15 QN N_11 GND GND mn15  l=0.13u w=0.26u m=1
M16 N_20 N_11 GND GND mn15  l=0.13u w=0.18u m=1
M17 N_3 N_2 VDD VDD mp15  l=0.13u w=0.42u m=1
M18 N_2 CKN VDD VDD mp15  l=0.13u w=0.46u m=1
M19 N_90 D VDD VDD mp15  l=0.13u w=0.38u m=1
M20 N_90 N_2 N_7 VDD mp15  l=0.13u w=0.38u m=1
M21 N_89 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_7 N_3 N_89 VDD mp15  l=0.13u w=0.17u m=1
M23 N_11 N_2 N_32 VDD mp15  l=0.13u w=0.17u m=1
M24 N_11 N_3 N_9 VDD mp15  l=0.13u w=0.46u m=1
M25 N_9 N_7 N_28 VDD mp15  l=0.13u w=0.45u m=1
M26 N_28 N_20 N_32 VDD mp15  l=0.13u w=0.17u m=1
M27 N_28 N_17 VDD VDD mp15  l=0.13u w=0.595u m=1
M28 VDD SN N_11 VDD mp15  l=0.13u w=0.28u m=1
M29 N_17 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M30 Q N_20 VDD VDD mp15  l=0.13u w=0.4u m=1
M31 QN N_11 VDD VDD mp15  l=0.13u w=0.4u m=1
M32 N_20 N_11 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends dfbfb0
* SPICE INPUT		Tue Jul 31 19:13:26 2018	dfbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb1
.subckt dfbfb1 GND QN Q VDD D SN RN CKN
M1 GND N_2 N_3 GND mn15  l=0.13u w=0.2u m=1
M2 GND CKN N_2 GND mn15  l=0.13u w=0.2u m=1
M3 QN N_14 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_7 N_14 GND GND mn15  l=0.13u w=0.28u m=1
M5 N_10 RN GND GND mn15  l=0.13u w=0.18u m=1
M6 Q N_7 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_23 D GND GND mn15  l=0.13u w=0.28u m=1
M8 N_13 N_2 N_22 GND mn15  l=0.13u w=0.17u m=1
M9 N_22 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M10 N_23 N_3 N_13 GND mn15  l=0.13u w=0.28u m=1
M11 N_16 N_13 N_15 GND mn15  l=0.13u w=0.4u m=1
M12 N_15 N_2 N_14 GND mn15  l=0.13u w=0.36u m=1
M13 N_14 N_3 N_24 GND mn15  l=0.13u w=0.17u m=1
M14 N_24 N_7 N_16 GND mn15  l=0.13u w=0.17u m=1
M15 N_14 N_10 N_16 GND mn15  l=0.13u w=0.28u m=1
M16 N_16 SN GND GND mn15  l=0.13u w=0.46u m=1
M17 N_3 N_2 VDD VDD mp15  l=0.13u w=0.51u m=1
M18 N_2 CKN VDD VDD mp15  l=0.13u w=0.51u m=1
M19 QN N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_7 N_14 VDD VDD mp15  l=0.13u w=0.37u m=1
M21 N_96 D VDD VDD mp15  l=0.13u w=0.42u m=1
M22 N_96 N_2 N_13 VDD mp15  l=0.13u w=0.42u m=1
M23 N_95 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 N_13 N_3 N_95 VDD mp15  l=0.13u w=0.17u m=1
M25 N_15 N_13 N_33 VDD mp15  l=0.13u w=0.295u m=1
M26 N_15 N_13 N_33 VDD mp15  l=0.13u w=0.295u m=1
M27 N_14 N_2 N_34 VDD mp15  l=0.13u w=0.17u m=1
M28 N_15 N_3 N_14 VDD mp15  l=0.13u w=0.56u m=1
M29 N_33 N_10 VDD VDD mp15  l=0.13u w=0.35u m=1
M30 N_33 N_10 VDD VDD mp15  l=0.13u w=0.35u m=1
M31 N_33 N_7 N_34 VDD mp15  l=0.13u w=0.17u m=1
M32 N_14 SN VDD VDD mp15  l=0.13u w=0.36u m=1
M33 N_10 RN VDD VDD mp15  l=0.13u w=0.28u m=1
M34 Q N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends dfbfb1
* SPICE INPUT		Tue Jul 31 19:13:40 2018	dfbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbfb2
.subckt dfbfb2 GND Q QN VDD RN SN D CKN
M1 GND CKN N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_25 D GND GND mn15  l=0.13u w=0.43u m=1
M3 N_25 N_2 N_6 GND mn15  l=0.13u w=0.43u m=1
M4 N_26 N_7 GND GND mn15  l=0.13u w=0.16u m=1
M5 GND N_4 N_2 GND mn15  l=0.13u w=0.22u m=1
M6 N_26 N_4 N_6 GND mn15  l=0.13u w=0.16u m=1
M7 N_9 N_6 N_7 GND mn15  l=0.13u w=0.305u m=1
M8 N_7 N_6 N_9 GND mn15  l=0.13u w=0.305u m=1
M9 N_8 N_4 N_7 GND mn15  l=0.13u w=0.45u m=1
M10 N_27 N_23 N_9 GND mn15  l=0.13u w=0.17u m=1
M11 N_8 N_2 N_27 GND mn15  l=0.13u w=0.17u m=1
M12 N_9 SN GND GND mn15  l=0.13u w=0.29u m=1
M13 GND SN N_9 GND mn15  l=0.13u w=0.29u m=1
M14 GND SN N_9 GND mn15  l=0.13u w=0.3u m=1
M15 N_8 N_19 N_9 GND mn15  l=0.13u w=0.36u m=1
M16 GND RN N_19 GND mn15  l=0.13u w=0.28u m=1
M17 Q N_23 GND GND mn15  l=0.13u w=0.46u m=1
M18 GND N_23 Q GND mn15  l=0.13u w=0.46u m=1
M19 GND N_8 QN GND mn15  l=0.13u w=0.46u m=1
M20 GND N_8 QN GND mn15  l=0.13u w=0.46u m=1
M21 GND N_8 N_23 GND mn15  l=0.13u w=0.36u m=1
M22 N_4 CKN VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_106 D VDD VDD mp15  l=0.13u w=0.64u m=1
M24 N_107 N_2 N_6 VDD mp15  l=0.13u w=0.16u m=1
M25 N_107 N_7 VDD VDD mp15  l=0.13u w=0.16u m=1
M26 VDD N_4 N_2 VDD mp15  l=0.13u w=0.55u m=1
M27 N_106 N_4 N_6 VDD mp15  l=0.13u w=0.64u m=1
M28 N_7 N_6 N_35 VDD mp15  l=0.13u w=0.45u m=1
M29 N_35 N_6 N_7 VDD mp15  l=0.13u w=0.45u m=1
M30 N_7 N_6 N_35 VDD mp15  l=0.13u w=0.44u m=1
M31 N_8 N_4 N_108 VDD mp15  l=0.13u w=0.17u m=1
M32 N_108 N_23 N_35 VDD mp15  l=0.13u w=0.17u m=1
M33 N_8 N_2 N_7 VDD mp15  l=0.13u w=0.56u m=1
M34 N_8 SN VDD VDD mp15  l=0.13u w=0.56u m=1
M35 N_35 N_19 VDD VDD mp15  l=0.13u w=0.45u m=1
M36 N_35 N_19 VDD VDD mp15  l=0.13u w=0.45u m=1
M37 N_35 N_19 VDD VDD mp15  l=0.13u w=0.44u m=1
M38 N_19 RN VDD VDD mp15  l=0.13u w=0.42u m=1
M39 VDD N_23 Q VDD mp15  l=0.13u w=0.69u m=1
M40 Q N_23 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 VDD N_8 QN VDD mp15  l=0.13u w=0.69u m=1
M42 VDD N_8 QN VDD mp15  l=0.13u w=0.69u m=1
M43 VDD N_8 N_23 VDD mp15  l=0.13u w=0.53u m=1
.ends dfbfb2
* SPICE INPUT		Tue Jul 31 19:13:55 2018	dfbrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb0
.subckt dfbrb0 GND Q QN VDD SN RN D CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.18u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_7 N_2 N_21 GND mn15  l=0.13u w=0.17u m=1
M4 N_21 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_22 N_4 N_7 GND mn15  l=0.13u w=0.26u m=1
M6 N_22 D GND GND mn15  l=0.13u w=0.26u m=1
M7 N_8 N_7 N_9 GND mn15  l=0.13u w=0.28u m=1
M8 N_11 N_2 N_9 GND mn15  l=0.13u w=0.28u m=1
M9 N_11 N_4 N_23 GND mn15  l=0.13u w=0.17u m=1
M10 N_23 N_17 N_8 GND mn15  l=0.13u w=0.17u m=1
M11 N_14 RN GND GND mn15  l=0.13u w=0.18u m=1
M12 Q N_17 GND GND mn15  l=0.13u w=0.26u m=1
M13 QN N_11 GND GND mn15  l=0.13u w=0.26u m=1
M14 N_17 N_11 GND GND mn15  l=0.13u w=0.18u m=1
M15 N_11 N_14 N_8 GND mn15  l=0.13u w=0.2u m=1
M16 N_8 SN GND GND mn15  l=0.13u w=0.37u m=1
M17 N_4 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M18 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M19 N_90 N_2 N_7 VDD mp15  l=0.13u w=0.37u m=1
M20 N_89 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M21 N_7 N_4 N_89 VDD mp15  l=0.13u w=0.17u m=1
M22 N_90 D VDD VDD mp15  l=0.13u w=0.37u m=1
M23 N_9 N_7 N_31 VDD mp15  l=0.13u w=0.46u m=1
M24 N_11 N_2 N_32 VDD mp15  l=0.13u w=0.17u m=1
M25 N_11 N_4 N_9 VDD mp15  l=0.13u w=0.46u m=1
M26 N_14 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M27 Q N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 QN N_11 VDD VDD mp15  l=0.13u w=0.4u m=1
M29 N_17 N_11 VDD VDD mp15  l=0.13u w=0.26u m=1
M30 N_31 N_17 N_32 VDD mp15  l=0.13u w=0.17u m=1
M31 N_31 N_14 VDD VDD mp15  l=0.13u w=0.585u m=1
M32 VDD SN N_11 VDD mp15  l=0.13u w=0.28u m=1
.ends dfbrb0
* SPICE INPUT		Tue Jul 31 19:14:08 2018	dfbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb1
.subckt dfbrb1 GND QN Q CK D SN RN VDD
M1 QN N_10 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 N_10 GND GND mn15  l=0.13u w=0.28u m=1
M3 Q N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_7 RN GND GND mn15  l=0.13u w=0.18u m=1
M5 N_9 SN GND GND mn15  l=0.13u w=0.46u m=1
M6 N_10 N_7 N_9 GND mn15  l=0.13u w=0.28u m=1
M7 N_10 N_21 N_22 GND mn15  l=0.13u w=0.17u m=1
M8 N_22 N_4 N_9 GND mn15  l=0.13u w=0.17u m=1
M9 N_9 N_18 N_13 GND mn15  l=0.13u w=0.4u m=1
M10 N_10 N_19 N_13 GND mn15  l=0.13u w=0.4u m=1
M11 N_18 N_19 N_23 GND mn15  l=0.13u w=0.17u m=1
M12 N_23 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M13 N_24 N_21 N_18 GND mn15  l=0.13u w=0.28u m=1
M14 N_24 D GND GND mn15  l=0.13u w=0.28u m=1
M15 GND N_21 N_19 GND mn15  l=0.13u w=0.17u m=1
M16 N_21 CK GND GND mn15  l=0.13u w=0.2u m=1
M17 QN N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_4 N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M19 Q N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_7 RN VDD VDD mp15  l=0.13u w=0.28u m=1
M21 N_10 SN VDD VDD mp15  l=0.13u w=0.37u m=1
M22 N_19 N_21 VDD VDD mp15  l=0.13u w=0.44u m=1
M23 N_21 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M24 N_31 N_4 N_30 VDD mp15  l=0.13u w=0.17u m=1
M25 N_31 N_7 VDD VDD mp15  l=0.13u w=0.35u m=1
M26 N_31 N_7 VDD VDD mp15  l=0.13u w=0.35u m=1
M27 N_13 N_18 N_31 VDD mp15  l=0.13u w=0.345u m=1
M28 N_13 N_18 N_31 VDD mp15  l=0.13u w=0.325u m=1
M29 N_10 N_19 N_30 VDD mp15  l=0.13u w=0.17u m=1
M30 N_13 N_21 N_10 VDD mp15  l=0.13u w=0.55u m=1
M31 N_95 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_18 N_21 N_95 VDD mp15  l=0.13u w=0.17u m=1
M33 N_96 N_19 N_18 VDD mp15  l=0.13u w=0.42u m=1
M34 N_96 D VDD VDD mp15  l=0.13u w=0.42u m=1
.ends dfbrb1
* SPICE INPUT		Tue Jul 31 19:14:22 2018	dfbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrb2
.subckt dfbrb2 GND Q QN RN SN VDD D CK
M1 N_5 CK GND GND mn15  l=0.13u w=0.28u m=1
M2 N_26 D GND GND mn15  l=0.13u w=0.43u m=1
M3 N_27 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M4 N_27 N_2 N_6 GND mn15  l=0.13u w=0.17u m=1
M5 N_26 N_5 N_6 GND mn15  l=0.13u w=0.43u m=1
M6 GND N_5 N_2 GND mn15  l=0.13u w=0.17u m=1
M7 N_28 N_24 N_7 GND mn15  l=0.13u w=0.17u m=1
M8 N_9 N_6 N_7 GND mn15  l=0.13u w=0.21u m=1
M9 N_7 N_6 N_9 GND mn15  l=0.13u w=0.21u m=1
M10 N_9 N_6 N_7 GND mn15  l=0.13u w=0.21u m=1
M11 N_12 N_2 N_9 GND mn15  l=0.13u w=0.42u m=1
M12 N_28 N_5 N_12 GND mn15  l=0.13u w=0.17u m=1
M13 N_16 RN GND GND mn15  l=0.13u w=0.28u m=1
M14 GND N_24 Q GND mn15  l=0.13u w=0.46u m=1
M15 GND N_24 Q GND mn15  l=0.13u w=0.46u m=1
M16 N_7 SN GND GND mn15  l=0.13u w=0.31u m=1
M17 GND SN N_7 GND mn15  l=0.13u w=0.31u m=1
M18 GND SN N_7 GND mn15  l=0.13u w=0.31u m=1
M19 N_12 N_16 N_7 GND mn15  l=0.13u w=0.37u m=1
M20 GND N_12 QN GND mn15  l=0.13u w=0.46u m=1
M21 GND N_12 QN GND mn15  l=0.13u w=0.46u m=1
M22 GND N_12 N_24 GND mn15  l=0.13u w=0.36u m=1
M23 VDD N_12 QN VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_12 QN VDD mp15  l=0.13u w=0.69u m=1
M25 N_24 N_12 VDD VDD mp15  l=0.13u w=0.54u m=1
M26 VDD RN N_16 VDD mp15  l=0.13u w=0.42u m=1
M27 Q N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_24 Q VDD mp15  l=0.13u w=0.69u m=1
M29 N_5 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M30 N_43 D VDD VDD mp15  l=0.13u w=0.63u m=1
M31 N_44 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_43 N_2 N_6 VDD mp15  l=0.13u w=0.63u m=1
M33 N_2 N_5 VDD VDD mp15  l=0.13u w=0.42u m=1
M34 N_44 N_5 N_6 VDD mp15  l=0.13u w=0.17u m=1
M35 N_36 N_24 N_45 VDD mp15  l=0.13u w=0.17u m=1
M36 N_12 SN VDD VDD mp15  l=0.13u w=0.58u m=1
M37 N_36 N_16 VDD VDD mp15  l=0.13u w=0.41u m=1
M38 N_36 N_16 VDD VDD mp15  l=0.13u w=0.41u m=1
M39 VDD N_16 N_36 VDD mp15  l=0.13u w=0.41u m=1
M40 N_9 N_6 N_36 VDD mp15  l=0.13u w=0.315u m=1
M41 N_9 N_6 N_36 VDD mp15  l=0.13u w=0.315u m=1
M42 N_9 N_6 N_36 VDD mp15  l=0.13u w=0.315u m=1
M43 N_9 N_6 N_36 VDD mp15  l=0.13u w=0.315u m=1
M44 N_45 N_2 N_12 VDD mp15  l=0.13u w=0.17u m=1
M45 N_12 N_5 N_9 VDD mp15  l=0.13u w=0.55u m=1
.ends dfbrb2
* SPICE INPUT		Tue Jul 31 19:14:36 2018	dfbrbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrbm
.subckt dfbrbm GND Q QN VDD RN D SN CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.2u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_21 D GND GND mn15  l=0.13u w=0.28u m=1
M4 N_22 N_2 N_7 GND mn15  l=0.13u w=0.17u m=1
M5 N_22 N_16 GND GND mn15  l=0.13u w=0.17u m=1
M6 N_21 N_4 N_7 GND mn15  l=0.13u w=0.28u m=1
M7 Q N_13 GND GND mn15  l=0.13u w=0.36u m=1
M8 N_10 RN GND GND mn15  l=0.13u w=0.17u m=1
M9 QN N_17 GND GND mn15  l=0.13u w=0.36u m=1
M10 N_13 N_17 GND GND mn15  l=0.13u w=0.22u m=1
M11 N_16 N_7 N_14 GND mn15  l=0.13u w=0.28u m=1
M12 N_17 N_2 N_16 GND mn15  l=0.13u w=0.28u m=1
M13 N_17 N_4 N_23 GND mn15  l=0.13u w=0.17u m=1
M14 N_23 N_13 N_14 GND mn15  l=0.13u w=0.17u m=1
M15 N_17 N_10 N_14 GND mn15  l=0.13u w=0.22u m=1
M16 N_14 SN GND GND mn15  l=0.13u w=0.46u m=1
M17 N_4 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M18 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M19 N_90 D VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_90 N_2 N_7 VDD mp15  l=0.13u w=0.42u m=1
M21 N_89 N_16 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_7 N_4 N_89 VDD mp15  l=0.13u w=0.17u m=1
M23 Q N_13 VDD VDD mp15  l=0.13u w=0.55u m=1
M24 N_10 RN VDD VDD mp15  l=0.13u w=0.24u m=1
M25 N_28 N_13 N_30 VDD mp15  l=0.13u w=0.17u m=1
M26 N_28 N_10 VDD VDD mp15  l=0.13u w=0.61u m=1
M27 N_17 SN VDD VDD mp15  l=0.13u w=0.31u m=1
M28 N_16 N_7 N_28 VDD mp15  l=0.13u w=0.54u m=1
M29 N_17 N_2 N_30 VDD mp15  l=0.13u w=0.17u m=1
M30 N_17 N_4 N_16 VDD mp15  l=0.13u w=0.44u m=1
M31 QN N_17 VDD VDD mp15  l=0.13u w=0.55u m=1
M32 N_13 N_17 VDD VDD mp15  l=0.13u w=0.31u m=1
.ends dfbrbm
* SPICE INPUT		Tue Jul 31 19:14:48 2018	dfbrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq0
.subckt dfbrq0 GND Q VDD RN SN D CK
M1 N_5 N_11 N_4 GND mn15  l=0.13u w=0.2u m=1
M2 N_5 SN GND GND mn15  l=0.13u w=0.37u m=1
M3 GND N_4 N_2 GND mn15  l=0.13u w=0.18u m=1
M4 N_8 CK GND GND mn15  l=0.13u w=0.18u m=1
M5 GND N_8 N_6 GND mn15  l=0.13u w=0.17u m=1
M6 Q N_2 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_11 RN GND GND mn15  l=0.13u w=0.18u m=1
M8 N_19 D GND GND mn15  l=0.13u w=0.26u m=1
M9 N_20 N_6 N_14 GND mn15  l=0.13u w=0.17u m=1
M10 N_20 N_16 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_14 N_8 N_19 GND mn15  l=0.13u w=0.26u m=1
M12 N_5 N_14 N_16 GND mn15  l=0.13u w=0.28u m=1
M13 N_4 N_6 N_16 GND mn15  l=0.13u w=0.28u m=1
M14 N_4 N_8 N_21 GND mn15  l=0.13u w=0.17u m=1
M15 N_21 N_2 N_5 GND mn15  l=0.13u w=0.17u m=1
M16 N_2 N_4 VDD VDD mp15  l=0.13u w=0.26u m=1
M17 Q N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_11 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M19 N_8 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M20 N_6 N_8 VDD VDD mp15  l=0.13u w=0.42u m=1
M21 N_28 N_2 N_29 VDD mp15  l=0.13u w=0.17u m=1
M22 N_28 N_11 VDD VDD mp15  l=0.13u w=0.585u m=1
M23 N_4 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M24 N_84 D VDD VDD mp15  l=0.13u w=0.37u m=1
M25 N_84 N_6 N_14 VDD mp15  l=0.13u w=0.37u m=1
M26 N_83 N_16 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_14 N_8 N_83 VDD mp15  l=0.13u w=0.17u m=1
M28 N_28 N_14 N_16 VDD mp15  l=0.13u w=0.45u m=1
M29 N_4 N_6 N_29 VDD mp15  l=0.13u w=0.17u m=1
M30 N_4 N_8 N_16 VDD mp15  l=0.13u w=0.46u m=1
.ends dfbrq0
* SPICE INPUT		Tue Jul 31 19:15:00 2018	dfbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq1
.subckt dfbrq1 GND Q VDD CK D SN RN
M1 N_19 N_16 GND GND mn15  l=0.13u w=0.17u m=1
M2 N_20 D GND GND mn15  l=0.13u w=0.28u m=1
M3 N_4 N_9 N_19 GND mn15  l=0.13u w=0.17u m=1
M4 N_20 N_11 N_4 GND mn15  l=0.13u w=0.28u m=1
M5 N_8 SN GND GND mn15  l=0.13u w=0.46u m=1
M6 N_8 N_14 N_7 GND mn15  l=0.13u w=0.28u m=1
M7 N_6 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_11 CK GND GND mn15  l=0.13u w=0.2u m=1
M9 GND N_11 N_9 GND mn15  l=0.13u w=0.17u m=1
M10 N_14 RN GND GND mn15  l=0.13u w=0.18u m=1
M11 Q N_6 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_7 N_11 N_21 GND mn15  l=0.13u w=0.17u m=1
M13 N_21 N_6 N_8 GND mn15  l=0.13u w=0.17u m=1
M14 N_7 N_9 N_16 GND mn15  l=0.13u w=0.41u m=1
M15 N_8 N_4 N_16 GND mn15  l=0.13u w=0.4u m=1
M16 N_30 N_14 VDD VDD mp15  l=0.13u w=0.35u m=1
M17 VDD N_14 N_30 VDD mp15  l=0.13u w=0.35u m=1
M18 N_35 N_16 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 N_36 D VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_4 N_11 N_35 VDD mp15  l=0.13u w=0.17u m=1
M21 N_36 N_9 N_4 VDD mp15  l=0.13u w=0.42u m=1
M22 N_11 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M23 N_9 N_11 VDD VDD mp15  l=0.13u w=0.44u m=1
M24 N_14 RN VDD VDD mp15  l=0.13u w=0.28u m=1
M25 Q N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_37 N_6 N_30 VDD mp15  l=0.13u w=0.17u m=1
M27 N_37 N_9 N_7 VDD mp15  l=0.13u w=0.17u m=1
M28 N_7 N_11 N_16 VDD mp15  l=0.13u w=0.57u m=1
M29 N_16 N_4 N_30 VDD mp15  l=0.13u w=0.39u m=1
M30 N_16 N_4 N_30 VDD mp15  l=0.13u w=0.28u m=1
M31 N_7 SN VDD VDD mp15  l=0.13u w=0.37u m=1
M32 N_6 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends dfbrq1
* SPICE INPUT		Tue Jul 31 19:15:12 2018	dfbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfbrq2
.subckt dfbrq2 GND Q VDD RN D CK SN
M1 GND CK N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_23 D GND GND mn15  l=0.13u w=0.43u m=1
M3 N_24 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M4 N_24 N_2 N_6 GND mn15  l=0.13u w=0.17u m=1
M5 N_23 N_4 N_6 GND mn15  l=0.13u w=0.43u m=1
M6 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M7 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M8 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND RN N_9 GND mn15  l=0.13u w=0.28u m=1
M10 N_8 N_17 GND GND mn15  l=0.13u w=0.37u m=1
M11 N_13 N_6 N_12 GND mn15  l=0.13u w=0.18u m=1
M12 N_12 N_6 N_13 GND mn15  l=0.13u w=0.26u m=1
M13 N_12 N_6 N_13 GND mn15  l=0.13u w=0.17u m=1
M14 N_17 N_2 N_13 GND mn15  l=0.13u w=0.42u m=1
M15 N_17 N_4 N_25 GND mn15  l=0.13u w=0.17u m=1
M16 N_25 N_8 N_12 GND mn15  l=0.13u w=0.17u m=1
M17 N_17 N_9 N_12 GND mn15  l=0.13u w=0.36u m=1
M18 N_12 SN GND GND mn15  l=0.13u w=0.305u m=1
M19 GND SN N_12 GND mn15  l=0.13u w=0.305u m=1
M20 GND SN N_12 GND mn15  l=0.13u w=0.3u m=1
M21 N_4 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_40 D VDD VDD mp15  l=0.13u w=0.63u m=1
M23 N_41 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 N_40 N_2 N_6 VDD mp15  l=0.13u w=0.63u m=1
M25 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M26 N_41 N_4 N_6 VDD mp15  l=0.13u w=0.17u m=1
M27 N_13 N_6 N_35 VDD mp15  l=0.13u w=0.31u m=1
M28 N_13 N_6 N_35 VDD mp15  l=0.13u w=0.31u m=1
M29 N_13 N_6 N_35 VDD mp15  l=0.13u w=0.31u m=1
M30 N_13 N_6 N_35 VDD mp15  l=0.13u w=0.31u m=1
M31 N_17 N_4 N_13 VDD mp15  l=0.13u w=0.55u m=1
M32 N_42 N_2 N_17 VDD mp15  l=0.13u w=0.17u m=1
M33 N_42 N_8 N_35 VDD mp15  l=0.13u w=0.17u m=1
M34 N_35 N_9 VDD VDD mp15  l=0.13u w=0.42u m=1
M35 N_35 N_9 VDD VDD mp15  l=0.13u w=0.42u m=1
M36 VDD N_9 N_35 VDD mp15  l=0.13u w=0.41u m=1
M37 N_17 SN VDD VDD mp15  l=0.13u w=0.56u m=1
M38 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M40 VDD RN N_9 VDD mp15  l=0.13u w=0.42u m=1
M41 N_8 N_17 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends dfbrq2
* SPICE INPUT		Tue Jul 31 19:15:24 2018	dfcfb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb0
.subckt dfcfb0 VDD Q QN GND RN D CKN
M1 GND CKN N_4 GND mn15  l=0.13u w=0.2u m=1
M2 N_29 D GND GND mn15  l=0.13u w=0.26u m=1
M3 N_29 N_2 N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_30 N_8 GND GND mn15  l=0.13u w=0.17u m=1
M5 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M6 N_30 N_4 N_5 GND mn15  l=0.13u w=0.17u m=1
M7 N_8 N_5 GND GND mn15  l=0.13u w=0.24u m=1
M8 GND N_15 N_9 GND mn15  l=0.13u w=0.18u m=1
M9 N_9 N_4 N_8 GND mn15  l=0.13u w=0.23u m=1
M10 N_31 N_2 N_9 GND mn15  l=0.13u w=0.17u m=1
M11 GND N_18 N_31 GND mn15  l=0.13u w=0.17u m=1
M12 QN N_9 GND GND mn15  l=0.13u w=0.26u m=1
M13 N_18 N_9 GND GND mn15  l=0.13u w=0.18u m=1
M14 N_15 RN GND GND mn15  l=0.13u w=0.17u m=1
M15 Q N_18 GND GND mn15  l=0.13u w=0.26u m=1
M16 N_4 CKN VDD VDD mp15  l=0.13u w=0.51u m=1
M17 N_19 D VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_20 N_2 N_5 VDD mp15  l=0.13u w=0.17u m=1
M19 N_20 N_8 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 VDD N_4 N_2 VDD mp15  l=0.13u w=0.42u m=1
M21 N_19 N_4 N_5 VDD mp15  l=0.13u w=0.4u m=1
M22 N_9 N_2 N_8 VDD mp15  l=0.13u w=0.44u m=1
M23 N_8 N_5 N_7 VDD mp15  l=0.13u w=0.45u m=1
M24 N_21 N_4 N_9 VDD mp15  l=0.13u w=0.17u m=1
M25 N_7 N_15 VDD VDD mp15  l=0.13u w=0.59u m=1
M26 N_21 N_18 N_7 VDD mp15  l=0.13u w=0.17u m=1
M27 N_15 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M28 VDD N_18 Q VDD mp15  l=0.13u w=0.4u m=1
M29 QN N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M30 N_18 N_9 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends dfcfb0
* SPICE INPUT		Tue Jul 31 19:15:39 2018	dfcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb1
.subckt dfcfb1 GND QN Q VDD CKN D RN
M1 GND CKN N_4 GND mn15  l=0.13u w=0.2u m=1
M2 N_19 D GND GND mn15  l=0.13u w=0.28u m=1
M3 N_19 N_2 N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_20 N_11 GND GND mn15  l=0.13u w=0.17u m=1
M5 GND N_4 N_2 GND mn15  l=0.13u w=0.2u m=1
M6 N_20 N_4 N_6 GND mn15  l=0.13u w=0.17u m=1
M7 QN N_10 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_9 N_10 GND GND mn15  l=0.13u w=0.27u m=1
M9 N_21 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M10 N_11 N_6 GND GND mn15  l=0.13u w=0.21u m=1
M11 GND N_6 N_11 GND mn15  l=0.13u w=0.2u m=1
M12 GND N_18 N_10 GND mn15  l=0.13u w=0.27u m=1
M13 N_11 N_4 N_10 GND mn15  l=0.13u w=0.37u m=1
M14 N_21 N_2 N_10 GND mn15  l=0.13u w=0.17u m=1
M15 Q N_9 GND GND mn15  l=0.13u w=0.43u m=1
M16 N_18 RN GND GND mn15  l=0.13u w=0.18u m=1
M17 QN N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_9 N_10 VDD VDD mp15  l=0.13u w=0.39u m=1
M19 N_83 N_9 N_29 VDD mp15  l=0.13u w=0.17u m=1
M20 N_83 N_4 N_10 VDD mp15  l=0.13u w=0.17u m=1
M21 N_29 N_18 VDD VDD mp15  l=0.13u w=0.665u m=1
M22 N_11 N_2 N_10 VDD mp15  l=0.13u w=0.285u m=1
M23 N_10 N_2 N_11 VDD mp15  l=0.13u w=0.285u m=1
M24 N_11 N_6 N_29 VDD mp15  l=0.13u w=0.58u m=1
M25 N_4 CKN VDD VDD mp15  l=0.13u w=0.51u m=1
M26 N_84 D VDD VDD mp15  l=0.13u w=0.42u m=1
M27 N_85 N_2 N_6 VDD mp15  l=0.13u w=0.17u m=1
M28 N_85 N_11 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 VDD N_4 N_2 VDD mp15  l=0.13u w=0.51u m=1
M30 N_84 N_4 N_6 VDD mp15  l=0.13u w=0.42u m=1
M31 Q N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 N_18 RN VDD VDD mp15  l=0.13u w=0.28u m=1
.ends dfcfb1
* SPICE INPUT		Tue Jul 31 19:15:53 2018	dfcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcfb2
.subckt dfcfb2 GND Q QN VDD RN D CKN
M1 GND CKN N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_23 D GND GND mn15  l=0.13u w=0.41u m=1
M3 N_23 N_2 N_6 GND mn15  l=0.13u w=0.41u m=1
M4 N_24 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M5 GND N_4 N_2 GND mn15  l=0.13u w=0.22u m=1
M6 N_24 N_4 N_6 GND mn15  l=0.13u w=0.17u m=1
M7 GND N_6 N_7 GND mn15  l=0.13u w=0.23u m=1
M8 GND N_6 N_7 GND mn15  l=0.13u w=0.23u m=1
M9 N_8 N_4 N_7 GND mn15  l=0.13u w=0.46u m=1
M10 N_8 N_17 GND GND mn15  l=0.13u w=0.18u m=1
M11 GND N_17 N_8 GND mn15  l=0.13u w=0.18u m=1
M12 N_25 N_2 N_8 GND mn15  l=0.13u w=0.17u m=1
M13 GND N_21 N_25 GND mn15  l=0.13u w=0.17u m=1
M14 GND RN N_17 GND mn15  l=0.13u w=0.28u m=1
M15 GND N_21 Q GND mn15  l=0.13u w=0.46u m=1
M16 GND N_21 Q GND mn15  l=0.13u w=0.43u m=1
M17 GND N_8 QN GND mn15  l=0.13u w=0.46u m=1
M18 GND N_8 QN GND mn15  l=0.13u w=0.46u m=1
M19 GND N_8 N_21 GND mn15  l=0.13u w=0.37u m=1
M20 N_4 CKN VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_101 D VDD VDD mp15  l=0.13u w=0.62u m=1
M22 N_101 N_4 N_6 VDD mp15  l=0.13u w=0.62u m=1
M23 N_102 N_2 N_6 VDD mp15  l=0.13u w=0.17u m=1
M24 N_102 N_7 VDD VDD mp15  l=0.13u w=0.17u m=1
M25 N_2 N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
M26 N_7 N_2 N_8 VDD mp15  l=0.13u w=0.35u m=1
M27 N_7 N_2 N_8 VDD mp15  l=0.13u w=0.35u m=1
M28 N_7 N_6 N_31 VDD mp15  l=0.13u w=0.46u m=1
M29 N_31 N_6 N_7 VDD mp15  l=0.13u w=0.44u m=1
M30 N_31 N_6 N_7 VDD mp15  l=0.13u w=0.44u m=1
M31 N_103 N_4 N_8 VDD mp15  l=0.13u w=0.17u m=1
M32 VDD N_17 N_31 VDD mp15  l=0.13u w=0.67u m=1
M33 N_31 N_17 VDD VDD mp15  l=0.13u w=0.67u m=1
M34 N_31 N_21 N_103 VDD mp15  l=0.13u w=0.17u m=1
M35 N_17 RN VDD VDD mp15  l=0.13u w=0.42u m=1
M36 Q N_21 VDD VDD mp15  l=0.13u w=0.69u m=1
M37 VDD N_21 Q VDD mp15  l=0.13u w=0.69u m=1
M38 VDD N_8 QN VDD mp15  l=0.13u w=0.69u m=1
M39 VDD N_8 QN VDD mp15  l=0.13u w=0.69u m=1
M40 VDD N_8 N_21 VDD mp15  l=0.13u w=0.55u m=1
.ends dfcfb2
* SPICE INPUT		Tue Jul 31 19:16:05 2018	dfcrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb0
.subckt dfcrb0 VDD Q QN GND RN D CK
M1 GND CK N_5 GND mn15  l=0.13u w=0.18u m=1
M2 N_77 D GND GND mn15  l=0.13u w=0.26u m=1
M3 N_77 N_5 N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_78 N_8 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_78 N_2 N_6 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_5 N_2 GND mn15  l=0.13u w=0.17u m=1
M7 N_8 N_6 GND GND mn15  l=0.13u w=0.24u m=1
M8 N_10 N_2 N_8 GND mn15  l=0.13u w=0.23u m=1
M9 N_79 N_5 N_10 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_16 N_10 GND mn15  l=0.13u w=0.18u m=1
M11 N_79 N_19 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_16 RN GND GND mn15  l=0.13u w=0.17u m=1
M13 Q N_19 GND GND mn15  l=0.13u w=0.26u m=1
M14 QN N_10 GND GND mn15  l=0.13u w=0.26u m=1
M15 N_19 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M16 N_5 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M17 N_20 D VDD VDD mp15  l=0.13u w=0.37u m=1
M18 N_21 N_8 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 N_20 N_2 N_6 VDD mp15  l=0.13u w=0.37u m=1
M20 VDD N_5 N_2 VDD mp15  l=0.13u w=0.42u m=1
M21 N_21 N_5 N_6 VDD mp15  l=0.13u w=0.17u m=1
M22 N_8 N_6 N_7 VDD mp15  l=0.13u w=0.2u m=1
M23 N_7 N_6 N_8 VDD mp15  l=0.13u w=0.2u m=1
M24 N_10 N_2 N_22 VDD mp15  l=0.13u w=0.17u m=1
M25 N_22 N_19 N_7 VDD mp15  l=0.13u w=0.17u m=1
M26 N_8 N_5 N_10 VDD mp15  l=0.13u w=0.44u m=1
M27 N_7 N_16 VDD VDD mp15  l=0.13u w=0.59u m=1
M28 N_16 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M29 Q N_19 VDD VDD mp15  l=0.13u w=0.4u m=1
M30 QN N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M31 N_19 N_10 VDD VDD mp15  l=0.13u w=0.28u m=1
.ends dfcrb0
* SPICE INPUT		Tue Jul 31 19:16:20 2018	dfcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb1
.subckt dfcrb1 GND QN Q VDD RN D CK
M1 QN N_11 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 N_11 GND GND mn15  l=0.13u w=0.28u m=1
M3 GND CK N_7 GND mn15  l=0.13u w=0.2u m=1
M4 N_19 D GND GND mn15  l=0.13u w=0.28u m=1
M5 N_19 N_7 N_9 GND mn15  l=0.13u w=0.28u m=1
M6 N_20 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M7 N_20 N_5 N_9 GND mn15  l=0.13u w=0.17u m=1
M8 GND N_7 N_5 GND mn15  l=0.13u w=0.17u m=1
M9 GND N_9 N_12 GND mn15  l=0.13u w=0.19u m=1
M10 N_12 N_9 GND GND mn15  l=0.13u w=0.18u m=1
M11 N_11 N_5 N_12 GND mn15  l=0.13u w=0.37u m=1
M12 N_21 N_7 N_11 GND mn15  l=0.13u w=0.17u m=1
M13 N_11 N_18 GND GND mn15  l=0.13u w=0.28u m=1
M14 N_21 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M15 N_18 RN GND GND mn15  l=0.13u w=0.2u m=1
M16 Q N_4 GND GND mn15  l=0.13u w=0.44u m=1
M17 QN N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_4 N_11 VDD VDD mp15  l=0.13u w=0.41u m=1
M19 N_7 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M20 N_82 D VDD VDD mp15  l=0.13u w=0.42u m=1
M21 N_83 N_12 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_82 N_5 N_9 VDD mp15  l=0.13u w=0.42u m=1
M23 VDD N_7 N_5 VDD mp15  l=0.13u w=0.42u m=1
M24 N_83 N_7 N_9 VDD mp15  l=0.13u w=0.17u m=1
M25 N_12 N_9 N_27 VDD mp15  l=0.13u w=0.35u m=1
M26 N_27 N_9 N_12 VDD mp15  l=0.13u w=0.35u m=1
M27 N_11 N_5 N_84 VDD mp15  l=0.13u w=0.17u m=1
M28 N_84 N_4 N_27 VDD mp15  l=0.13u w=0.17u m=1
M29 N_11 N_7 N_12 VDD mp15  l=0.13u w=0.52u m=1
M30 N_27 N_18 VDD VDD mp15  l=0.13u w=0.35u m=1
M31 VDD N_18 N_27 VDD mp15  l=0.13u w=0.35u m=1
M32 N_18 RN VDD VDD mp15  l=0.13u w=0.29u m=1
M33 Q N_4 VDD VDD mp15  l=0.13u w=0.68u m=1
.ends dfcrb1
* SPICE INPUT		Tue Jul 31 19:16:32 2018	dfcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrb2
.subckt dfcrb2 GND QN Q VDD RN D CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.22u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.19u m=1
M3 GND D N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_19 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M5 N_20 N_2 N_8 GND mn15  l=0.13u w=0.17u m=1
M6 N_20 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M7 N_11 N_2 N_10 GND mn15  l=0.13u w=0.38u m=1
M8 N_10 N_8 N_21 GND mn15  l=0.13u w=0.45u m=1
M9 N_19 N_4 N_8 GND mn15  l=0.13u w=0.28u m=1
M10 N_22 N_4 N_11 GND mn15  l=0.13u w=0.17u m=1
M11 N_23 N_17 N_22 GND mn15  l=0.13u w=0.17u m=1
M12 N_21 RN GND GND mn15  l=0.13u w=0.45u m=1
M13 N_23 RN GND GND mn15  l=0.13u w=0.17u m=1
M14 GND N_17 QN GND mn15  l=0.13u w=0.46u m=1
M15 GND N_17 QN GND mn15  l=0.13u w=0.46u m=1
M16 GND N_11 Q GND mn15  l=0.13u w=0.46u m=1
M17 GND N_11 Q GND mn15  l=0.13u w=0.46u m=1
M18 GND N_11 N_17 GND mn15  l=0.13u w=0.37u m=1
M19 N_4 CK VDD VDD mp15  l=0.13u w=0.55u m=1
M20 N_2 N_4 VDD VDD mp15  l=0.13u w=0.49u m=1
M21 N_6 D VDD VDD mp15  l=0.13u w=0.42u m=1
M22 N_37 N_6 VDD VDD mp15  l=0.13u w=0.41u m=1
M23 N_37 N_2 N_8 VDD mp15  l=0.13u w=0.41u m=1
M24 N_38 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M25 N_10 N_8 VDD VDD mp15  l=0.13u w=0.21u m=1
M26 VDD N_8 N_10 VDD mp15  l=0.13u w=0.16u m=1
M27 N_10 N_8 VDD VDD mp15  l=0.13u w=0.16u m=1
M28 N_11 N_4 N_10 VDD mp15  l=0.13u w=0.59u m=1
M29 N_38 N_4 N_8 VDD mp15  l=0.13u w=0.17u m=1
M30 N_39 N_2 N_11 VDD mp15  l=0.13u w=0.28u m=1
M31 N_39 N_17 VDD VDD mp15  l=0.13u w=0.28u m=1
M32 N_11 RN VDD VDD mp15  l=0.13u w=0.56u m=1
M33 N_10 RN VDD VDD mp15  l=0.13u w=0.37u m=1
M34 VDD RN N_10 VDD mp15  l=0.13u w=0.16u m=1
M35 QN N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 VDD N_17 QN VDD mp15  l=0.13u w=0.69u m=1
M37 VDD N_11 Q VDD mp15  l=0.13u w=0.69u m=1
M38 VDD N_11 Q VDD mp15  l=0.13u w=0.69u m=1
M39 N_17 N_11 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends dfcrb2
* SPICE INPUT		Tue Jul 31 19:16:45 2018	dfcrbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrbm
.subckt dfcrbm GND Q QN VDD RN D CK
M1 GND CK N_4 GND mn15  l=0.13u w=0.19u m=1
M2 N_19 D GND GND mn15  l=0.13u w=0.28u m=1
M3 N_19 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_20 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_20 N_2 N_6 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M7 GND N_6 N_9 GND mn15  l=0.13u w=0.14u m=1
M8 N_9 N_6 GND GND mn15  l=0.13u w=0.14u m=1
M9 N_7 N_2 N_9 GND mn15  l=0.13u w=0.28u m=1
M10 N_21 N_4 N_7 GND mn15  l=0.13u w=0.17u m=1
M11 GND N_15 N_7 GND mn15  l=0.13u w=0.22u m=1
M12 N_21 N_18 GND GND mn15  l=0.13u w=0.17u m=1
M13 N_15 RN GND GND mn15  l=0.13u w=0.17u m=1
M14 Q N_18 GND GND mn15  l=0.13u w=0.36u m=1
M15 QN N_7 GND GND mn15  l=0.13u w=0.36u m=1
M16 N_18 N_7 GND GND mn15  l=0.13u w=0.22u m=1
M17 N_4 CK VDD VDD mp15  l=0.13u w=0.49u m=1
M18 N_82 D VDD VDD mp15  l=0.13u w=0.42u m=1
M19 N_83 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 N_82 N_2 N_6 VDD mp15  l=0.13u w=0.42u m=1
M21 VDD N_4 N_2 VDD mp15  l=0.13u w=0.42u m=1
M22 N_83 N_4 N_6 VDD mp15  l=0.13u w=0.17u m=1
M23 N_9 N_6 N_28 VDD mp15  l=0.13u w=0.28u m=1
M24 N_28 N_6 N_9 VDD mp15  l=0.13u w=0.28u m=1
M25 N_7 N_2 N_84 VDD mp15  l=0.13u w=0.17u m=1
M26 N_84 N_18 N_28 VDD mp15  l=0.13u w=0.17u m=1
M27 N_9 N_4 N_7 VDD mp15  l=0.13u w=0.46u m=1
M28 N_28 N_15 VDD VDD mp15  l=0.13u w=0.325u m=1
M29 VDD N_15 N_28 VDD mp15  l=0.13u w=0.325u m=1
M30 N_15 RN VDD VDD mp15  l=0.13u w=0.24u m=1
M31 Q N_18 VDD VDD mp15  l=0.13u w=0.55u m=1
M32 QN N_7 VDD VDD mp15  l=0.13u w=0.55u m=1
M33 N_18 N_7 VDD VDD mp15  l=0.13u w=0.31u m=1
.ends dfcrbm
* SPICE INPUT		Tue Jul 31 19:16:56 2018	dfcrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq0
.subckt dfcrq0 GND Q D VDD RN CK
M1 Q N_13 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M3 GND N_7 N_5 GND mn15  l=0.13u w=0.17u m=1
M4 N_7 CK GND GND mn15  l=0.13u w=0.17u m=1
M5 N_11 N_7 N_16 GND mn15  l=0.13u w=0.17u m=1
M6 N_19 N_7 N_13 GND mn15  l=0.13u w=0.17u m=1
M7 N_17 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_14 N_11 N_18 GND mn15  l=0.13u w=0.28u m=1
M9 GND D N_9 GND mn15  l=0.13u w=0.175u m=1
M10 N_16 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_17 N_5 N_11 GND mn15  l=0.13u w=0.17u m=1
M12 N_18 RN GND GND mn15  l=0.13u w=0.28u m=1
M13 N_15 RN GND GND mn15  l=0.13u w=0.17u m=1
M14 N_19 N_4 N_15 GND mn15  l=0.13u w=0.17u m=1
M15 N_14 N_5 N_13 GND mn15  l=0.13u w=0.28u m=1
M16 N_5 N_7 VDD VDD mp15  l=0.13u w=0.28u m=1
M17 N_7 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M18 N_33 N_7 N_11 VDD mp15  l=0.13u w=0.17u m=1
M19 N_33 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 N_14 N_11 VDD VDD mp15  l=0.13u w=0.31u m=1
M21 VDD D N_9 VDD mp15  l=0.13u w=0.26u m=1
M22 N_32 N_9 VDD VDD mp15  l=0.13u w=0.28u m=1
M23 VDD RN N_14 VDD mp15  l=0.13u w=0.31u m=1
M24 N_11 N_5 N_32 VDD mp15  l=0.13u w=0.28u m=1
M25 Q N_13 VDD VDD mp15  l=0.13u w=0.4u m=1
M26 N_4 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_13 N_7 N_14 VDD mp15  l=0.13u w=0.28u m=1
M28 N_34 N_5 N_13 VDD mp15  l=0.13u w=0.28u m=1
M29 N_13 RN VDD VDD mp15  l=0.13u w=0.28u m=1
M30 N_34 N_4 VDD VDD mp15  l=0.13u w=0.28u m=1
.ends dfcrq0
* SPICE INPUT		Tue Jul 31 19:17:08 2018	dfcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq1
.subckt dfcrq1 GND Q VDD RN D CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.2u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.2u m=1
M3 GND D N_6 GND mn15  l=0.13u w=0.175u m=1
M4 N_16 N_6 GND GND mn15  l=0.13u w=0.3u m=1
M5 N_17 N_2 N_8 GND mn15  l=0.13u w=0.17u m=1
M6 N_10 N_8 N_18 GND mn15  l=0.13u w=0.36u m=1
M7 N_11 N_2 N_10 GND mn15  l=0.13u w=0.31u m=1
M8 N_16 N_4 N_8 GND mn15  l=0.13u w=0.3u m=1
M9 N_19 N_4 N_11 GND mn15  l=0.13u w=0.17u m=1
M10 N_18 RN GND GND mn15  l=0.13u w=0.36u m=1
M11 N_15 RN GND GND mn15  l=0.13u w=0.17u m=1
M12 N_19 N_14 N_15 GND mn15  l=0.13u w=0.17u m=1
M13 N_17 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M14 Q N_11 GND GND mn15  l=0.13u w=0.46u m=1
M15 N_14 N_11 GND GND mn15  l=0.13u w=0.28u m=1
M16 N_4 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M17 N_2 N_4 VDD VDD mp15  l=0.13u w=0.51u m=1
M18 Q N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_14 N_11 VDD VDD mp15  l=0.13u w=0.28u m=1
M20 VDD D N_6 VDD mp15  l=0.13u w=0.28u m=1
M21 N_32 N_6 VDD VDD mp15  l=0.13u w=0.42u m=1
M22 N_8 N_2 N_32 VDD mp15  l=0.13u w=0.42u m=1
M23 N_10 N_8 VDD VDD mp15  l=0.13u w=0.18u m=1
M24 VDD N_8 N_10 VDD mp15  l=0.13u w=0.17u m=1
M25 N_11 N_4 N_10 VDD mp15  l=0.13u w=0.5u m=1
M26 N_33 N_4 N_8 VDD mp15  l=0.13u w=0.17u m=1
M27 N_34 N_2 N_11 VDD mp15  l=0.13u w=0.28u m=1
M28 N_11 RN VDD VDD mp15  l=0.13u w=0.34u m=1
M29 N_10 RN VDD VDD mp15  l=0.13u w=0.35u m=1
M30 N_34 N_14 VDD VDD mp15  l=0.13u w=0.28u m=1
M31 N_33 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
.ends dfcrq1
* SPICE INPUT		Tue Jul 31 19:17:22 2018	dfcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq2
.subckt dfcrq2 GND Q VDD RN D CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.27u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.22u m=1
M3 GND D N_6 GND mn15  l=0.13u w=0.23u m=1
M4 N_17 N_6 GND GND mn15  l=0.13u w=0.35u m=1
M5 N_18 N_2 N_8 GND mn15  l=0.13u w=0.17u m=1
M6 N_18 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M7 N_11 N_2 N_10 GND mn15  l=0.13u w=0.36u m=1
M8 N_10 N_8 N_19 GND mn15  l=0.13u w=0.44u m=1
M9 N_8 N_4 N_17 GND mn15  l=0.13u w=0.35u m=1
M10 N_21 N_4 N_11 GND mn15  l=0.13u w=0.17u m=1
M11 N_21 N_14 N_20 GND mn15  l=0.13u w=0.17u m=1
M12 N_19 RN GND GND mn15  l=0.13u w=0.44u m=1
M13 N_20 RN GND GND mn15  l=0.13u w=0.17u m=1
M14 Q N_11 GND GND mn15  l=0.13u w=0.305u m=1
M15 Q N_11 GND GND mn15  l=0.13u w=0.305u m=1
M16 Q N_11 GND GND mn15  l=0.13u w=0.3u m=1
M17 GND N_11 N_14 GND mn15  l=0.13u w=0.28u m=1
M18 N_4 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M19 N_2 N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
M20 N_6 D VDD VDD mp15  l=0.13u w=0.35u m=1
M21 N_34 N_6 VDD VDD mp15  l=0.13u w=0.52u m=1
M22 N_8 N_2 N_34 VDD mp15  l=0.13u w=0.52u m=1
M23 N_35 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 N_10 N_8 VDD VDD mp15  l=0.13u w=0.2u m=1
M25 VDD N_8 N_10 VDD mp15  l=0.13u w=0.17u m=1
M26 N_10 N_8 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_11 N_4 N_10 VDD mp15  l=0.13u w=0.53u m=1
M28 N_35 N_4 N_8 VDD mp15  l=0.13u w=0.17u m=1
M29 VDD N_11 Q VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_11 Q VDD mp15  l=0.13u w=0.69u m=1
M31 N_14 N_11 VDD VDD mp15  l=0.13u w=0.28u m=1
M32 N_36 N_2 N_11 VDD mp15  l=0.13u w=0.28u m=1
M33 VDD N_14 N_36 VDD mp15  l=0.13u w=0.28u m=1
M34 VDD RN N_10 VDD mp15  l=0.13u w=0.27u m=1
M35 N_10 RN VDD VDD mp15  l=0.13u w=0.27u m=1
M36 VDD RN N_11 VDD mp15  l=0.13u w=0.19u m=1
M37 N_11 RN VDD VDD mp15  l=0.13u w=0.28u m=1
.ends dfcrq2
* SPICE INPUT		Tue Jul 31 19:17:37 2018	dfcrq3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrq3
.subckt dfcrq3 VDD Q GND RN D CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.28u m=1
M2 GND N_4 N_3 GND mn15  l=0.13u w=0.22u m=1
M3 GND D N_8 GND mn15  l=0.13u w=0.28u m=1
M4 N_34 N_8 GND GND mn15  l=0.13u w=0.36u m=1
M5 N_9 N_3 N_33 GND mn15  l=0.13u w=0.17u m=1
M6 N_33 N_6 GND GND mn15  l=0.13u w=0.17u m=1
M7 N_9 N_4 N_34 GND mn15  l=0.13u w=0.36u m=1
M8 N_28 N_9 N_6 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 N_4 N_30 GND mn15  l=0.13u w=0.17u m=1
M10 N_6 N_3 N_12 GND mn15  l=0.13u w=0.46u m=1
M11 N_28 N_18 N_30 GND mn15  l=0.13u w=0.17u m=1
M12 N_28 RN GND GND mn15  l=0.13u w=0.42u m=1
M13 N_28 RN GND GND mn15  l=0.13u w=0.42u m=1
M14 Q N_12 GND GND mn15  l=0.13u w=0.46u m=1
M15 Q N_12 GND GND mn15  l=0.13u w=0.46u m=1
M16 Q N_12 GND GND mn15  l=0.13u w=0.46u m=1
M17 GND N_12 N_18 GND mn15  l=0.13u w=0.17u m=1
M18 N_4 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_3 N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
M20 N_8 D VDD VDD mp15  l=0.13u w=0.42u m=1
M21 N_21 N_8 VDD VDD mp15  l=0.13u w=0.51u m=1
M22 N_21 N_3 N_9 VDD mp15  l=0.13u w=0.51u m=1
M23 N_22 N_6 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 N_6 N_9 VDD VDD mp15  l=0.13u w=0.35u m=1
M25 VDD N_9 N_6 VDD mp15  l=0.13u w=0.35u m=1
M26 N_22 N_4 N_9 VDD mp15  l=0.13u w=0.17u m=1
M27 N_6 N_4 N_12 VDD mp15  l=0.13u w=0.35u m=1
M28 N_12 N_4 N_6 VDD mp15  l=0.13u w=0.35u m=1
M29 N_23 N_3 N_12 VDD mp15  l=0.13u w=0.17u m=1
M30 N_23 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M31 N_12 RN VDD VDD mp15  l=0.13u w=0.72u m=1
M32 Q N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M33 Q N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M34 Q N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_12 N_18 VDD mp15  l=0.13u w=0.17u m=1
.ends dfcrq3
* SPICE INPUT		Tue Jul 31 19:17:50 2018	dfcrqm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfcrqm
.subckt dfcrqm VDD Q GND RN D CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.2u m=1
M2 GND N_4 N_3 GND mn15  l=0.13u w=0.17u m=1
M3 N_31 RN GND GND mn15  l=0.13u w=0.29u m=1
M4 N_28 RN GND GND mn15  l=0.13u w=0.17u m=1
M5 GND D N_7 GND mn15  l=0.13u w=0.175u m=1
M6 N_29 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M7 N_30 N_3 N_9 GND mn15  l=0.13u w=0.17u m=1
M8 N_30 N_6 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_31 N_9 N_6 GND mn15  l=0.13u w=0.29u m=1
M10 N_32 N_17 N_28 GND mn15  l=0.13u w=0.17u m=1
M11 N_29 N_4 N_9 GND mn15  l=0.13u w=0.28u m=1
M12 N_32 N_4 N_12 GND mn15  l=0.13u w=0.17u m=1
M13 N_12 N_3 N_6 GND mn15  l=0.13u w=0.28u m=1
M14 Q N_12 GND GND mn15  l=0.13u w=0.36u m=1
M15 N_17 N_12 GND GND mn15  l=0.13u w=0.28u m=1
M16 N_4 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M17 N_3 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M18 VDD RN N_6 VDD mp15  l=0.13u w=0.33u m=1
M19 VDD D N_7 VDD mp15  l=0.13u w=0.28u m=1
M20 N_18 N_7 VDD VDD mp15  l=0.13u w=0.37u m=1
M21 N_18 N_3 N_9 VDD mp15  l=0.13u w=0.37u m=1
M22 N_19 N_6 VDD VDD mp15  l=0.13u w=0.17u m=1
M23 N_6 N_9 VDD VDD mp15  l=0.13u w=0.33u m=1
M24 N_19 N_4 N_9 VDD mp15  l=0.13u w=0.17u m=1
M25 N_12 RN VDD VDD mp15  l=0.13u w=0.28u m=1
M26 N_20 N_17 VDD VDD mp15  l=0.13u w=0.28u m=1
M27 N_6 N_4 N_12 VDD mp15  l=0.13u w=0.37u m=1
M28 N_20 N_3 N_12 VDD mp15  l=0.13u w=0.28u m=1
M29 Q N_12 VDD VDD mp15  l=0.13u w=0.55u m=1
M30 N_17 N_12 VDD VDD mp15  l=0.13u w=0.28u m=1
.ends dfcrqm
* SPICE INPUT		Tue Jul 31 19:18:03 2018	dfnfb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb0
.subckt dfnfb0 VDD QN Q GND D CKN
M1 GND CKN N_5 GND mn15  l=0.13u w=0.17u m=1
M2 N_26 D GND GND mn15  l=0.13u w=0.18u m=1
M3 N_26 N_9 N_6 GND mn15  l=0.13u w=0.18u m=1
M4 N_27 N_2 GND GND mn15  l=0.13u w=0.17u m=1
M5 GND N_6 N_2 GND mn15  l=0.13u w=0.18u m=1
M6 N_27 N_5 N_6 GND mn15  l=0.13u w=0.17u m=1
M7 N_28 N_2 GND GND mn15  l=0.13u w=0.18u m=1
M8 N_11 N_5 N_28 GND mn15  l=0.13u w=0.18u m=1
M9 GND N_5 N_9 GND mn15  l=0.13u w=0.17u m=1
M10 N_29 N_9 N_11 GND mn15  l=0.13u w=0.17u m=1
M11 QN N_14 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_29 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M13 Q N_11 GND GND mn15  l=0.13u w=0.26u m=1
M14 N_14 N_11 GND GND mn15  l=0.13u w=0.18u m=1
M15 N_5 CKN VDD VDD mp15  l=0.13u w=0.42u m=1
M16 N_15 D VDD VDD mp15  l=0.13u w=0.52u m=1
M17 N_15 N_5 N_6 VDD mp15  l=0.13u w=0.52u m=1
M18 N_16 N_9 N_6 VDD mp15  l=0.13u w=0.17u m=1
M19 N_16 N_2 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 VDD N_6 N_2 VDD mp15  l=0.13u w=0.26u m=1
M21 N_17 N_2 VDD VDD mp15  l=0.13u w=0.27u m=1
M22 N_17 N_9 N_11 VDD mp15  l=0.13u w=0.27u m=1
M23 VDD N_5 N_9 VDD mp15  l=0.13u w=0.42u m=1
M24 N_18 N_5 N_11 VDD mp15  l=0.13u w=0.17u m=1
M25 VDD N_14 QN VDD mp15  l=0.13u w=0.4u m=1
M26 N_18 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 Q N_11 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_14 N_11 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends dfnfb0
* SPICE INPUT		Tue Jul 31 19:18:17 2018	dfnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb1
.subckt dfnfb1 GND Q QN VDD D CKN
M1 GND CKN N_4 GND mn15  l=0.13u w=0.2u m=1
M2 N_15 D GND GND mn15  l=0.13u w=0.28u m=1
M3 N_15 N_12 N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_16 N_3 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_3 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M6 N_16 N_4 N_6 GND mn15  l=0.13u w=0.17u m=1
M7 Q N_14 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_9 N_14 GND GND mn15  l=0.13u w=0.28u m=1
M9 N_18 N_12 N_14 GND mn15  l=0.13u w=0.17u m=1
M10 N_17 N_4 N_14 GND mn15  l=0.13u w=0.36u m=1
M11 QN N_9 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_18 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M13 GND N_4 N_12 GND mn15  l=0.13u w=0.17u m=1
M14 N_17 N_3 GND GND mn15  l=0.13u w=0.36u m=1
M15 N_4 CKN VDD VDD mp15  l=0.13u w=0.51u m=1
M16 N_72 D VDD VDD mp15  l=0.13u w=0.42u m=1
M17 N_72 N_4 N_6 VDD mp15  l=0.13u w=0.42u m=1
M18 N_73 N_12 N_6 VDD mp15  l=0.13u w=0.17u m=1
M19 N_73 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 N_3 N_6 VDD VDD mp15  l=0.13u w=0.39u m=1
M21 N_75 N_4 N_14 VDD mp15  l=0.13u w=0.17u m=1
M22 QN N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_75 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 VDD N_4 N_12 VDD mp15  l=0.13u w=0.42u m=1
M25 N_74 N_3 VDD VDD mp15  l=0.13u w=0.57u m=1
M26 N_74 N_12 N_14 VDD mp15  l=0.13u w=0.57u m=1
M27 Q N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 N_9 N_14 VDD VDD mp15  l=0.13u w=0.41u m=1
.ends dfnfb1
* SPICE INPUT		Tue Jul 31 19:18:30 2018	dfnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfb2
.subckt dfnfb2 GND QN Q VDD D CKN
M1 GND CKN N_4 GND mn15  l=0.13u w=0.27u m=1
M2 N_17 D GND GND mn15  l=0.13u w=0.41u m=1
M3 N_17 N_9 N_6 GND mn15  l=0.13u w=0.41u m=1
M4 N_18 N_4 N_6 GND mn15  l=0.13u w=0.17u m=1
M5 N_18 N_2 GND GND mn15  l=0.13u w=0.17u m=1
M6 GND N_6 N_2 GND mn15  l=0.13u w=0.41u m=1
M7 GND N_4 N_9 GND mn15  l=0.13u w=0.22u m=1
M8 N_19 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M9 N_19 N_4 N_11 GND mn15  l=0.13u w=0.46u m=1
M10 N_20 N_9 N_11 GND mn15  l=0.13u w=0.17u m=1
M11 GND N_15 QN GND mn15  l=0.13u w=0.46u m=1
M12 GND N_15 QN GND mn15  l=0.13u w=0.46u m=1
M13 N_20 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M14 GND N_11 Q GND mn15  l=0.13u w=0.46u m=1
M15 GND N_11 Q GND mn15  l=0.13u w=0.46u m=1
M16 GND N_11 N_15 GND mn15  l=0.13u w=0.36u m=1
M17 N_4 CKN VDD VDD mp15  l=0.13u w=0.67u m=1
M18 N_79 D VDD VDD mp15  l=0.13u w=0.63u m=1
M19 N_79 N_4 N_6 VDD mp15  l=0.13u w=0.63u m=1
M20 N_80 N_9 N_6 VDD mp15  l=0.13u w=0.17u m=1
M21 N_80 N_2 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_2 N_6 VDD VDD mp15  l=0.13u w=0.63u m=1
M23 VDD N_4 N_9 VDD mp15  l=0.13u w=0.55u m=1
M24 N_81 N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_81 N_9 N_11 VDD mp15  l=0.13u w=0.69u m=1
M26 N_82 N_4 N_11 VDD mp15  l=0.13u w=0.17u m=1
M27 QN N_15 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_15 QN VDD mp15  l=0.13u w=0.69u m=1
M29 N_82 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 VDD N_11 Q VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_11 Q VDD mp15  l=0.13u w=0.69u m=1
M32 N_15 N_11 VDD VDD mp15  l=0.13u w=0.53u m=1
.ends dfnfb2
* SPICE INPUT		Tue Jul 31 19:18:41 2018	dfnfq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfq0
.subckt dfnfq0 VDD Q GND CKN D
M1 Q N_8 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 N_8 GND GND mn15  l=0.13u w=0.18u m=1
M3 N_8 N_6 N_25 GND mn15  l=0.13u w=0.17u m=1
M4 N_26 N_11 N_8 GND mn15  l=0.13u w=0.18u m=1
M5 GND N_11 N_6 GND mn15  l=0.13u w=0.17u m=1
M6 N_26 N_10 GND GND mn15  l=0.13u w=0.18u m=1
M7 N_25 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_28 N_11 N_13 GND mn15  l=0.13u w=0.17u m=1
M9 GND N_13 N_10 GND mn15  l=0.13u w=0.18u m=1
M10 N_28 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_27 N_6 N_13 GND mn15  l=0.13u w=0.18u m=1
M12 N_27 D GND GND mn15  l=0.13u w=0.18u m=1
M13 GND CKN N_11 GND mn15  l=0.13u w=0.17u m=1
M14 Q N_8 VDD VDD mp15  l=0.13u w=0.4u m=1
M15 N_4 N_8 VDD VDD mp15  l=0.13u w=0.26u m=1
M16 VDD N_11 N_6 VDD mp15  l=0.13u w=0.42u m=1
M17 N_8 N_11 N_14 VDD mp15  l=0.13u w=0.17u m=1
M18 N_15 N_6 N_8 VDD mp15  l=0.13u w=0.27u m=1
M19 N_15 N_10 VDD VDD mp15  l=0.13u w=0.27u m=1
M20 N_14 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M21 N_10 N_13 VDD VDD mp15  l=0.13u w=0.26u m=1
M22 N_17 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M23 N_17 N_6 N_13 VDD mp15  l=0.13u w=0.17u m=1
M24 N_16 N_11 N_13 VDD mp15  l=0.13u w=0.52u m=1
M25 N_16 D VDD VDD mp15  l=0.13u w=0.52u m=1
M26 VDD CKN N_11 VDD mp15  l=0.13u w=0.42u m=1
.ends dfnfq0
* SPICE INPUT		Tue Jul 31 19:18:54 2018	dfnfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfq1
.subckt dfnfq1 GND Q D CKN VDD
M1 Q N_13 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 N_13 GND GND mn15  l=0.13u w=0.27u m=1
M3 GND CKN N_7 GND mn15  l=0.13u w=0.19u m=1
M4 N_14 D GND GND mn15  l=0.13u w=0.27u m=1
M5 N_15 N_7 N_9 GND mn15  l=0.13u w=0.17u m=1
M6 N_14 N_11 N_9 GND mn15  l=0.13u w=0.27u m=1
M7 N_6 N_9 GND GND mn15  l=0.13u w=0.27u m=1
M8 N_15 N_6 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_17 N_6 GND GND mn15  l=0.13u w=0.36u m=1
M10 GND N_7 N_11 GND mn15  l=0.13u w=0.16u m=1
M11 N_17 N_7 N_13 GND mn15  l=0.13u w=0.36u m=1
M12 N_13 N_11 N_16 GND mn15  l=0.13u w=0.17u m=1
M13 N_16 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M14 Q N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_4 N_13 VDD VDD mp15  l=0.13u w=0.39u m=1
M16 N_7 CKN VDD VDD mp15  l=0.13u w=0.49u m=1
M17 N_30 D VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_30 N_7 N_9 VDD mp15  l=0.13u w=0.4u m=1
M19 N_31 N_11 N_9 VDD mp15  l=0.13u w=0.17u m=1
M20 VDD N_9 N_6 VDD mp15  l=0.13u w=0.37u m=1
M21 N_31 N_6 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_32 N_6 VDD VDD mp15  l=0.13u w=0.57u m=1
M23 VDD N_7 N_11 VDD mp15  l=0.13u w=0.4u m=1
M24 N_33 N_7 N_13 VDD mp15  l=0.13u w=0.17u m=1
M25 N_32 N_11 N_13 VDD mp15  l=0.13u w=0.57u m=1
M26 N_33 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
.ends dfnfq1
* SPICE INPUT		Tue Jul 31 19:19:09 2018	dfnfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnfq2
.subckt dfnfq2 VDD Q GND D CKN
M1 GND N_14 Q GND mn15  l=0.13u w=0.46u m=1
M2 GND N_14 Q GND mn15  l=0.13u w=0.46u m=1
M3 GND N_14 N_9 GND mn15  l=0.13u w=0.36u m=1
M4 GND CKN N_5 GND mn15  l=0.13u w=0.27u m=1
M5 N_26 D GND GND mn15  l=0.13u w=0.41u m=1
M6 N_26 N_12 N_6 GND mn15  l=0.13u w=0.41u m=1
M7 N_27 N_5 N_6 GND mn15  l=0.13u w=0.17u m=1
M8 N_27 N_3 GND GND mn15  l=0.13u w=0.17u m=1
M9 GND N_6 N_3 GND mn15  l=0.13u w=0.41u m=1
M10 N_28 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M11 GND N_5 N_12 GND mn15  l=0.13u w=0.22u m=1
M12 N_29 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_14 N_12 N_28 GND mn15  l=0.13u w=0.17u m=1
M14 N_29 N_5 N_14 GND mn15  l=0.13u w=0.46u m=1
M15 N_5 CKN VDD VDD mp15  l=0.13u w=0.67u m=1
M16 N_15 D VDD VDD mp15  l=0.13u w=0.63u m=1
M17 N_15 N_5 N_6 VDD mp15  l=0.13u w=0.63u m=1
M18 N_16 N_12 N_6 VDD mp15  l=0.13u w=0.17u m=1
M19 N_16 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 N_3 N_6 VDD VDD mp15  l=0.13u w=0.63u m=1
M21 VDD N_14 Q VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_14 Q VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_14 N_9 VDD mp15  l=0.13u w=0.53u m=1
M24 N_17 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M25 VDD N_5 N_12 VDD mp15  l=0.13u w=0.55u m=1
M26 N_18 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_18 N_12 N_14 VDD mp15  l=0.13u w=0.69u m=1
M28 N_14 N_5 N_17 VDD mp15  l=0.13u w=0.17u m=1
.ends dfnfq2
* SPICE INPUT		Tue Jul 31 19:19:23 2018	dfnrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb0
.subckt dfnrb0 GND Q QN CK D VDD
M1 Q N_9 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 N_9 GND GND mn15  l=0.13u w=0.18u m=1
M3 QN N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_16 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_16 N_11 N_9 GND mn15  l=0.13u w=0.17u m=1
M6 N_15 N_7 N_9 GND mn15  l=0.13u w=0.17u m=1
M7 N_15 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M8 GND N_11 N_7 GND mn15  l=0.13u w=0.17u m=1
M9 N_18 N_7 N_13 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_13 N_10 GND mn15  l=0.13u w=0.18u m=1
M11 GND CK N_11 GND mn15  l=0.13u w=0.17u m=1
M12 N_18 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M13 N_17 N_11 N_13 GND mn15  l=0.13u w=0.18u m=1
M14 N_17 D GND GND mn15  l=0.13u w=0.18u m=1
M15 Q N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_4 N_9 VDD VDD mp15  l=0.13u w=0.26u m=1
M17 QN N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_27 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 N_26 N_11 N_9 VDD mp15  l=0.13u w=0.27u m=1
M20 N_27 N_7 N_9 VDD mp15  l=0.13u w=0.17u m=1
M21 N_26 N_10 VDD VDD mp15  l=0.13u w=0.27u m=1
M22 N_7 N_11 VDD VDD mp15  l=0.13u w=0.42u m=1
M23 N_28 N_7 N_13 VDD mp15  l=0.13u w=0.52u m=1
M24 VDD N_13 N_10 VDD mp15  l=0.13u w=0.26u m=1
M25 N_29 N_11 N_13 VDD mp15  l=0.13u w=0.17u m=1
M26 N_11 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M27 N_29 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 N_28 D VDD VDD mp15  l=0.13u w=0.52u m=1
.ends dfnrb0
* SPICE INPUT		Tue Jul 31 19:19:39 2018	dfnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb1
.subckt dfnrb1 GND Q QN CK D VDD
M1 Q N_9 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M3 QN N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_16 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_16 N_11 N_9 GND mn15  l=0.13u w=0.17u m=1
M6 N_15 N_7 N_9 GND mn15  l=0.13u w=0.41u m=1
M7 N_15 N_10 GND GND mn15  l=0.13u w=0.41u m=1
M8 GND N_11 N_7 GND mn15  l=0.13u w=0.2u m=1
M9 N_18 N_7 N_13 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_13 N_10 GND mn15  l=0.13u w=0.28u m=1
M11 N_18 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_13 N_11 N_17 GND mn15  l=0.13u w=0.28u m=1
M13 N_17 D GND GND mn15  l=0.13u w=0.28u m=1
M14 GND CK N_11 GND mn15  l=0.13u w=0.2u m=1
M15 Q N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_4 N_9 VDD VDD mp15  l=0.13u w=0.41u m=1
M17 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_72 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 N_71 N_11 N_9 VDD mp15  l=0.13u w=0.62u m=1
M20 N_72 N_7 N_9 VDD mp15  l=0.13u w=0.17u m=1
M21 N_71 N_10 VDD VDD mp15  l=0.13u w=0.62u m=1
M22 VDD N_11 N_7 VDD mp15  l=0.13u w=0.51u m=1
M23 N_73 N_7 N_13 VDD mp15  l=0.13u w=0.42u m=1
M24 VDD N_13 N_10 VDD mp15  l=0.13u w=0.41u m=1
M25 N_74 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M26 N_74 N_11 N_13 VDD mp15  l=0.13u w=0.17u m=1
M27 N_73 D VDD VDD mp15  l=0.13u w=0.42u m=1
M28 N_11 CK VDD VDD mp15  l=0.13u w=0.51u m=1
.ends dfnrb1
* SPICE INPUT		Tue Jul 31 19:19:55 2018	dfnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrb2
.subckt dfnrb2 GND Q QN VDD D CK
M1 N_18 N_5 N_6 GND mn15  l=0.13u w=0.41u m=1
M2 N_19 N_14 N_6 GND mn15  l=0.13u w=0.17u m=1
M3 N_5 CK GND GND mn15  l=0.13u w=0.27u m=1
M4 N_3 N_6 GND GND mn15  l=0.13u w=0.205u m=1
M5 GND N_6 N_3 GND mn15  l=0.13u w=0.205u m=1
M6 N_18 D GND GND mn15  l=0.13u w=0.41u m=1
M7 N_19 N_3 GND GND mn15  l=0.13u w=0.17u m=1
M8 Q N_16 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_16 Q GND mn15  l=0.13u w=0.46u m=1
M10 GND N_16 N_10 GND mn15  l=0.13u w=0.37u m=1
M11 GND N_5 N_14 GND mn15  l=0.13u w=0.22u m=1
M12 N_20 N_3 GND GND mn15  l=0.13u w=0.41u m=1
M13 N_21 N_5 N_16 GND mn15  l=0.13u w=0.17u m=1
M14 N_20 N_14 N_16 GND mn15  l=0.13u w=0.41u m=1
M15 GND N_10 QN GND mn15  l=0.13u w=0.46u m=1
M16 GND N_10 QN GND mn15  l=0.13u w=0.46u m=1
M17 GND N_10 N_21 GND mn15  l=0.13u w=0.17u m=1
M18 N_33 N_14 N_6 VDD mp15  l=0.13u w=0.63u m=1
M19 N_34 N_5 N_6 VDD mp15  l=0.13u w=0.17u m=1
M20 N_5 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M21 N_3 N_6 VDD VDD mp15  l=0.13u w=0.315u m=1
M22 VDD N_6 N_3 VDD mp15  l=0.13u w=0.315u m=1
M23 N_33 D VDD VDD mp15  l=0.13u w=0.63u m=1
M24 N_34 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M25 VDD N_5 N_14 VDD mp15  l=0.13u w=0.55u m=1
M26 N_35 N_3 VDD VDD mp15  l=0.13u w=0.62u m=1
M27 N_35 N_5 N_16 VDD mp15  l=0.13u w=0.62u m=1
M28 VDD N_10 QN VDD mp15  l=0.13u w=0.69u m=1
M29 QN N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_10 N_36 VDD mp15  l=0.13u w=0.17u m=1
M31 N_36 N_14 N_16 VDD mp15  l=0.13u w=0.17u m=1
M32 VDD N_16 Q VDD mp15  l=0.13u w=0.69u m=1
M33 VDD N_16 Q VDD mp15  l=0.13u w=0.69u m=1
M34 N_10 N_16 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends dfnrb2
* SPICE INPUT		Tue Jul 31 19:20:13 2018	dfnrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq0
.subckt dfnrq0 VDD Q GND D CK
M1 GND N_6 N_2 GND mn15  l=0.13u w=0.18u m=1
M2 N_26 N_2 GND GND mn15  l=0.13u w=0.17u m=1
M3 N_26 N_9 N_6 GND mn15  l=0.13u w=0.17u m=1
M4 GND CK N_5 GND mn15  l=0.13u w=0.17u m=1
M5 N_25 D GND GND mn15  l=0.13u w=0.18u m=1
M6 N_25 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M7 N_27 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_10 N_5 N_27 GND mn15  l=0.13u w=0.17u m=1
M9 N_28 N_9 N_10 GND mn15  l=0.13u w=0.17u m=1
M10 N_28 N_2 GND GND mn15  l=0.13u w=0.17u m=1
M11 GND N_5 N_9 GND mn15  l=0.13u w=0.17u m=1
M12 Q N_10 GND GND mn15  l=0.13u w=0.26u m=1
M13 N_13 N_10 GND GND mn15  l=0.13u w=0.18u m=1
M14 VDD N_6 N_2 VDD mp15  l=0.13u w=0.26u m=1
M15 N_15 N_2 VDD VDD mp15  l=0.13u w=0.17u m=1
M16 N_14 N_9 N_6 VDD mp15  l=0.13u w=0.52u m=1
M17 N_5 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M18 N_14 D VDD VDD mp15  l=0.13u w=0.52u m=1
M19 N_15 N_5 N_6 VDD mp15  l=0.13u w=0.17u m=1
M20 N_16 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M21 N_10 N_9 N_16 VDD mp15  l=0.13u w=0.17u m=1
M22 N_10 N_5 N_17 VDD mp15  l=0.13u w=0.27u m=1
M23 N_17 N_2 VDD VDD mp15  l=0.13u w=0.27u m=1
M24 N_9 N_5 VDD VDD mp15  l=0.13u w=0.42u m=1
M25 Q N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M26 N_13 N_10 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends dfnrq0
* SPICE INPUT		Tue Jul 31 19:20:26 2018	dfnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq1
.subckt dfnrq1 GND Q VDD D CK
M1 GND CK N_3 GND mn15  l=0.13u w=0.2u m=1
M2 N_14 D GND GND mn15  l=0.13u w=0.28u m=1
M3 N_5 N_3 N_14 GND mn15  l=0.13u w=0.28u m=1
M4 N_15 N_2 GND GND mn15  l=0.13u w=0.17u m=1
M5 GND N_5 N_2 GND mn15  l=0.13u w=0.28u m=1
M6 N_15 N_8 N_5 GND mn15  l=0.13u w=0.17u m=1
M7 GND N_3 N_8 GND mn15  l=0.13u w=0.2u m=1
M8 N_17 N_2 GND GND mn15  l=0.13u w=0.36u m=1
M9 N_17 N_8 N_10 GND mn15  l=0.13u w=0.36u m=1
M10 N_10 N_3 N_16 GND mn15  l=0.13u w=0.17u m=1
M11 N_16 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M12 Q N_10 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_13 N_10 GND GND mn15  l=0.13u w=0.28u m=1
M14 N_3 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M15 N_29 D VDD VDD mp15  l=0.13u w=0.42u m=1
M16 N_30 N_3 N_5 VDD mp15  l=0.13u w=0.17u m=1
M17 N_30 N_2 VDD VDD mp15  l=0.13u w=0.17u m=1
M18 VDD N_5 N_2 VDD mp15  l=0.13u w=0.41u m=1
M19 N_29 N_8 N_5 VDD mp15  l=0.13u w=0.42u m=1
M20 VDD N_3 N_8 VDD mp15  l=0.13u w=0.51u m=1
M21 N_32 N_2 VDD VDD mp15  l=0.13u w=0.52u m=1
M22 N_32 N_3 N_10 VDD mp15  l=0.13u w=0.52u m=1
M23 N_10 N_8 N_31 VDD mp15  l=0.13u w=0.17u m=1
M24 N_31 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M25 Q N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_13 N_10 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends dfnrq1
* SPICE INPUT		Tue Jul 31 19:20:39 2018	dfnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfnrq2
.subckt dfnrq2 VDD Q GND D CK
M1 N_27 N_12 N_6 GND mn15  l=0.13u w=0.17u m=1
M2 GND N_3 N_27 GND mn15  l=0.13u w=0.17u m=1
M3 Q N_6 GND GND mn15  l=0.13u w=0.46u m=1
M4 Q N_6 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 N_6 GND GND mn15  l=0.13u w=0.36u m=1
M6 GND N_12 N_4 GND mn15  l=0.13u w=0.22u m=1
M7 N_26 N_4 N_6 GND mn15  l=0.13u w=0.41u m=1
M8 N_26 N_10 GND GND mn15  l=0.13u w=0.41u m=1
M9 N_12 CK GND GND mn15  l=0.13u w=0.27u m=1
M10 N_28 D GND GND mn15  l=0.13u w=0.41u m=1
M11 N_28 N_12 N_13 GND mn15  l=0.13u w=0.41u m=1
M12 N_29 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M13 N_10 N_13 GND GND mn15  l=0.13u w=0.205u m=1
M14 GND N_13 N_10 GND mn15  l=0.13u w=0.205u m=1
M15 N_29 N_4 N_13 GND mn15  l=0.13u w=0.17u m=1
M16 N_16 N_4 N_6 VDD mp15  l=0.13u w=0.17u m=1
M17 N_15 N_12 N_6 VDD mp15  l=0.13u w=0.62u m=1
M18 VDD N_3 N_16 VDD mp15  l=0.13u w=0.17u m=1
M19 N_3 N_6 VDD VDD mp15  l=0.13u w=0.53u m=1
M20 Q N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 Q N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_12 N_4 VDD mp15  l=0.13u w=0.55u m=1
M23 N_15 N_10 VDD VDD mp15  l=0.13u w=0.62u m=1
M24 N_12 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M25 N_17 D VDD VDD mp15  l=0.13u w=0.63u m=1
M26 N_18 N_12 N_13 VDD mp15  l=0.13u w=0.17u m=1
M27 N_18 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 N_10 N_13 VDD VDD mp15  l=0.13u w=0.31u m=1
M29 VDD N_13 N_10 VDD mp15  l=0.13u w=0.32u m=1
M30 N_17 N_4 N_13 VDD mp15  l=0.13u w=0.63u m=1
.ends dfnrq2
* SPICE INPUT		Tue Jul 31 19:20:52 2018	dfpfb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb0
.subckt dfpfb0 VDD Q QN GND SN D CKN
M1 GND CKN N_4 GND mn15  l=0.13u w=0.17u m=1
M2 N_29 D GND GND mn15  l=0.13u w=0.26u m=1
M3 N_29 N_2 N_5 GND mn15  l=0.13u w=0.26u m=1
M4 GND N_9 N_30 GND mn15  l=0.13u w=0.17u m=1
M5 N_30 N_4 N_5 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M7 QN N_10 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_16 N_10 GND GND mn15  l=0.13u w=0.18u m=1
M9 N_9 N_5 N_26 GND mn15  l=0.13u w=0.31u m=1
M10 N_10 N_4 N_9 GND mn15  l=0.13u w=0.28u m=1
M11 N_31 N_16 N_26 GND mn15  l=0.13u w=0.17u m=1
M12 N_10 N_2 N_31 GND mn15  l=0.13u w=0.17u m=1
M13 N_26 SN GND GND mn15  l=0.13u w=0.37u m=1
M14 Q N_16 GND GND mn15  l=0.13u w=0.26u m=1
M15 N_4 CKN VDD VDD mp15  l=0.13u w=0.44u m=1
M16 N_17 D VDD VDD mp15  l=0.13u w=0.38u m=1
M17 N_18 N_2 N_5 VDD mp15  l=0.13u w=0.17u m=1
M18 N_18 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 VDD N_4 N_2 VDD mp15  l=0.13u w=0.42u m=1
M20 N_17 N_4 N_5 VDD mp15  l=0.13u w=0.38u m=1
M21 N_9 N_5 VDD VDD mp15  l=0.13u w=0.39u m=1
M22 N_10 N_4 N_19 VDD mp15  l=0.13u w=0.17u m=1
M23 N_19 N_16 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 N_10 N_2 N_9 VDD mp15  l=0.13u w=0.42u m=1
M25 N_10 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M26 Q N_16 VDD VDD mp15  l=0.13u w=0.4u m=1
M27 QN N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_16 N_10 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends dfpfb0
* SPICE INPUT		Tue Jul 31 19:21:05 2018	dfpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb1
.subckt dfpfb1 GND Q QN VDD SN D CKN
M1 GND CKN N_3 GND mn15  l=0.13u w=0.2u m=1
M2 N_17 D GND GND mn15  l=0.13u w=0.28u m=1
M3 N_17 N_2 N_5 GND mn15  l=0.13u w=0.28u m=1
M4 GND N_9 N_18 GND mn15  l=0.13u w=0.17u m=1
M5 N_18 N_3 N_5 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_3 N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_9 N_5 N_7 GND mn15  l=0.13u w=0.4u m=1
M8 N_10 N_3 N_9 GND mn15  l=0.13u w=0.36u m=1
M9 N_19 N_16 N_7 GND mn15  l=0.13u w=0.17u m=1
M10 N_10 N_2 N_19 GND mn15  l=0.13u w=0.17u m=1
M11 N_7 SN GND GND mn15  l=0.13u w=0.46u m=1
M12 Q N_16 GND GND mn15  l=0.13u w=0.46u m=1
M13 QN N_10 GND GND mn15  l=0.13u w=0.46u m=1
M14 N_16 N_10 GND GND mn15  l=0.13u w=0.28u m=1
M15 N_3 CKN VDD VDD mp15  l=0.13u w=0.51u m=1
M16 N_31 D VDD VDD mp15  l=0.13u w=0.42u m=1
M17 N_32 N_2 N_5 VDD mp15  l=0.13u w=0.17u m=1
M18 N_32 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 N_31 N_3 N_5 VDD mp15  l=0.13u w=0.42u m=1
M20 VDD N_3 N_2 VDD mp15  l=0.13u w=0.51u m=1
M21 N_9 N_5 VDD VDD mp15  l=0.13u w=0.25u m=1
M22 VDD N_5 N_9 VDD mp15  l=0.13u w=0.25u m=1
M23 N_10 N_3 N_33 VDD mp15  l=0.13u w=0.17u m=1
M24 N_33 N_16 VDD VDD mp15  l=0.13u w=0.17u m=1
M25 N_10 N_2 N_9 VDD mp15  l=0.13u w=0.565u m=1
M26 N_10 SN VDD VDD mp15  l=0.13u w=0.35u m=1
M27 Q N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 QN N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 N_16 N_10 VDD VDD mp15  l=0.13u w=0.41u m=1
.ends dfpfb1
* SPICE INPUT		Tue Jul 31 19:21:18 2018	dfpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfpfb2
.subckt dfpfb2 GND Q QN VDD SN D CKN
M1 N_4 CKN GND GND mn15  l=0.13u w=0.27u m=1
M2 N_20 D GND GND mn15  l=0.13u w=0.36u m=1
M3 N_21 N_4 N_5 GND mn15  l=0.13u w=0.17u m=1
M4 GND N_4 N_2 GND mn15  l=0.13u w=0.22u m=1
M5 N_20 N_2 N_5 GND mn15  l=0.13u w=0.36u m=1
M6 GND N_9 N_21 GND mn15  l=0.13u w=0.17u m=1
M7 N_9 N_5 N_7 GND mn15  l=0.13u w=0.46u m=1
M8 N_10 N_4 N_9 GND mn15  l=0.13u w=0.46u m=1
M9 N_22 N_16 N_7 GND mn15  l=0.13u w=0.17u m=1
M10 N_10 N_2 N_22 GND mn15  l=0.13u w=0.17u m=1
M11 GND SN N_7 GND mn15  l=0.13u w=0.46u m=1
M12 GND SN N_7 GND mn15  l=0.13u w=0.46u m=1
M13 GND N_10 QN GND mn15  l=0.13u w=0.46u m=1
M14 QN N_10 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_10 N_16 GND mn15  l=0.13u w=0.37u m=1
M16 GND N_16 Q GND mn15  l=0.13u w=0.46u m=1
M17 GND N_16 Q GND mn15  l=0.13u w=0.46u m=1
M18 N_4 CKN VDD VDD mp15  l=0.13u w=0.67u m=1
M19 N_33 D VDD VDD mp15  l=0.13u w=0.55u m=1
M20 VDD N_4 N_2 VDD mp15  l=0.13u w=0.55u m=1
M21 N_33 N_4 N_5 VDD mp15  l=0.13u w=0.55u m=1
M22 N_34 N_2 N_5 VDD mp15  l=0.13u w=0.17u m=1
M23 N_34 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 VDD N_5 N_9 VDD mp15  l=0.13u w=0.405u m=1
M25 VDD N_5 N_9 VDD mp15  l=0.13u w=0.405u m=1
M26 N_10 N_4 N_35 VDD mp15  l=0.13u w=0.17u m=1
M27 N_35 N_16 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 N_10 N_2 N_9 VDD mp15  l=0.13u w=0.565u m=1
M29 N_10 SN VDD VDD mp15  l=0.13u w=0.56u m=1
M30 QN N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 QN N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 N_16 N_10 VDD VDD mp15  l=0.13u w=0.55u m=1
M33 VDD N_16 Q VDD mp15  l=0.13u w=0.69u m=1
M34 VDD N_16 Q VDD mp15  l=0.13u w=0.69u m=1
.ends dfpfb2
* SPICE INPUT		Tue Jul 31 19:21:31 2018	dfprb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb0
.subckt dfprb0 VDD Q QN GND SN D CK
M1 GND CK N_5 GND mn15  l=0.13u w=0.2u m=1
M2 N_30 D GND GND mn15  l=0.13u w=0.18u m=1
M3 N_30 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M4 N_31 N_8 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_31 N_2 N_6 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_5 N_2 GND mn15  l=0.13u w=0.17u m=1
M7 N_8 N_6 N_26 GND mn15  l=0.13u w=0.16u m=1
M8 N_26 N_6 N_8 GND mn15  l=0.13u w=0.15u m=1
M9 N_8 N_2 N_10 GND mn15  l=0.13u w=0.3u m=1
M10 N_32 N_17 N_26 GND mn15  l=0.13u w=0.17u m=1
M11 N_10 N_5 N_32 GND mn15  l=0.13u w=0.17u m=1
M12 Q N_17 GND GND mn15  l=0.13u w=0.26u m=1
M13 N_26 SN GND GND mn15  l=0.13u w=0.31u m=1
M14 QN N_10 GND GND mn15  l=0.13u w=0.26u m=1
M15 N_17 N_10 GND GND mn15  l=0.13u w=0.18u m=1
M16 N_5 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M17 N_18 D VDD VDD mp15  l=0.13u w=0.28u m=1
M18 N_19 N_8 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 N_18 N_2 N_6 VDD mp15  l=0.13u w=0.28u m=1
M20 VDD N_5 N_2 VDD mp15  l=0.13u w=0.42u m=1
M21 N_19 N_5 N_6 VDD mp15  l=0.13u w=0.17u m=1
M22 N_8 N_6 VDD VDD mp15  l=0.13u w=0.2u m=1
M23 VDD N_6 N_8 VDD mp15  l=0.13u w=0.18u m=1
M24 N_20 N_2 N_10 VDD mp15  l=0.13u w=0.17u m=1
M25 N_20 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M26 N_8 N_5 N_10 VDD mp15  l=0.13u w=0.39u m=1
M27 VDD N_17 Q VDD mp15  l=0.13u w=0.4u m=1
M28 N_10 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M29 QN N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M30 N_17 N_10 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends dfprb0
* SPICE INPUT		Tue Jul 31 19:21:45 2018	dfprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb1
.subckt dfprb1 GND QN Q VDD SN D CK
M1 QN N_9 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_5 N_14 N_6 GND mn15  l=0.13u w=0.21u m=1
M4 N_6 N_14 N_5 GND mn15  l=0.13u w=0.21u m=1
M5 N_9 N_12 N_19 GND mn15  l=0.13u w=0.17u m=1
M6 N_19 N_4 N_5 GND mn15  l=0.13u w=0.17u m=1
M7 N_9 N_10 N_6 GND mn15  l=0.13u w=0.4u m=1
M8 GND CK N_12 GND mn15  l=0.13u w=0.2u m=1
M9 GND N_12 N_10 GND mn15  l=0.13u w=0.17u m=1
M10 N_20 D GND GND mn15  l=0.13u w=0.28u m=1
M11 N_21 N_6 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_20 N_12 N_14 GND mn15  l=0.13u w=0.28u m=1
M13 N_21 N_10 N_14 GND mn15  l=0.13u w=0.17u m=1
M14 N_5 SN GND GND mn15  l=0.13u w=0.32u m=1
M15 N_5 SN GND GND mn15  l=0.13u w=0.32u m=1
M16 Q N_4 GND GND mn15  l=0.13u w=0.46u m=1
M17 N_6 N_14 VDD VDD mp15  l=0.13u w=0.225u m=1
M18 VDD N_14 N_6 VDD mp15  l=0.13u w=0.225u m=1
M19 N_9 N_12 N_6 VDD mp15  l=0.13u w=0.565u m=1
M20 N_33 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M21 N_33 N_10 N_9 VDD mp15  l=0.13u w=0.17u m=1
M22 QN N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_4 N_9 VDD VDD mp15  l=0.13u w=0.41u m=1
M24 N_12 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M25 VDD N_12 N_10 VDD mp15  l=0.13u w=0.42u m=1
M26 N_35 N_12 N_14 VDD mp15  l=0.13u w=0.17u m=1
M27 N_34 D VDD VDD mp15  l=0.13u w=0.42u m=1
M28 N_35 N_6 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_34 N_10 N_14 VDD mp15  l=0.13u w=0.42u m=1
M30 N_9 SN VDD VDD mp15  l=0.13u w=0.37u m=1
M31 Q N_4 VDD VDD mp15  l=0.13u w=0.35u m=1
M32 VDD N_4 Q VDD mp15  l=0.13u w=0.35u m=1
.ends dfprb1
* SPICE INPUT		Tue Jul 31 19:21:58 2018	dfprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprb2
.subckt dfprb2 VDD Q QN GND SN D CK
M1 GND N_11 QN GND mn15  l=0.13u w=0.46u m=1
M2 GND N_11 QN GND mn15  l=0.13u w=0.46u m=1
M3 GND N_11 N_20 GND mn15  l=0.13u w=0.37u m=1
M4 N_33 D GND GND mn15  l=0.13u w=0.43u m=1
M5 N_33 N_4 N_5 GND mn15  l=0.13u w=0.43u m=1
M6 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M7 N_4 CK GND GND mn15  l=0.13u w=0.27u m=1
M8 N_34 N_2 N_5 GND mn15  l=0.13u w=0.17u m=1
M9 N_34 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M10 N_30 N_5 N_9 GND mn15  l=0.13u w=0.215u m=1
M11 N_9 N_5 N_30 GND mn15  l=0.13u w=0.215u m=1
M12 N_9 N_5 N_30 GND mn15  l=0.13u w=0.2u m=1
M13 N_35 N_4 N_11 GND mn15  l=0.13u w=0.17u m=1
M14 N_30 N_20 N_35 GND mn15  l=0.13u w=0.17u m=1
M15 GND SN N_30 GND mn15  l=0.13u w=0.31u m=1
M16 N_30 SN GND GND mn15  l=0.13u w=0.31u m=1
M17 N_30 SN GND GND mn15  l=0.13u w=0.3u m=1
M18 N_11 N_2 N_9 GND mn15  l=0.13u w=0.46u m=1
M19 GND N_20 Q GND mn15  l=0.13u w=0.46u m=1
M20 GND N_20 Q GND mn15  l=0.13u w=0.46u m=1
M21 N_21 D VDD VDD mp15  l=0.13u w=0.64u m=1
M22 VDD N_4 N_2 VDD mp15  l=0.13u w=0.42u m=1
M23 N_22 N_4 N_5 VDD mp15  l=0.13u w=0.17u m=1
M24 N_21 N_2 N_5 VDD mp15  l=0.13u w=0.64u m=1
M25 N_4 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M26 VDD N_9 N_22 VDD mp15  l=0.13u w=0.17u m=1
M27 N_9 N_5 VDD VDD mp15  l=0.13u w=0.325u m=1
M28 N_9 N_5 VDD VDD mp15  l=0.13u w=0.325u m=1
M29 N_11 N_4 N_9 VDD mp15  l=0.13u w=0.565u m=1
M30 N_23 N_2 N_11 VDD mp15  l=0.13u w=0.17u m=1
M31 N_23 N_20 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_11 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M33 N_11 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M34 Q N_20 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_20 Q VDD mp15  l=0.13u w=0.69u m=1
M36 VDD N_11 QN VDD mp15  l=0.13u w=0.69u m=1
M37 VDD N_11 QN VDD mp15  l=0.13u w=0.69u m=1
M38 N_20 N_11 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends dfprb2
* SPICE INPUT		Tue Jul 31 19:22:11 2018	dfprq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq0
.subckt dfprq0 VDD Q GND SN D CK
M1 Q N_13 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M3 N_7 CK GND GND mn15  l=0.13u w=0.18u m=1
M4 GND N_7 N_6 GND mn15  l=0.13u w=0.17u m=1
M5 GND D N_16 GND mn15  l=0.13u w=0.17u m=1
M6 N_77 N_16 GND GND mn15  l=0.13u w=0.17u m=1
M7 N_78 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_13 N_6 N_10 GND mn15  l=0.13u w=0.22u m=1
M9 N_78 N_6 N_18 GND mn15  l=0.13u w=0.17u m=1
M10 N_10 N_18 GND GND mn15  l=0.13u w=0.23u m=1
M11 N_77 N_7 N_18 GND mn15  l=0.13u w=0.17u m=1
M12 N_13 N_7 N_76 GND mn15  l=0.13u w=0.17u m=1
M13 N_76 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M14 N_13 N_9 GND GND mn15  l=0.13u w=0.18u m=1
M15 GND SN N_9 GND mn15  l=0.13u w=0.17u m=1
M16 Q N_13 VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_4 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M18 N_7 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M19 N_6 N_7 VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_10 N_18 N_11 VDD mp15  l=0.13u w=0.21u m=1
M21 N_11 N_18 N_10 VDD mp15  l=0.13u w=0.21u m=1
M22 N_13 N_7 N_10 VDD mp15  l=0.13u w=0.42u m=1
M23 N_22 N_6 N_13 VDD mp15  l=0.13u w=0.17u m=1
M24 N_11 N_4 N_22 VDD mp15  l=0.13u w=0.17u m=1
M25 N_11 N_9 VDD VDD mp15  l=0.13u w=0.57u m=1
M26 N_9 SN VDD VDD mp15  l=0.13u w=0.26u m=1
M27 VDD D N_16 VDD mp15  l=0.13u w=0.28u m=1
M28 N_24 N_16 VDD VDD mp15  l=0.13u w=0.36u m=1
M29 N_24 N_6 N_18 VDD mp15  l=0.13u w=0.36u m=1
M30 N_23 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M31 N_18 N_7 N_23 VDD mp15  l=0.13u w=0.17u m=1
.ends dfprq0
* SPICE INPUT		Tue Jul 31 19:22:26 2018	dfprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq1
.subckt dfprq1 GND Q VDD SN D CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.2u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 Q N_14 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_7 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M5 GND D N_9 GND mn15  l=0.13u w=0.175u m=1
M6 N_19 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M7 N_20 N_2 N_11 GND mn15  l=0.13u w=0.17u m=1
M8 N_20 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_14 N_2 N_13 GND mn15  l=0.13u w=0.255u m=1
M10 N_13 N_11 GND GND mn15  l=0.13u w=0.28u m=1
M11 N_19 N_4 N_11 GND mn15  l=0.13u w=0.28u m=1
M12 N_14 N_4 N_18 GND mn15  l=0.13u w=0.17u m=1
M13 N_18 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M14 GND SN N_15 GND mn15  l=0.13u w=0.18u m=1
M15 GND N_15 N_14 GND mn15  l=0.13u w=0.28u m=1
M16 N_4 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M17 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M18 Q N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_7 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 VDD D N_9 VDD mp15  l=0.13u w=0.28u m=1
M21 N_81 N_9 VDD VDD mp15  l=0.13u w=0.42u m=1
M22 N_11 N_2 N_81 VDD mp15  l=0.13u w=0.42u m=1
M23 N_80 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 N_11 N_4 N_80 VDD mp15  l=0.13u w=0.17u m=1
M25 N_26 N_11 N_13 VDD mp15  l=0.13u w=0.32u m=1
M26 N_26 N_11 N_13 VDD mp15  l=0.13u w=0.32u m=1
M27 N_14 N_4 N_13 VDD mp15  l=0.13u w=0.42u m=1
M28 N_82 N_2 N_14 VDD mp15  l=0.13u w=0.17u m=1
M29 N_26 N_7 N_82 VDD mp15  l=0.13u w=0.17u m=1
M30 N_15 SN VDD VDD mp15  l=0.13u w=0.26u m=1
M31 N_26 N_15 VDD VDD mp15  l=0.13u w=0.7u m=1
.ends dfprq1
* SPICE INPUT		Tue Jul 31 19:22:39 2018	dfprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprq2
.subckt dfprq2 GND Q SN VDD D CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.28u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.23u m=1
M3 N_8 D GND GND mn15  l=0.13u w=0.28u m=1
M4 N_21 N_8 GND GND mn15  l=0.13u w=0.36u m=1
M5 N_22 N_2 N_9 GND mn15  l=0.13u w=0.17u m=1
M6 N_22 N_6 GND GND mn15  l=0.13u w=0.17u m=1
M7 GND N_9 N_6 GND mn15  l=0.13u w=0.41u m=1
M8 N_9 N_4 N_21 GND mn15  l=0.13u w=0.36u m=1
M9 N_6 N_2 N_5 GND mn15  l=0.13u w=0.4u m=1
M10 N_5 N_4 N_11 GND mn15  l=0.13u w=0.17u m=1
M11 GND SN N_13 GND mn15  l=0.13u w=0.24u m=1
M12 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M14 GND N_5 N_15 GND mn15  l=0.13u w=0.17u m=1
M15 N_5 N_13 GND GND mn15  l=0.13u w=0.37u m=1
M16 N_11 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M17 N_4 CK VDD VDD mp15  l=0.13u w=0.66u m=1
M18 VDD N_4 N_2 VDD mp15  l=0.13u w=0.55u m=1
M19 N_13 SN VDD VDD mp15  l=0.13u w=0.34u m=1
M20 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_5 N_15 VDD mp15  l=0.13u w=0.17u m=1
M23 N_8 D VDD VDD mp15  l=0.13u w=0.42u m=1
M24 N_34 N_8 VDD VDD mp15  l=0.13u w=0.53u m=1
M25 N_34 N_2 N_9 VDD mp15  l=0.13u w=0.53u m=1
M26 N_33 N_6 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_9 N_4 N_33 VDD mp15  l=0.13u w=0.17u m=1
M28 N_27 N_13 VDD VDD mp15  l=0.13u w=0.61u m=1
M29 VDD N_13 N_27 VDD mp15  l=0.13u w=0.46u m=1
M30 N_6 N_9 N_27 VDD mp15  l=0.13u w=0.27u m=1
M31 N_6 N_9 N_27 VDD mp15  l=0.13u w=0.27u m=1
M32 N_6 N_9 N_27 VDD mp15  l=0.13u w=0.27u m=1
M33 N_6 N_9 N_27 VDD mp15  l=0.13u w=0.27u m=1
M34 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.59u m=1
M35 N_35 N_2 N_5 VDD mp15  l=0.13u w=0.17u m=1
M36 N_27 N_15 N_35 VDD mp15  l=0.13u w=0.17u m=1
.ends dfprq2
* SPICE INPUT		Tue Jul 31 19:22:52 2018	dfprqm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfprqm
.subckt dfprqm VDD Q GND SN D CK
M1 GND N_4 N_3 GND mn15  l=0.13u w=0.17u m=1
M2 N_4 CK GND GND mn15  l=0.13u w=0.18u m=1
M3 GND D N_6 GND mn15  l=0.13u w=0.175u m=1
M4 N_31 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M5 GND N_14 N_32 GND mn15  l=0.13u w=0.17u m=1
M6 N_14 N_8 GND GND mn15  l=0.13u w=0.28u m=1
M7 N_32 N_3 N_8 GND mn15  l=0.13u w=0.17u m=1
M8 N_17 N_3 N_14 GND mn15  l=0.13u w=0.28u m=1
M9 N_31 N_4 N_8 GND mn15  l=0.13u w=0.28u m=1
M10 N_17 N_4 N_30 GND mn15  l=0.13u w=0.17u m=1
M11 N_30 N_11 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_11 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M13 Q N_17 GND GND mn15  l=0.13u w=0.36u m=1
M14 GND SN N_12 GND mn15  l=0.13u w=0.17u m=1
M15 N_17 N_12 GND GND mn15  l=0.13u w=0.24u m=1
M16 N_3 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M17 N_4 CK VDD VDD mp15  l=0.13u w=0.45u m=1
M18 VDD D N_6 VDD mp15  l=0.13u w=0.28u m=1
M19 N_20 N_6 VDD VDD mp15  l=0.13u w=0.37u m=1
M20 N_8 N_3 N_20 VDD mp15  l=0.13u w=0.37u m=1
M21 N_19 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_8 N_4 N_19 VDD mp15  l=0.13u w=0.17u m=1
M23 Q N_17 VDD VDD mp15  l=0.13u w=0.55u m=1
M24 N_11 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M25 N_14 N_8 N_15 VDD mp15  l=0.13u w=0.21u m=1
M26 N_15 N_8 N_14 VDD mp15  l=0.13u w=0.21u m=1
M27 N_17 N_4 N_14 VDD mp15  l=0.13u w=0.39u m=1
M28 N_21 N_3 N_17 VDD mp15  l=0.13u w=0.17u m=1
M29 VDD SN N_12 VDD mp15  l=0.13u w=0.24u m=1
M30 N_15 N_11 N_21 VDD mp15  l=0.13u w=0.17u m=1
M31 N_15 N_12 VDD VDD mp15  l=0.13u w=0.59u m=1
.ends dfprqm
* SPICE INPUT		Tue Jul 31 19:23:04 2018	dfscrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfscrq0
.subckt dfscrq0 VDD Q GND RN D CK
M1 GND CK N_4 GND mn15  l=0.13u w=0.17u m=1
M2 N_25 D GND GND mn15  l=0.13u w=0.26u m=1
M3 N_3 RN N_25 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 N_4 N_3 GND mn15  l=0.13u w=0.28u m=1
M5 GND N_5 N_26 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_7 N_5 GND mn15  l=0.13u w=0.18u m=1
M7 N_26 N_11 N_7 GND mn15  l=0.13u w=0.17u m=1
M8 GND N_4 N_11 GND mn15  l=0.13u w=0.17u m=1
M9 N_27 N_5 GND GND mn15  l=0.13u w=0.17u m=1
M10 N_27 N_11 N_13 GND mn15  l=0.13u w=0.17u m=1
M11 N_28 N_4 N_13 GND mn15  l=0.13u w=0.17u m=1
M12 N_28 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M13 Q N_13 GND GND mn15  l=0.13u w=0.26u m=1
M14 N_14 N_13 GND GND mn15  l=0.13u w=0.18u m=1
M15 N_4 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M16 N_3 D VDD VDD mp15  l=0.13u w=0.35u m=1
M17 N_3 RN VDD VDD mp15  l=0.13u w=0.35u m=1
M18 N_15 N_4 N_7 VDD mp15  l=0.13u w=0.17u m=1
M19 N_15 N_5 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 VDD N_7 N_5 VDD mp15  l=0.13u w=0.26u m=1
M21 N_3 N_11 N_7 VDD mp15  l=0.13u w=0.42u m=1
M22 VDD N_4 N_11 VDD mp15  l=0.13u w=0.42u m=1
M23 N_16 N_5 VDD VDD mp15  l=0.13u w=0.27u m=1
M24 N_13 N_4 N_16 VDD mp15  l=0.13u w=0.27u m=1
M25 N_17 N_11 N_13 VDD mp15  l=0.13u w=0.17u m=1
M26 N_17 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 Q N_13 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_14 N_13 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends dfscrq0
* SPICE INPUT		Tue Jul 31 19:23:17 2018	dfscrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfscrq1
.subckt dfscrq1 GND Q VDD D RN CK
M1 GND CK N_3 GND mn15  l=0.13u w=0.2u m=1
M2 N_15 RN GND GND mn15  l=0.13u w=0.26u m=1
M3 N_5 D N_15 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 N_3 N_5 GND mn15  l=0.13u w=0.28u m=1
M5 GND N_2 N_16 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_6 N_2 GND mn15  l=0.13u w=0.28u m=1
M7 N_16 N_9 N_6 GND mn15  l=0.13u w=0.17u m=1
M8 GND N_3 N_9 GND mn15  l=0.13u w=0.2u m=1
M9 N_18 N_9 N_11 GND mn15  l=0.13u w=0.36u m=1
M10 N_11 N_3 N_17 GND mn15  l=0.13u w=0.17u m=1
M11 N_17 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_18 N_2 GND GND mn15  l=0.13u w=0.36u m=1
M13 Q N_11 GND GND mn15  l=0.13u w=0.46u m=1
M14 N_14 N_11 GND GND mn15  l=0.13u w=0.28u m=1
M15 N_3 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M16 VDD RN N_5 VDD mp15  l=0.13u w=0.35u m=1
M17 N_5 D VDD VDD mp15  l=0.13u w=0.35u m=1
M18 N_30 N_3 N_6 VDD mp15  l=0.13u w=0.17u m=1
M19 N_30 N_2 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 VDD N_6 N_2 VDD mp15  l=0.13u w=0.41u m=1
M21 N_6 N_9 N_5 VDD mp15  l=0.13u w=0.42u m=1
M22 VDD N_3 N_9 VDD mp15  l=0.13u w=0.51u m=1
M23 N_32 N_3 N_11 VDD mp15  l=0.13u w=0.52u m=1
M24 N_11 N_9 N_31 VDD mp15  l=0.13u w=0.17u m=1
M25 N_31 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M26 N_32 N_2 VDD VDD mp15  l=0.13u w=0.52u m=1
M27 Q N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 N_14 N_11 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends dfscrq1
* SPICE INPUT		Tue Jul 31 19:23:30 2018	dfscrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dfscrq2
.subckt dfscrq2 GND Q VDD CK RN D
M1 N_5 CK GND GND mn15  l=0.13u w=0.27u m=1
M2 N_16 RN GND GND mn15  l=0.13u w=0.46u m=1
M3 N_16 D N_6 GND mn15  l=0.13u w=0.46u m=1
M4 N_7 N_5 N_6 GND mn15  l=0.13u w=0.41u m=1
M5 GND N_3 N_17 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_7 N_3 GND mn15  l=0.13u w=0.205u m=1
M7 N_3 N_7 GND GND mn15  l=0.13u w=0.205u m=1
M8 N_17 N_11 N_7 GND mn15  l=0.13u w=0.17u m=1
M9 GND N_5 N_11 GND mn15  l=0.13u w=0.22u m=1
M10 N_18 N_11 N_13 GND mn15  l=0.13u w=0.41u m=1
M11 N_19 N_5 N_13 GND mn15  l=0.13u w=0.17u m=1
M12 GND N_10 N_19 GND mn15  l=0.13u w=0.17u m=1
M13 Q N_13 GND GND mn15  l=0.13u w=0.46u m=1
M14 Q N_13 GND GND mn15  l=0.13u w=0.46u m=1
M15 N_10 N_13 GND GND mn15  l=0.13u w=0.36u m=1
M16 N_18 N_3 GND GND mn15  l=0.13u w=0.41u m=1
M17 N_5 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M18 VDD RN N_6 VDD mp15  l=0.13u w=0.61u m=1
M19 N_6 D VDD VDD mp15  l=0.13u w=0.61u m=1
M20 N_31 N_5 N_7 VDD mp15  l=0.13u w=0.17u m=1
M21 N_31 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_3 N_7 VDD VDD mp15  l=0.13u w=0.31u m=1
M23 N_3 N_7 VDD VDD mp15  l=0.13u w=0.32u m=1
M24 N_7 N_11 N_6 VDD mp15  l=0.13u w=0.63u m=1
M25 N_11 N_5 VDD VDD mp15  l=0.13u w=0.55u m=1
M26 N_33 N_11 N_13 VDD mp15  l=0.13u w=0.17u m=1
M27 N_32 N_5 N_13 VDD mp15  l=0.13u w=0.62u m=1
M28 VDD N_10 N_33 VDD mp15  l=0.13u w=0.17u m=1
M29 Q N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 Q N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 N_10 N_13 VDD VDD mp15  l=0.13u w=0.53u m=1
M32 N_32 N_3 VDD VDD mp15  l=0.13u w=0.62u m=1
.ends dfscrq2
* SPICE INPUT		Tue Jul 31 19:23:44 2018	dl01d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d1
.subckt dl01d1 VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.14u m=1
M2 GND N_4 N_3 GND mn15  l=0.13u w=0.14u m=1
M3 N_7 N_3 GND GND mn15  l=0.13u w=0.14u m=1
M4 GND N_7 Y GND mn15  l=0.13u w=0.2u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.49u m=1
M6 N_3 N_4 VDD VDD mp15  l=0.13u w=0.49u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.13u w=0.49u m=1
M8 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends dl01d1
* SPICE INPUT		Tue Jul 31 19:23:56 2018	dl01d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01d2
.subckt dl01d2 Y VDD GND A
M1 N_8 A GND GND mn15  l=0.13u w=0.14u m=1
M2 GND N_8 N_7 GND mn15  l=0.13u w=0.14u m=1
M3 GND N_7 N_4 GND mn15  l=0.13u w=0.14u m=1
M4 Y N_4 GND GND mn15  l=0.13u w=0.24u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.24u m=1
M6 VDD N_7 N_4 VDD mp15  l=0.13u w=0.49u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_8 A VDD VDD mp15  l=0.13u w=0.49u m=1
M10 N_7 N_8 VDD VDD mp15  l=0.13u w=0.49u m=1
.ends dl01d2
* SPICE INPUT		Tue Jul 31 19:24:09 2018	dl01dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl01dm
.subckt dl01dm VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.14u m=1
M2 GND N_4 N_3 GND mn15  l=0.13u w=0.14u m=1
M3 N_7 N_3 GND GND mn15  l=0.13u w=0.14u m=1
M4 GND N_7 Y GND mn15  l=0.13u w=0.18u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.49u m=1
M6 N_3 N_4 VDD VDD mp15  l=0.13u w=0.49u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.13u w=0.49u m=1
M8 Y N_7 VDD VDD mp15  l=0.13u w=0.63u m=1
.ends dl01dm
* SPICE INPUT		Tue Jul 31 19:24:22 2018	dl02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d1
.subckt dl02d1 VDD Y GND A
M1 N_4 A GND GND mn15  l=0.13u w=0.14u m=1
M2 GND N_4 N_3 GND mn15  l=0.26u w=0.14u m=1
M3 N_7 N_3 GND GND mn15  l=0.26u w=0.14u m=1
M4 GND N_7 Y GND mn15  l=0.13u w=0.2u m=1
M5 N_4 A VDD VDD mp15  l=0.13u w=0.49u m=1
M6 N_3 N_4 VDD VDD mp15  l=0.26u w=0.49u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.26u w=0.49u m=1
M8 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends dl02d1
* SPICE INPUT		Tue Jul 31 19:24:35 2018	dl02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dl02d2
.subckt dl02d2 VDD Y GND A
M1 GND N_3 N_7 GND mn15  l=0.26u w=0.14u m=1
M2 GND N_7 Y GND mn15  l=0.13u w=0.34u m=1
M3 GND N_7 Y GND mn15  l=0.13u w=0.14u m=1
M4 N_4 A GND GND mn15  l=0.13u w=0.14u m=1
M5 GND N_4 N_3 GND mn15  l=0.26u w=0.14u m=1
M6 N_4 A VDD VDD mp15  l=0.13u w=0.49u m=1
M7 N_3 N_4 VDD VDD mp15  l=0.26u w=0.49u m=1
M8 VDD N_3 N_7 VDD mp15  l=0.26u w=0.49u m=1
M9 VDD N_7 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_7 Y VDD mp15  l=0.13u w=0.69u m=1
.ends dl02d2
* SPICE INPUT		Tue Jul 31 19:24:48 2018	dmnrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dmnrq0
.subckt dmnrq0 GND Q VDD CK D1 S0 D0
M1 GND S0 N_4 GND mn15  l=0.13u w=0.18u m=1
M2 N_18 D0 GND GND mn15  l=0.13u w=0.18u m=1
M3 N_18 N_4 N_6 GND mn15  l=0.13u w=0.18u m=1
M4 N_19 S0 N_6 GND mn15  l=0.13u w=0.18u m=1
M5 N_19 D1 GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.17u m=1
M7 N_20 N_12 N_9 GND mn15  l=0.13u w=0.17u m=1
M8 N_20 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M9 GND N_9 N_7 GND mn15  l=0.13u w=0.18u m=1
M10 N_6 N_2 N_9 GND mn15  l=0.13u w=0.28u m=1
M11 GND N_2 N_12 GND mn15  l=0.13u w=0.17u m=1
M12 N_22 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M13 N_22 N_12 N_14 GND mn15  l=0.13u w=0.17u m=1
M14 N_14 N_2 N_21 GND mn15  l=0.13u w=0.17u m=1
M15 N_21 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M16 Q N_14 GND GND mn15  l=0.13u w=0.26u m=1
M17 N_17 N_14 GND GND mn15  l=0.13u w=0.18u m=1
M18 N_4 S0 VDD VDD mp15  l=0.13u w=0.26u m=1
M19 N_39 D0 VDD VDD mp15  l=0.13u w=0.28u m=1
M20 N_39 S0 N_6 VDD mp15  l=0.13u w=0.28u m=1
M21 N_40 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M22 N_40 D1 VDD VDD mp15  l=0.13u w=0.28u m=1
M23 N_2 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M24 N_6 N_12 N_9 VDD mp15  l=0.13u w=0.42u m=1
M25 N_41 N_7 VDD VDD mp15  l=0.13u w=0.17u m=1
M26 VDD N_9 N_7 VDD mp15  l=0.13u w=0.26u m=1
M27 N_41 N_2 N_9 VDD mp15  l=0.13u w=0.17u m=1
M28 N_12 N_2 VDD VDD mp15  l=0.13u w=0.42u m=1
M29 N_43 N_7 VDD VDD mp15  l=0.13u w=0.27u m=1
M30 N_14 N_12 N_42 VDD mp15  l=0.13u w=0.17u m=1
M31 N_14 N_2 N_43 VDD mp15  l=0.13u w=0.27u m=1
M32 N_42 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M33 VDD N_14 Q VDD mp15  l=0.13u w=0.4u m=1
M34 N_17 N_14 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends dmnrq0
* SPICE INPUT		Tue Jul 31 19:25:01 2018	dmnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dmnrq1
.subckt dmnrq1 GND Q VDD CK D1 S0 D0
M1 N_5 N_6 N_18 GND mn15  l=0.13u w=0.17u m=1
M2 N_19 N_3 N_5 GND mn15  l=0.13u w=0.36u m=1
M3 GND N_6 N_3 GND mn15  l=0.13u w=0.2u m=1
M4 N_18 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_19 N_15 GND GND mn15  l=0.13u w=0.36u m=1
M6 GND S0 N_8 GND mn15  l=0.13u w=0.17u m=1
M7 N_20 D0 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_20 N_8 N_10 GND mn15  l=0.13u w=0.28u m=1
M9 N_21 S0 N_10 GND mn15  l=0.13u w=0.28u m=1
M10 N_21 D1 GND GND mn15  l=0.13u w=0.28u m=1
M11 GND CK N_6 GND mn15  l=0.13u w=0.2u m=1
M12 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_13 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M14 N_10 N_6 N_16 GND mn15  l=0.13u w=0.28u m=1
M15 N_15 N_16 GND GND mn15  l=0.13u w=0.28u m=1
M16 N_22 N_3 N_16 GND mn15  l=0.13u w=0.17u m=1
M17 N_22 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M18 VDD S0 N_8 VDD mp15  l=0.13u w=0.24u m=1
M19 N_39 D0 VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_10 S0 N_39 VDD mp15  l=0.13u w=0.42u m=1
M21 N_40 N_8 N_10 VDD mp15  l=0.13u w=0.42u m=1
M22 N_40 D1 VDD VDD mp15  l=0.13u w=0.42u m=1
M23 N_6 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M24 N_41 N_6 N_16 VDD mp15  l=0.13u w=0.17u m=1
M25 VDD N_16 N_15 VDD mp15  l=0.13u w=0.42u m=1
M26 N_10 N_3 N_16 VDD mp15  l=0.13u w=0.42u m=1
M27 N_41 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 N_43 N_6 N_5 VDD mp15  l=0.13u w=0.52u m=1
M29 N_5 N_3 N_42 VDD mp15  l=0.13u w=0.17u m=1
M30 N_3 N_6 VDD VDD mp15  l=0.13u w=0.51u m=1
M31 N_42 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_43 N_15 VDD VDD mp15  l=0.13u w=0.52u m=1
M33 VDD N_5 Q VDD mp15  l=0.13u w=0.69u m=1
M34 N_13 N_5 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends dmnrq1
* SPICE INPUT		Tue Jul 31 19:25:14 2018	dmnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=dmnrq2
.subckt dmnrq2 GND Q VDD CK D1 S0 D0
M1 GND S0 N_4 GND mn15  l=0.13u w=0.24u m=1
M2 N_19 D0 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_6 N_4 N_19 GND mn15  l=0.13u w=0.28u m=1
M4 N_20 S0 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_20 D1 GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 CK GND GND mn15  l=0.13u w=0.28u m=1
M7 N_21 N_18 GND GND mn15  l=0.13u w=0.41u m=1
M8 N_21 N_13 N_10 GND mn15  l=0.13u w=0.41u m=1
M9 N_22 N_3 N_10 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_8 N_22 GND mn15  l=0.13u w=0.17u m=1
M11 Q N_10 GND GND mn15  l=0.13u w=0.46u m=1
M12 Q N_10 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_8 N_10 GND GND mn15  l=0.13u w=0.37u m=1
M14 N_23 N_13 N_16 GND mn15  l=0.13u w=0.17u m=1
M15 N_16 N_3 N_6 GND mn15  l=0.13u w=0.41u m=1
M16 GND N_18 N_23 GND mn15  l=0.13u w=0.17u m=1
M17 N_18 N_16 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_18 N_16 GND GND mn15  l=0.13u w=0.15u m=1
M19 GND N_3 N_13 GND mn15  l=0.13u w=0.23u m=1
M20 VDD S0 N_4 VDD mp15  l=0.13u w=0.37u m=1
M21 N_41 D0 VDD VDD mp15  l=0.13u w=0.42u m=1
M22 N_6 S0 N_41 VDD mp15  l=0.13u w=0.42u m=1
M23 N_42 N_4 N_6 VDD mp15  l=0.13u w=0.42u m=1
M24 N_42 D1 VDD VDD mp15  l=0.13u w=0.42u m=1
M25 N_3 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M26 N_16 N_13 N_6 VDD mp15  l=0.13u w=0.63u m=1
M27 N_43 N_3 N_16 VDD mp15  l=0.13u w=0.17u m=1
M28 N_43 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 VDD N_16 N_18 VDD mp15  l=0.13u w=0.63u m=1
M30 VDD N_3 N_13 VDD mp15  l=0.13u w=0.57u m=1
M31 N_44 N_18 VDD VDD mp15  l=0.13u w=0.62u m=1
M32 N_44 N_3 N_10 VDD mp15  l=0.13u w=0.62u m=1
M33 N_45 N_13 N_10 VDD mp15  l=0.13u w=0.17u m=1
M34 VDD N_8 N_45 VDD mp15  l=0.13u w=0.17u m=1
M35 N_8 N_10 VDD VDD mp15  l=0.13u w=0.55u m=1
M36 Q N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M37 Q N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends dmnrq2
* SPICE INPUT		Tue Jul 31 19:26:49 2018	fillercap16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap16
.subckt fillercap16 GND VDD
M1 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M2 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M3 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M4 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
.ends fillercap16
* SPICE INPUT		Tue Jul 31 19:27:11 2018	fillercap3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap3
.subckt fillercap3 VDD GND
M1 VDD GND VDD VDD mp15  l=0.33u w=0.69u m=1
.ends fillercap3
* SPICE INPUT		Tue Jul 31 19:27:24 2018	fillercap32
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap32
.subckt fillercap32 GND VDD
M1 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M2 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M3 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M4 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M5 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M6 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M7 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M8 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M9 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M10 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
.ends fillercap32
* SPICE INPUT		Tue Jul 31 19:27:37 2018	fillercap4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap4
.subckt fillercap4 VDD GND
M1 VDD GND VDD VDD mp15  l=0.67u w=0.69u m=1
.ends fillercap4
* SPICE INPUT		Tue Jul 31 19:27:50 2018	fillercap6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap6
.subckt fillercap6 VDD GND
M1 VDD GND VDD VDD mp15  l=0.33u w=1.22u m=1
.ends fillercap6
* SPICE INPUT		Tue Jul 31 19:28:03 2018	fillercap64
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap64
.subckt fillercap64 GND VDD
M1 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M2 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M3 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M4 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M5 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M6 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M7 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M8 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M9 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M10 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M11 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M12 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M13 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M14 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M15 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M16 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M17 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M18 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M19 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M20 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M21 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
M22 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
.ends fillercap64
* SPICE INPUT		Tue Jul 31 19:28:16 2018	fillercap8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=fillercap8
.subckt fillercap8 VDD GND
M1 VDD GND VDD VDD mp15  l=0.67u w=1.22u m=1
.ends fillercap8
* SPICE INPUT		Tue Jul 31 19:28:38 2018	inv0d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d0
.subckt inv0d0 GND VDD Y A
M1 Y A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends inv0d0
* SPICE INPUT		Tue Jul 31 19:28:51 2018	inv0d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d1
.subckt inv0d1 GND VDD Y A
M1 Y A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d1
* SPICE INPUT		Tue Jul 31 19:29:04 2018	inv0d12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d12
.subckt inv0d12 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A Y GND mn15  l=0.13u w=0.46u m=1
M8 Y A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND A Y GND mn15  l=0.13u w=0.46u m=1
M10 Y A GND GND mn15  l=0.13u w=0.46u m=1
M11 GND A Y GND mn15  l=0.13u w=0.46u m=1
M12 Y A GND GND mn15  l=0.13u w=0.46u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d12
* SPICE INPUT		Tue Jul 31 19:29:17 2018	inv0d16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d16
.subckt inv0d16 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A Y GND mn15  l=0.13u w=0.46u m=1
M8 Y A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND A Y GND mn15  l=0.13u w=0.46u m=1
M10 Y A GND GND mn15  l=0.13u w=0.46u m=1
M11 GND A Y GND mn15  l=0.13u w=0.46u m=1
M12 Y A GND GND mn15  l=0.13u w=0.46u m=1
M13 GND A Y GND mn15  l=0.13u w=0.46u m=1
M14 Y A GND GND mn15  l=0.13u w=0.46u m=1
M15 GND A Y GND mn15  l=0.13u w=0.46u m=1
M16 Y A GND GND mn15  l=0.13u w=0.46u m=1
M17 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M31 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d16
* SPICE INPUT		Tue Jul 31 19:29:30 2018	inv0d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d2
.subckt inv0d2 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M4 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d2
* SPICE INPUT		Tue Jul 31 19:29:42 2018	inv0d20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d20
.subckt inv0d20 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A Y GND mn15  l=0.13u w=0.46u m=1
M8 Y A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND A Y GND mn15  l=0.13u w=0.46u m=1
M10 Y A GND GND mn15  l=0.13u w=0.46u m=1
M11 GND A Y GND mn15  l=0.13u w=0.46u m=1
M12 Y A GND GND mn15  l=0.13u w=0.46u m=1
M13 GND A Y GND mn15  l=0.13u w=0.46u m=1
M14 Y A GND GND mn15  l=0.13u w=0.46u m=1
M15 GND A Y GND mn15  l=0.13u w=0.46u m=1
M16 Y A GND GND mn15  l=0.13u w=0.46u m=1
M17 GND A Y GND mn15  l=0.13u w=0.46u m=1
M18 Y A GND GND mn15  l=0.13u w=0.46u m=1
M19 GND A Y GND mn15  l=0.13u w=0.46u m=1
M20 Y A GND GND mn15  l=0.13u w=0.46u m=1
M21 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M31 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M33 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M34 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M35 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M36 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M37 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M38 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M39 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M40 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d20
* SPICE INPUT		Tue Jul 31 19:29:55 2018	inv0d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d3
.subckt inv0d3 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y A GND GND mn15  l=0.13u w=0.46u m=1
M4 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M5 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d3
* SPICE INPUT		Tue Jul 31 19:30:08 2018	inv0d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d4
.subckt inv0d4 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M6 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d4
* SPICE INPUT		Tue Jul 31 19:30:21 2018	inv0d5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d5
.subckt inv0d5 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A Y GND mn15  l=0.13u w=0.46u m=1
M5 Y A GND GND mn15  l=0.13u w=0.46u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d5
* SPICE INPUT		Tue Jul 31 19:30:34 2018	inv0d6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d6
.subckt inv0d6 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d6
* SPICE INPUT		Tue Jul 31 19:30:47 2018	inv0d7
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d7
.subckt inv0d7 GND Y VDD A
M1 Y A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A Y GND mn15  l=0.13u w=0.46u m=1
M5 Y A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A Y GND mn15  l=0.13u w=0.46u m=1
M7 Y A GND GND mn15  l=0.13u w=0.46u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d7
* SPICE INPUT		Tue Jul 31 19:31:00 2018	inv0d8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0d8
.subckt inv0d8 Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.46u m=1
M2 GND A Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A Y GND mn15  l=0.13u w=0.46u m=1
M4 Y A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A Y GND mn15  l=0.13u w=0.46u m=1
M6 Y A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND A Y GND mn15  l=0.13u w=0.46u m=1
M8 Y A GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends inv0d8
* SPICE INPUT		Tue Jul 31 19:31:13 2018	inv0dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0dm
.subckt inv0dm GND VDD Y A
M1 Y A GND GND mn15  l=0.13u w=0.36u m=1
M2 Y A VDD VDD mp15  l=0.13u w=0.55u m=1
.ends inv0dm
* SPICE INPUT		Tue Jul 31 19:31:26 2018	inv0dp
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=inv0dp
.subckt inv0dp Y GND VDD A
M1 GND A Y GND mn15  l=0.13u w=0.355u m=1
M2 GND A Y GND mn15  l=0.13u w=0.355u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
M4 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
.ends inv0dp
* SPICE INPUT		Tue Jul 31 19:31:40 2018	invod8d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invod8d1
.subckt invod8d1 GND Y0 Y6 Y5 Y2 Y1 Y7 Y4 Y3 VDD A
M1 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y0 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y6 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 Y5 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 Y1 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y2 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y7 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M8 Y4 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y3 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M10 VDD A N_4 VDD mp15  l=0.13u w=0.69u m=1
.ends invod8d1
* SPICE INPUT		Tue Jul 31 19:31:52 2018	invtld0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld0
.subckt invtld0 GND Y VDD A E
M1 GND E N_3 GND mn15  l=0.13u w=0.26u m=1
M2 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y E N_6 GND mn15  l=0.13u w=0.26u m=1
M4 Y E N_7 GND mn15  l=0.13u w=0.26u m=1
M5 GND A N_6 GND mn15  l=0.13u w=0.26u m=1
M6 VDD E N_3 VDD mp15  l=0.13u w=0.4u m=1
M7 N_14 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 Y N_3 N_13 VDD mp15  l=0.13u w=0.4u m=1
M9 Y N_3 N_14 VDD mp15  l=0.13u w=0.4u m=1
M10 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends invtld0
* SPICE INPUT		Tue Jul 31 19:32:06 2018	invtld1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld1
.subckt invtld1 Y VDD GND A E
M1 GND E N_3 GND mn15  l=0.13u w=0.31u m=1
M2 GND A N_13 GND mn15  l=0.13u w=0.46u m=1
M3 Y E N_15 GND mn15  l=0.13u w=0.46u m=1
M4 Y E N_13 GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_15 GND mn15  l=0.13u w=0.46u m=1
M6 VDD E N_3 VDD mp15  l=0.13u w=0.46u m=1
M7 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_7 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M9 Y N_3 N_8 VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends invtld1
* SPICE INPUT		Tue Jul 31 19:32:19 2018	invtld12
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld12
.subckt invtld12 GND Y VDD E A
M1 GND E N_2 GND mn15  l=0.13u w=0.42u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.31u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.31u m=1
M4 N_7 N_5 GND GND mn15  l=0.13u w=0.455u m=1
M5 N_7 N_5 GND GND mn15  l=0.13u w=0.45u m=1
M6 N_7 N_5 GND GND mn15  l=0.13u w=0.45u m=1
M7 N_7 N_5 GND GND mn15  l=0.13u w=0.45u m=1
M8 N_7 N_5 GND GND mn15  l=0.13u w=0.415u m=1
M9 N_6 E N_7 GND mn15  l=0.13u w=0.4u m=1
M10 N_6 E N_7 GND mn15  l=0.13u w=0.405u m=1
M11 N_7 E N_6 GND mn15  l=0.13u w=0.395u m=1
M12 GND N_2 N_7 GND mn15  l=0.13u w=0.37u m=1
M13 N_7 N_2 GND GND mn15  l=0.13u w=0.37u m=1
M14 N_7 N_2 GND GND mn15  l=0.13u w=0.37u m=1
M15 Y N_7 GND GND mn15  l=0.13u w=0.43u m=1
M16 GND N_7 Y GND mn15  l=0.13u w=0.4u m=1
M17 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M18 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M19 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M20 GND N_7 Y GND mn15  l=0.13u w=0.42u m=1
M21 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M22 GND N_7 Y GND mn15  l=0.13u w=0.42u m=1
M23 Y N_7 GND GND mn15  l=0.13u w=0.4u m=1
M24 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M25 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M26 Y N_7 GND GND mn15  l=0.13u w=0.42u m=1
M27 Y N_7 GND GND mn15  l=0.13u w=0.37u m=1
M28 N_2 E VDD VDD mp15  l=0.13u w=0.63u m=1
M29 N_5 A VDD VDD mp15  l=0.13u w=0.47u m=1
M30 N_5 A VDD VDD mp15  l=0.13u w=0.47u m=1
M31 VDD N_6 Y VDD mp15  l=0.13u w=0.72u m=1
M32 VDD N_6 Y VDD mp15  l=0.13u w=0.72u m=1
M33 Y N_6 VDD VDD mp15  l=0.13u w=0.72u m=1
M34 VDD N_6 Y VDD mp15  l=0.13u w=0.72u m=1
M35 Y N_6 VDD VDD mp15  l=0.13u w=0.72u m=1
M36 VDD N_6 Y VDD mp15  l=0.13u w=0.71u m=1
M37 VDD N_6 Y VDD mp15  l=0.13u w=0.71u m=1
M38 Y N_6 VDD VDD mp15  l=0.13u w=0.71u m=1
M39 VDD N_6 Y VDD mp15  l=0.13u w=0.68u m=1
M40 VDD N_6 Y VDD mp15  l=0.13u w=0.64u m=1
M41 VDD N_6 Y VDD mp15  l=0.13u w=0.64u m=1
M42 VDD N_6 Y VDD mp15  l=0.13u w=0.59u m=1
M43 N_6 N_5 VDD VDD mp15  l=0.13u w=0.54u m=1
M44 N_6 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M45 N_6 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M46 N_6 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M47 N_6 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M48 N_6 E VDD VDD mp15  l=0.13u w=0.57u m=1
M49 N_6 E VDD VDD mp15  l=0.13u w=0.57u m=1
M50 VDD E N_6 VDD mp15  l=0.13u w=0.48u m=1
M51 N_7 N_2 N_6 VDD mp15  l=0.13u w=0.76u m=1
M52 N_6 N_2 N_7 VDD mp15  l=0.13u w=0.78u m=1
M53 N_7 N_2 N_6 VDD mp15  l=0.13u w=0.78u m=1
.ends invtld12
* SPICE INPUT		Tue Jul 31 19:32:33 2018	invtld16
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld16
.subckt invtld16 GND Y A VDD E
M1 N_3 N_16 GND GND mn15  l=0.13u w=0.37u m=1
M2 N_3 N_16 GND GND mn15  l=0.13u w=0.37u m=1
M3 GND N_16 N_3 GND mn15  l=0.13u w=0.37u m=1
M4 N_3 N_16 GND GND mn15  l=0.13u w=0.35u m=1
M5 GND N_5 N_3 GND mn15  l=0.13u w=0.41u m=1
M6 GND N_5 N_3 GND mn15  l=0.13u w=0.44u m=1
M7 GND N_5 N_3 GND mn15  l=0.13u w=0.44u m=1
M8 N_3 N_5 GND GND mn15  l=0.13u w=0.44u m=1
M9 GND N_5 N_3 GND mn15  l=0.13u w=0.44u m=1
M10 N_3 N_5 GND GND mn15  l=0.13u w=0.39u m=1
M11 N_3 N_5 GND GND mn15  l=0.13u w=0.37u m=1
M12 GND A N_5 GND mn15  l=0.13u w=0.39u m=1
M13 N_5 A GND GND mn15  l=0.13u w=0.39u m=1
M14 GND E N_16 GND mn15  l=0.13u w=0.44u m=1
M15 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M16 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M17 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M18 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M19 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M20 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M21 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M22 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M23 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M24 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M25 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M26 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M27 Y N_3 GND GND mn15  l=0.13u w=0.39u m=1
M28 GND N_3 Y GND mn15  l=0.13u w=0.39u m=1
M29 Y N_3 GND GND mn15  l=0.13u w=0.39u m=1
M30 Y N_3 GND GND mn15  l=0.13u w=0.39u m=1
M31 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M32 N_37 E N_3 GND mn15  l=0.13u w=0.55u m=1
M33 N_3 E N_37 GND mn15  l=0.13u w=0.55u m=1
M34 N_3 E N_37 GND mn15  l=0.13u w=0.46u m=1
M35 N_37 E VDD VDD mp15  l=0.13u w=0.76u m=1
M36 N_37 E VDD VDD mp15  l=0.13u w=0.76u m=1
M37 VDD E N_37 VDD mp15  l=0.13u w=0.67u m=1
M38 N_16 E VDD VDD mp15  l=0.13u w=0.67u m=1
M39 N_37 N_5 VDD VDD mp15  l=0.13u w=0.63u m=1
M40 VDD N_5 N_37 VDD mp15  l=0.13u w=0.63u m=1
M41 N_37 N_5 VDD VDD mp15  l=0.13u w=0.63u m=1
M42 VDD N_5 N_37 VDD mp15  l=0.13u w=0.63u m=1
M43 N_37 N_5 VDD VDD mp15  l=0.13u w=0.63u m=1
M44 VDD N_5 N_37 VDD mp15  l=0.13u w=0.63u m=1
M45 N_37 N_5 VDD VDD mp15  l=0.13u w=0.62u m=1
M46 VDD A N_5 VDD mp15  l=0.13u w=0.59u m=1
M47 N_5 A VDD VDD mp15  l=0.13u w=0.59u m=1
M48 N_3 N_16 N_37 VDD mp15  l=0.13u w=0.54u m=1
M49 N_37 N_16 N_3 VDD mp15  l=0.13u w=0.54u m=1
M50 N_37 N_16 N_3 VDD mp15  l=0.13u w=0.54u m=1
M51 N_3 N_16 N_37 VDD mp15  l=0.13u w=0.54u m=1
M52 N_37 N_16 N_3 VDD mp15  l=0.13u w=0.54u m=1
M53 N_37 N_16 N_3 VDD mp15  l=0.13u w=0.4u m=1
M54 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M55 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M56 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M57 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M58 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M59 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M60 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M61 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M62 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M63 Y N_37 VDD VDD mp15  l=0.13u w=0.69u m=1
M64 VDD N_37 Y VDD mp15  l=0.13u w=0.69u m=1
M65 Y N_37 VDD VDD mp15  l=0.13u w=0.64u m=1
M66 Y N_37 VDD VDD mp15  l=0.13u w=0.61u m=1
M67 VDD N_37 Y VDD mp15  l=0.13u w=0.55u m=1
M68 Y N_37 VDD VDD mp15  l=0.13u w=0.55u m=1
M69 VDD N_37 Y VDD mp15  l=0.13u w=0.55u m=1
M70 Y N_37 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends invtld16
* SPICE INPUT		Tue Jul 31 19:32:46 2018	invtld2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld2
.subckt invtld2 GND Y VDD E A
M1 N_3 E GND GND mn15  l=0.13u w=0.46u m=1
M2 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_5 E Y GND mn15  l=0.13u w=0.42u m=1
M7 N_5 E Y GND mn15  l=0.13u w=0.57u m=1
M8 N_5 E Y GND mn15  l=0.13u w=0.57u m=1
M9 Y E N_5 GND mn15  l=0.13u w=0.29u m=1
M10 VDD E N_3 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD A N_14 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_14 VDD mp15  l=0.13u w=0.69u m=1
M13 N_14 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_14 VDD mp15  l=0.13u w=0.69u m=1
M15 Y N_3 N_14 VDD mp15  l=0.13u w=0.57u m=1
M16 Y N_3 N_14 VDD mp15  l=0.13u w=0.57u m=1
M17 Y N_3 N_14 VDD mp15  l=0.13u w=0.57u m=1
M18 N_14 N_3 Y VDD mp15  l=0.13u w=0.57u m=1
M19 Y N_3 N_14 VDD mp15  l=0.13u w=0.46u m=1
.ends invtld2
* SPICE INPUT		Tue Jul 31 19:33:00 2018	invtld20
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld20
.subckt invtld20 GND Y VDD E A
M1 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M2 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_25 GND GND mn15  l=0.13u w=0.4u m=1
M4 Y N_25 GND GND mn15  l=0.13u w=0.4u m=1
M5 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M8 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_25 GND GND mn15  l=0.13u w=0.385u m=1
M10 Y N_25 GND GND mn15  l=0.13u w=0.315u m=1
M11 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M12 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M13 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M14 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M15 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M16 Y N_25 GND GND mn15  l=0.13u w=0.4u m=1
M17 Y N_25 GND GND mn15  l=0.13u w=0.4u m=1
M18 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M19 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M20 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M21 Y N_25 GND GND mn15  l=0.13u w=0.46u m=1
M22 N_25 E N_24 GND mn15  l=0.13u w=0.56u m=1
M23 N_25 E N_24 GND mn15  l=0.13u w=0.56u m=1
M24 N_25 E N_24 GND mn15  l=0.13u w=0.56u m=1
M25 N_24 E N_25 GND mn15  l=0.13u w=0.27u m=1
M26 GND A N_32 GND mn15  l=0.13u w=0.46u m=1
M27 N_32 A GND GND mn15  l=0.13u w=0.46u m=1
M28 GND N_32 N_25 GND mn15  l=0.13u w=0.46u m=1
M29 N_25 N_32 GND GND mn15  l=0.13u w=0.46u m=1
M30 GND N_32 N_25 GND mn15  l=0.13u w=0.46u m=1
M31 N_25 N_32 GND GND mn15  l=0.13u w=0.46u m=1
M32 GND N_32 N_25 GND mn15  l=0.13u w=0.46u m=1
M33 N_25 N_32 GND GND mn15  l=0.13u w=0.46u m=1
M34 GND N_32 N_25 GND mn15  l=0.13u w=0.46u m=1
M35 N_25 N_32 GND GND mn15  l=0.13u w=0.46u m=1
M36 GND E N_29 GND mn15  l=0.13u w=0.46u m=1
M37 N_25 N_29 GND GND mn15  l=0.13u w=0.46u m=1
M38 N_25 N_29 GND GND mn15  l=0.13u w=0.46u m=1
M39 GND N_29 N_25 GND mn15  l=0.13u w=0.46u m=1
M40 N_25 N_29 GND GND mn15  l=0.13u w=0.46u m=1
M41 VDD A N_32 VDD mp15  l=0.13u w=0.69u m=1
M42 N_32 A VDD VDD mp15  l=0.13u w=0.69u m=1
M43 VDD N_32 N_24 VDD mp15  l=0.13u w=0.69u m=1
M44 N_24 N_32 VDD VDD mp15  l=0.13u w=0.69u m=1
M45 VDD N_32 N_24 VDD mp15  l=0.13u w=0.69u m=1
M46 N_24 N_32 VDD VDD mp15  l=0.13u w=0.69u m=1
M47 VDD N_32 N_24 VDD mp15  l=0.13u w=0.69u m=1
M48 N_24 N_32 VDD VDD mp15  l=0.13u w=0.69u m=1
M49 VDD N_32 N_24 VDD mp15  l=0.13u w=0.69u m=1
M50 N_24 N_32 VDD VDD mp15  l=0.13u w=0.69u m=1
M51 N_29 E VDD VDD mp15  l=0.13u w=0.69u m=1
M52 N_24 E VDD VDD mp15  l=0.13u w=0.69u m=1
M53 N_24 E VDD VDD mp15  l=0.13u w=0.69u m=1
M54 VDD E N_24 VDD mp15  l=0.13u w=0.69u m=1
M55 N_24 E VDD VDD mp15  l=0.13u w=0.69u m=1
M56 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.58u m=1
M57 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.58u m=1
M58 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.58u m=1
M59 N_24 N_29 N_25 VDD mp15  l=0.13u w=0.58u m=1
M60 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.58u m=1
M61 N_24 N_29 N_25 VDD mp15  l=0.13u w=0.58u m=1
M62 N_25 N_29 N_24 VDD mp15  l=0.13u w=0.4u m=1
M63 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M64 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M65 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M66 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M67 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M68 Y N_24 VDD VDD mp15  l=0.13u w=0.665u m=1
M69 Y N_24 VDD VDD mp15  l=0.13u w=0.665u m=1
M70 VDD N_24 Y VDD mp15  l=0.13u w=0.665u m=1
M71 Y N_24 VDD VDD mp15  l=0.13u w=0.665u m=1
M72 VDD N_24 Y VDD mp15  l=0.13u w=0.65u m=1
M73 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M74 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M75 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M76 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M77 Y N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M78 VDD N_24 Y VDD mp15  l=0.13u w=0.69u m=1
M79 Y N_24 VDD VDD mp15  l=0.13u w=0.61u m=1
M80 VDD N_24 Y VDD mp15  l=0.13u w=0.57u m=1
M81 Y N_24 VDD VDD mp15  l=0.13u w=0.57u m=1
M82 VDD N_24 Y VDD mp15  l=0.13u w=0.57u m=1
M83 Y N_24 VDD VDD mp15  l=0.13u w=0.57u m=1
.ends invtld20
* SPICE INPUT		Tue Jul 31 19:33:13 2018	invtld3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld3
.subckt invtld3 GND Y VDD E A
M1 N_4 A GND GND mn15  l=0.13u w=0.3u m=1
M2 N_3 N_4 GND GND mn15  l=0.13u w=0.56u m=1
M3 GND N_5 N_3 GND mn15  l=0.13u w=0.28u m=1
M4 GND E N_5 GND mn15  l=0.13u w=0.3u m=1
M5 N_7 E N_3 GND mn15  l=0.13u w=0.3u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M8 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M9 VDD A N_4 VDD mp15  l=0.13u w=0.42u m=1
M10 VDD N_4 N_7 VDD mp15  l=0.13u w=0.42u m=1
M11 VDD N_4 N_7 VDD mp15  l=0.13u w=0.41u m=1
M12 N_3 N_5 N_7 VDD mp15  l=0.13u w=0.58u m=1
M13 VDD E N_7 VDD mp15  l=0.13u w=0.41u m=1
M14 VDD E N_5 VDD mp15  l=0.13u w=0.42u m=1
M15 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 Y N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends invtld3
* SPICE INPUT		Tue Jul 31 19:33:26 2018	invtld4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld4
.subckt invtld4 Y GND E A VDD
M1 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_8 E GND GND mn15  l=0.13u w=0.3u m=1
M6 N_9 A GND GND mn15  l=0.13u w=0.34u m=1
M7 N_13 N_9 GND GND mn15  l=0.13u w=0.37u m=1
M8 N_13 N_9 GND GND mn15  l=0.13u w=0.37u m=1
M9 N_13 N_8 GND GND mn15  l=0.13u w=0.37u m=1
M10 N_13 E N_10 GND mn15  l=0.13u w=0.39u m=1
M11 N_8 E VDD VDD mp15  l=0.13u w=0.4u m=1
M12 N_9 A VDD VDD mp15  l=0.13u w=0.48u m=1
M13 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_9 N_10 VDD mp15  l=0.13u w=0.55u m=1
M18 N_10 N_9 VDD VDD mp15  l=0.13u w=0.55u m=1
M19 VDD E N_10 VDD mp15  l=0.13u w=0.55u m=1
M20 N_13 N_8 N_10 VDD mp15  l=0.13u w=0.64u m=1
.ends invtld4
* SPICE INPUT		Tue Jul 31 19:33:40 2018	invtld6
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld6
.subckt invtld6 GND Y VDD E A
M1 N_4 A GND GND mn15  l=0.13u w=0.39u m=1
M2 N_3 E GND GND mn15  l=0.13u w=0.3u m=1
M3 GND N_4 N_5 GND mn15  l=0.13u w=0.37u m=1
M4 N_5 N_4 GND GND mn15  l=0.13u w=0.37u m=1
M5 N_5 N_4 GND GND mn15  l=0.13u w=0.37u m=1
M6 N_6 E N_5 GND mn15  l=0.13u w=0.59u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_5 N_3 GND GND mn15  l=0.13u w=0.55u m=1
M14 N_4 A VDD VDD mp15  l=0.13u w=0.58u m=1
M15 N_3 E VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_6 N_4 VDD VDD mp15  l=0.13u w=0.57u m=1
M17 N_6 N_4 VDD VDD mp15  l=0.13u w=0.64u m=1
M18 N_6 N_4 VDD VDD mp15  l=0.13u w=0.45u m=1
M19 N_6 E VDD VDD mp15  l=0.13u w=0.41u m=1
M20 VDD E N_6 VDD mp15  l=0.13u w=0.41u m=1
M21 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.595u m=1
M22 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.565u m=1
M23 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M28 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends invtld6
* SPICE INPUT		Tue Jul 31 19:33:52 2018	invtld8
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtld8
.subckt invtld8 GND Y VDD E A
M1 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 E GND GND mn15  l=0.13u w=0.39u m=1
M3 N_5 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_5 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_10 E N_5 GND mn15  l=0.13u w=0.41u m=1
M7 N_5 E N_10 GND mn15  l=0.13u w=0.38u m=1
M8 GND N_3 N_5 GND mn15  l=0.13u w=0.345u m=1
M9 GND N_3 N_5 GND mn15  l=0.13u w=0.345u m=1
M10 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M13 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M14 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M15 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M16 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M17 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M18 N_4 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 VDD E N_3 VDD mp15  l=0.13u w=0.58u m=1
M20 N_10 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_10 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_10 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_10 E VDD VDD mp15  l=0.13u w=0.605u m=1
M24 VDD E N_10 VDD mp15  l=0.13u w=0.415u m=1
M25 N_5 N_3 N_10 VDD mp15  l=0.13u w=0.77u m=1
M26 N_5 N_3 N_10 VDD mp15  l=0.13u w=0.77u m=1
M27 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M33 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M34 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends invtld8
* SPICE INPUT		Tue Jul 31 19:34:05 2018	invtldm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=invtldm
.subckt invtldm VDD Y A E GND
M1 Y E N_13 GND mn15  l=0.13u w=0.47u m=1
M2 N_14 E Y GND mn15  l=0.13u w=0.24u m=1
M3 N_3 E GND GND mn15  l=0.13u w=0.26u m=1
M4 N_14 A GND GND mn15  l=0.13u w=0.24u m=1
M5 GND A N_13 GND mn15  l=0.13u w=0.47u m=1
M6 N_3 E VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_7 A VDD VDD mp15  l=0.13u w=0.55u m=1
M8 N_7 N_3 Y VDD mp15  l=0.13u w=0.55u m=1
M9 Y N_3 N_6 VDD mp15  l=0.13u w=0.55u m=1
M10 N_6 A VDD VDD mp15  l=0.13u w=0.55u m=1
.ends invtldm
* SPICE INPUT		Tue Jul 31 19:34:18 2018	labhb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=labhb0
.subckt labhb0 GND QN Q D SN RN VDD G
M1 N_4 G GND GND mn15  l=0.13u w=0.17u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_7 N_2 N_6 GND mn15  l=0.13u w=0.17u m=1
M4 N_6 D N_5 GND mn15  l=0.13u w=0.18u m=1
M5 N_5 RN GND GND mn15  l=0.13u w=0.34u m=1
M6 N_18 N_4 N_7 GND mn15  l=0.13u w=0.17u m=1
M7 N_7 N_8 GND GND mn15  l=0.13u w=0.18u m=1
M8 GND SN N_8 GND mn15  l=0.13u w=0.18u m=1
M9 N_18 N_17 N_5 GND mn15  l=0.13u w=0.17u m=1
M10 QN N_17 GND GND mn15  l=0.13u w=0.26u m=1
M11 Q N_7 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_17 N_7 GND GND mn15  l=0.13u w=0.18u m=1
M13 N_4 G VDD VDD mp15  l=0.13u w=0.42u m=1
M14 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M15 N_22 D N_6 VDD mp15  l=0.13u w=0.33u m=1
M16 N_7 RN N_22 VDD mp15  l=0.13u w=0.3u m=1
M17 N_7 N_2 N_67 VDD mp15  l=0.13u w=0.17u m=1
M18 N_7 N_4 N_6 VDD mp15  l=0.13u w=0.42u m=1
M19 N_67 N_17 N_22 VDD mp15  l=0.13u w=0.17u m=1
M20 N_22 N_8 VDD VDD mp15  l=0.13u w=0.54u m=1
M21 N_8 SN VDD VDD mp15  l=0.13u w=0.26u m=1
M22 Q N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M23 N_17 N_7 VDD VDD mp15  l=0.13u w=0.26u m=1
M24 QN N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends labhb0
* SPICE INPUT		Tue Jul 31 19:34:32 2018	labhb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=labhb1
.subckt labhb1 GND QN Q VDD SN RN D G
M1 N_4 G GND GND mn15  l=0.13u w=0.2u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.2u m=1
M3 N_8 N_2 N_7 GND mn15  l=0.13u w=0.46u m=1
M4 N_10 D N_7 GND mn15  l=0.13u w=0.35u m=1
M5 N_10 RN GND GND mn15  l=0.13u w=0.35u m=1
M6 N_10 RN GND GND mn15  l=0.13u w=0.14u m=1
M7 N_8 N_4 N_18 GND mn15  l=0.13u w=0.17u m=1
M8 N_8 N_14 GND GND mn15  l=0.13u w=0.27u m=1
M9 N_14 SN GND GND mn15  l=0.13u w=0.14u m=1
M10 N_14 SN GND GND mn15  l=0.13u w=0.14u m=1
M11 QN N_17 GND GND mn15  l=0.13u w=0.43u m=1
M12 N_18 N_17 N_10 GND mn15  l=0.13u w=0.17u m=1
M13 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M14 N_17 N_8 GND GND mn15  l=0.13u w=0.28u m=1
M15 N_4 G VDD VDD mp15  l=0.13u w=0.51u m=1
M16 N_2 N_4 VDD VDD mp15  l=0.13u w=0.51u m=1
M17 N_22 D N_7 VDD mp15  l=0.13u w=0.52u m=1
M18 N_8 RN N_22 VDD mp15  l=0.13u w=0.39u m=1
M19 N_8 N_2 N_71 VDD mp15  l=0.13u w=0.17u m=1
M20 N_8 N_4 N_7 VDD mp15  l=0.13u w=0.65u m=1
M21 N_71 N_17 N_22 VDD mp15  l=0.13u w=0.17u m=1
M22 N_22 N_14 VDD VDD mp15  l=0.13u w=0.63u m=1
M23 N_14 SN VDD VDD mp15  l=0.13u w=0.195u m=1
M24 N_14 SN VDD VDD mp15  l=0.13u w=0.195u m=1
M25 QN N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_17 N_8 VDD VDD mp15  l=0.13u w=0.36u m=1
.ends labhb1
* SPICE INPUT		Tue Jul 31 19:34:45 2018	labhb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=labhb2
.subckt labhb2 GND QN Q VDD SN RN D G
M1 N_4 G GND GND mn15  l=0.13u w=0.27u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_6 D N_5 GND mn15  l=0.13u w=0.225u m=1
M4 N_5 D N_6 GND mn15  l=0.13u w=0.235u m=1
M5 N_5 N_2 N_8 GND mn15  l=0.13u w=0.24u m=1
M6 N_8 N_2 N_5 GND mn15  l=0.13u w=0.21u m=1
M7 N_25 N_4 N_8 GND mn15  l=0.13u w=0.17u m=1
M8 GND RN N_6 GND mn15  l=0.13u w=0.23u m=1
M9 N_6 RN GND GND mn15  l=0.13u w=0.23u m=1
M10 N_25 N_23 N_6 GND mn15  l=0.13u w=0.17u m=1
M11 GND N_19 N_8 GND mn15  l=0.13u w=0.185u m=1
M12 N_8 N_19 GND GND mn15  l=0.13u w=0.185u m=1
M13 GND SN N_19 GND mn15  l=0.13u w=0.14u m=1
M14 N_19 SN GND GND mn15  l=0.13u w=0.14u m=1
M15 GND N_23 QN GND mn15  l=0.13u w=0.46u m=1
M16 GND N_23 QN GND mn15  l=0.13u w=0.43u m=1
M17 GND N_8 Q GND mn15  l=0.13u w=0.46u m=1
M18 GND N_8 Q GND mn15  l=0.13u w=0.46u m=1
M19 GND N_8 N_23 GND mn15  l=0.13u w=0.37u m=1
M20 N_4 G VDD VDD mp15  l=0.13u w=0.67u m=1
M21 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M22 N_5 N_4 N_8 VDD mp15  l=0.13u w=0.56u m=1
M23 N_5 N_4 N_8 VDD mp15  l=0.13u w=0.56u m=1
M24 N_5 D N_29 VDD mp15  l=0.13u w=0.29u m=1
M25 N_5 D N_29 VDD mp15  l=0.13u w=0.29u m=1
M26 N_5 D N_29 VDD mp15  l=0.13u w=0.29u m=1
M27 N_5 D N_29 VDD mp15  l=0.13u w=0.29u m=1
M28 N_98 N_2 N_8 VDD mp15  l=0.13u w=0.17u m=1
M29 N_29 RN N_8 VDD mp15  l=0.13u w=0.54u m=1
M30 N_98 N_23 N_29 VDD mp15  l=0.13u w=0.17u m=1
M31 N_29 N_19 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 N_29 N_19 VDD VDD mp15  l=0.13u w=0.69u m=1
M33 N_19 SN VDD VDD mp15  l=0.13u w=0.21u m=1
M34 VDD SN N_19 VDD mp15  l=0.13u w=0.21u m=1
M35 QN N_23 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 VDD N_23 QN VDD mp15  l=0.13u w=0.69u m=1
M37 VDD N_8 Q VDD mp15  l=0.13u w=0.69u m=1
M38 VDD N_8 Q VDD mp15  l=0.13u w=0.69u m=1
M39 VDD N_8 N_23 VDD mp15  l=0.13u w=0.55u m=1
.ends labhb2
* SPICE INPUT		Tue Jul 31 19:34:58 2018	labhb3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=labhb3
.subckt labhb3 VDD QN Q GND SN RN D G
M1 N_4 G GND GND mn15  l=0.13u w=0.23u m=1
M2 GND N_4 N_3 GND mn15  l=0.13u w=0.17u m=1
M3 N_5 N_3 N_6 GND mn15  l=0.13u w=0.24u m=1
M4 N_5 N_3 N_6 GND mn15  l=0.13u w=0.24u m=1
M5 N_6 N_3 N_5 GND mn15  l=0.13u w=0.24u m=1
M6 N_34 D N_6 GND mn15  l=0.13u w=0.24u m=1
M7 N_34 D N_6 GND mn15  l=0.13u w=0.24u m=1
M8 N_6 D N_34 GND mn15  l=0.13u w=0.24u m=1
M9 N_37 N_4 N_5 GND mn15  l=0.13u w=0.17u m=1
M10 N_34 RN GND GND mn15  l=0.13u w=0.28u m=1
M11 N_34 RN GND GND mn15  l=0.13u w=0.27u m=1
M12 N_34 RN GND GND mn15  l=0.13u w=0.27u m=1
M13 N_21 SN GND GND mn15  l=0.13u w=0.16u m=1
M14 GND SN N_21 GND mn15  l=0.13u w=0.15u m=1
M15 QN N_27 GND GND mn15  l=0.13u w=0.455u m=1
M16 QN N_27 GND GND mn15  l=0.13u w=0.455u m=1
M17 N_34 N_27 N_37 GND mn15  l=0.13u w=0.17u m=1
M18 QN N_27 GND GND mn15  l=0.13u w=0.43u m=1
M19 GND N_21 N_5 GND mn15  l=0.13u w=0.185u m=1
M20 N_5 N_21 GND GND mn15  l=0.13u w=0.235u m=1
M21 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M22 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M23 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M24 GND N_5 N_27 GND mn15  l=0.13u w=0.39u m=1
M25 N_4 G VDD VDD mp15  l=0.13u w=0.55u m=1
M26 N_3 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M27 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.56u m=1
M28 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.56u m=1
M29 N_6 D N_8 VDD mp15  l=0.13u w=0.29u m=1
M30 N_6 D N_8 VDD mp15  l=0.13u w=0.29u m=1
M31 N_6 D N_8 VDD mp15  l=0.13u w=0.29u m=1
M32 N_6 D N_8 VDD mp15  l=0.13u w=0.29u m=1
M33 N_5 N_3 N_29 VDD mp15  l=0.13u w=0.17u m=1
M34 N_8 RN N_5 VDD mp15  l=0.13u w=0.58u m=1
M35 N_21 SN VDD VDD mp15  l=0.13u w=0.23u m=1
M36 VDD SN N_21 VDD mp15  l=0.13u w=0.23u m=1
M37 QN N_27 VDD VDD mp15  l=0.13u w=0.69u m=1
M38 QN N_27 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 QN N_27 VDD VDD mp15  l=0.13u w=0.69u m=1
M40 N_29 N_27 N_8 VDD mp15  l=0.13u w=0.17u m=1
M41 N_8 N_21 VDD VDD mp15  l=0.13u w=0.46u m=1
M42 N_8 N_21 VDD VDD mp15  l=0.13u w=0.46u m=1
M43 VDD N_21 N_8 VDD mp15  l=0.13u w=0.48u m=1
M44 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M45 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M46 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M47 N_27 N_5 VDD VDD mp15  l=0.13u w=0.58u m=1
.ends labhb3
* SPICE INPUT		Tue Jul 31 19:35:11 2018	lablb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb0
.subckt lablb0 GND Q QN SN D VDD RN GN
M1 N_4 GN GND GND mn15  l=0.13u w=0.17u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 Q N_12 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 N_12 GND GND mn15  l=0.13u w=0.18u m=1
M5 QN N_7 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_10 SN GND GND mn15  l=0.13u w=0.17u m=1
M7 N_18 N_7 N_14 GND mn15  l=0.13u w=0.17u m=1
M8 N_12 N_10 GND GND mn15  l=0.13u w=0.18u m=1
M9 N_18 N_2 N_12 GND mn15  l=0.13u w=0.17u m=1
M10 N_14 RN GND GND mn15  l=0.13u w=0.27u m=1
M11 N_12 N_4 N_15 GND mn15  l=0.13u w=0.27u m=1
M12 N_14 D N_15 GND mn15  l=0.13u w=0.27u m=1
M13 N_4 GN VDD VDD mp15  l=0.13u w=0.42u m=1
M14 VDD N_4 N_2 VDD mp15  l=0.13u w=0.42u m=1
M15 Q N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_7 N_12 VDD VDD mp15  l=0.13u w=0.26u m=1
M17 QN N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_10 SN VDD VDD mp15  l=0.13u w=0.26u m=1
M19 N_20 N_10 VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_20 D N_15 VDD mp15  l=0.13u w=0.42u m=1
M21 N_68 N_7 N_20 VDD mp15  l=0.13u w=0.17u m=1
M22 N_12 N_2 N_15 VDD mp15  l=0.13u w=0.4u m=1
M23 N_12 N_4 N_68 VDD mp15  l=0.13u w=0.17u m=1
M24 N_12 RN N_20 VDD mp15  l=0.13u w=0.3u m=1
.ends lablb0
* SPICE INPUT		Tue Jul 31 19:35:23 2018	lablb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb1
.subckt lablb1 GND Q QN VDD GN D RN SN
M1 N_4 GN GND GND mn15  l=0.13u w=0.17u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_7 N_4 N_5 GND mn15  l=0.13u w=0.37u m=1
M4 N_6 D N_5 GND mn15  l=0.13u w=0.37u m=1
M5 Q N_7 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_10 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M7 N_6 RN GND GND mn15  l=0.13u w=0.4u m=1
M8 N_18 N_2 N_7 GND mn15  l=0.13u w=0.17u m=1
M9 N_18 N_10 N_6 GND mn15  l=0.13u w=0.17u m=1
M10 N_7 N_17 GND GND mn15  l=0.13u w=0.26u m=1
M11 QN N_10 GND GND mn15  l=0.13u w=0.43u m=1
M12 N_17 SN GND GND mn15  l=0.13u w=0.19u m=1
M13 N_4 GN VDD VDD mp15  l=0.13u w=0.42u m=1
M14 VDD N_4 N_2 VDD mp15  l=0.13u w=0.42u m=1
M15 N_25 D N_5 VDD mp15  l=0.13u w=0.51u m=1
M16 N_7 RN N_25 VDD mp15  l=0.13u w=0.37u m=1
M17 N_7 N_4 N_69 VDD mp15  l=0.13u w=0.17u m=1
M18 N_7 N_2 N_5 VDD mp15  l=0.13u w=0.44u m=1
M19 N_7 N_2 N_5 VDD mp15  l=0.13u w=0.44u m=1
M20 N_69 N_10 N_25 VDD mp15  l=0.13u w=0.17u m=1
M21 N_25 N_17 VDD VDD mp15  l=0.13u w=0.62u m=1
M22 QN N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_17 SN VDD VDD mp15  l=0.13u w=0.3u m=1
M24 Q N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_10 N_7 VDD VDD mp15  l=0.13u w=0.36u m=1
.ends lablb1
* SPICE INPUT		Tue Jul 31 19:35:36 2018	lablb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb2
.subckt lablb2 GND QN Q D VDD SN RN GN
M1 N_4 GN GND GND mn15  l=0.13u w=0.22u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.22u m=1
M3 N_7 RN GND GND mn15  l=0.13u w=0.36u m=1
M4 N_7 RN GND GND mn15  l=0.13u w=0.36u m=1
M5 N_23 N_2 N_5 GND mn15  l=0.13u w=0.17u m=1
M6 N_7 N_21 N_23 GND mn15  l=0.13u w=0.17u m=1
M7 N_7 D N_9 GND mn15  l=0.13u w=0.72u m=1
M8 N_5 N_4 N_9 GND mn15  l=0.13u w=0.63u m=1
M9 GND N_17 N_5 GND mn15  l=0.13u w=0.185u m=1
M10 N_5 N_17 GND GND mn15  l=0.13u w=0.185u m=1
M11 GND SN N_17 GND mn15  l=0.13u w=0.185u m=1
M12 N_17 SN GND GND mn15  l=0.13u w=0.185u m=1
M13 GND N_21 QN GND mn15  l=0.13u w=0.455u m=1
M14 GND N_21 QN GND mn15  l=0.13u w=0.435u m=1
M15 GND N_5 Q GND mn15  l=0.13u w=0.46u m=1
M16 GND N_5 Q GND mn15  l=0.13u w=0.46u m=1
M17 GND N_5 N_21 GND mn15  l=0.13u w=0.36u m=1
M18 N_4 GN VDD VDD mp15  l=0.13u w=0.55u m=1
M19 VDD N_4 N_2 VDD mp15  l=0.13u w=0.55u m=1
M20 N_5 RN N_28 VDD mp15  l=0.13u w=0.27u m=1
M21 N_5 RN N_28 VDD mp15  l=0.13u w=0.27u m=1
M22 N_88 N_4 N_5 VDD mp15  l=0.13u w=0.17u m=1
M23 N_28 N_21 N_88 VDD mp15  l=0.13u w=0.17u m=1
M24 N_9 D N_28 VDD mp15  l=0.13u w=0.63u m=1
M25 N_9 D N_28 VDD mp15  l=0.13u w=0.63u m=1
M26 N_5 N_2 N_9 VDD mp15  l=0.13u w=1.25u m=1
M27 N_28 N_17 VDD VDD mp15  l=0.13u w=0.63u m=1
M28 VDD N_17 N_28 VDD mp15  l=0.13u w=0.63u m=1
M29 N_17 SN VDD VDD mp15  l=0.13u w=0.55u m=1
M30 VDD N_21 QN VDD mp15  l=0.13u w=0.69u m=1
M31 QN N_21 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 VDD N_5 Q VDD mp15  l=0.13u w=0.69u m=1
M33 VDD N_5 Q VDD mp15  l=0.13u w=0.69u m=1
M34 N_21 N_5 VDD VDD mp15  l=0.13u w=0.52u m=1
.ends lablb2
* SPICE INPUT		Tue Jul 31 19:35:49 2018	lablb3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lablb3
.subckt lablb3 GND Q QN D VDD GN SN RN
M1 Q N_14 GND GND mn15  l=0.13u w=0.46u m=1
M2 Q N_14 GND GND mn15  l=0.13u w=0.46u m=1
M3 Q N_14 GND GND mn15  l=0.13u w=0.46u m=1
M4 GND N_14 N_5 GND mn15  l=0.13u w=0.285u m=1
M5 N_5 N_14 GND GND mn15  l=0.13u w=0.285u m=1
M6 N_10 GN GND GND mn15  l=0.13u w=0.27u m=1
M7 N_9 N_10 GND GND mn15  l=0.13u w=0.27u m=1
M8 QN N_5 GND GND mn15  l=0.13u w=0.455u m=1
M9 QN N_5 GND GND mn15  l=0.13u w=0.455u m=1
M10 QN N_5 GND GND mn15  l=0.13u w=0.43u m=1
M11 GND SN N_16 GND mn15  l=0.13u w=0.185u m=1
M12 N_16 SN GND GND mn15  l=0.13u w=0.185u m=1
M13 GND N_16 N_14 GND mn15  l=0.13u w=0.23u m=1
M14 N_14 N_16 GND GND mn15  l=0.13u w=0.23u m=1
M15 N_14 N_10 N_19 GND mn15  l=0.13u w=0.74u m=1
M16 N_20 D N_19 GND mn15  l=0.13u w=0.85u m=1
M17 N_20 N_5 N_26 GND mn15  l=0.13u w=0.17u m=1
M18 N_26 N_9 N_14 GND mn15  l=0.13u w=0.17u m=1
M19 N_20 RN GND GND mn15  l=0.13u w=0.425u m=1
M20 N_20 RN GND GND mn15  l=0.13u w=0.425u m=1
M21 QN N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 QN N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 QN N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_16 SN VDD VDD mp15  l=0.13u w=0.56u m=1
M25 N_31 N_16 VDD VDD mp15  l=0.13u w=0.63u m=1
M26 VDD N_16 N_31 VDD mp15  l=0.13u w=0.63u m=1
M27 N_31 N_5 N_100 VDD mp15  l=0.13u w=0.17u m=1
M28 N_14 RN N_31 VDD mp15  l=0.13u w=0.315u m=1
M29 N_14 RN N_31 VDD mp15  l=0.13u w=0.315u m=1
M30 N_100 N_10 N_14 VDD mp15  l=0.13u w=0.17u m=1
M31 N_10 GN VDD VDD mp15  l=0.13u w=0.67u m=1
M32 VDD N_10 N_9 VDD mp15  l=0.13u w=0.67u m=1
M33 Q N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M34 Q N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 Q N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 N_5 N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M37 N_5 N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M38 N_14 N_9 N_19 VDD mp15  l=0.13u w=1.34u m=1
M39 N_19 D N_31 VDD mp15  l=0.13u w=0.67u m=1
M40 N_19 D N_31 VDD mp15  l=0.13u w=0.67u m=1
.ends lablb3
* SPICE INPUT		Tue Jul 31 19:36:02 2018	lachb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb0
.subckt lachb0 GND QN Q VDD RN D G
M1 N_4 G GND GND mn15  l=0.13u w=0.17u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_7 N_2 N_5 GND mn15  l=0.13u w=0.18u m=1
M4 N_15 D N_7 GND mn15  l=0.13u w=0.18u m=1
M5 N_15 RN GND GND mn15  l=0.13u w=0.18u m=1
M6 N_16 RN GND GND mn15  l=0.13u w=0.17u m=1
M7 N_14 N_4 N_5 GND mn15  l=0.13u w=0.17u m=1
M8 N_16 N_13 N_14 GND mn15  l=0.13u w=0.17u m=1
M9 QN N_13 GND GND mn15  l=0.13u w=0.26u m=1
M10 Q N_5 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_13 N_5 GND GND mn15  l=0.13u w=0.18u m=1
M12 N_4 G VDD VDD mp15  l=0.13u w=0.42u m=1
M13 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M14 N_7 D VDD VDD mp15  l=0.13u w=0.37u m=1
M15 N_5 RN VDD VDD mp15  l=0.13u w=0.22u m=1
M16 N_25 N_2 N_5 VDD mp15  l=0.13u w=0.17u m=1
M17 N_7 N_4 N_5 VDD mp15  l=0.13u w=0.28u m=1
M18 N_25 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 QN N_13 VDD VDD mp15  l=0.13u w=0.4u m=1
M20 Q N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_13 N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends lachb0
* SPICE INPUT		Tue Jul 31 19:36:15 2018	lachb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb1
.subckt lachb1 GND Q QN VDD G RN D
M1 N_4 G GND GND mn15  l=0.13u w=0.17u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_7 N_2 N_5 GND mn15  l=0.13u w=0.28u m=1
M4 N_15 D N_7 GND mn15  l=0.13u w=0.37u m=1
M5 N_15 RN GND GND mn15  l=0.13u w=0.37u m=1
M6 N_16 RN GND GND mn15  l=0.13u w=0.17u m=1
M7 N_14 N_4 N_5 GND mn15  l=0.13u w=0.17u m=1
M8 N_16 N_11 N_14 GND mn15  l=0.13u w=0.17u m=1
M9 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_11 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M11 QN N_11 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_4 G VDD VDD mp15  l=0.13u w=0.42u m=1
M13 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M14 N_7 D VDD VDD mp15  l=0.13u w=0.47u m=1
M15 N_5 RN VDD VDD mp15  l=0.13u w=0.37u m=1
M16 N_26 N_2 N_5 VDD mp15  l=0.13u w=0.17u m=1
M17 N_7 N_4 N_5 VDD mp15  l=0.13u w=0.42u m=1
M18 N_26 N_11 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 QN N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_11 N_5 VDD VDD mp15  l=0.13u w=0.37u m=1
.ends lachb1
* SPICE INPUT		Tue Jul 31 19:36:29 2018	lachb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb2
.subckt lachb2 GND QN Q VDD RN D G
M1 N_4 G GND GND mn15  l=0.13u w=0.17u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_6 N_2 N_5 GND mn15  l=0.13u w=0.225u m=1
M4 N_5 N_2 N_6 GND mn15  l=0.13u w=0.225u m=1
M5 N_17 D N_6 GND mn15  l=0.13u w=0.46u m=1
M6 N_17 RN GND GND mn15  l=0.13u w=0.46u m=1
M7 N_18 RN GND GND mn15  l=0.13u w=0.17u m=1
M8 N_16 N_4 N_5 GND mn15  l=0.13u w=0.17u m=1
M9 N_18 N_12 N_16 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_5 Q GND mn15  l=0.13u w=0.46u m=1
M11 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M12 GND N_5 N_12 GND mn15  l=0.13u w=0.36u m=1
M13 GND N_12 QN GND mn15  l=0.13u w=0.46u m=1
M14 GND N_12 QN GND mn15  l=0.13u w=0.46u m=1
M15 N_4 G VDD VDD mp15  l=0.13u w=0.42u m=1
M16 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M17 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.315u m=1
M18 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.315u m=1
M19 N_6 D VDD VDD mp15  l=0.13u w=0.63u m=1
M20 N_5 RN VDD VDD mp15  l=0.13u w=0.5u m=1
M21 N_5 N_2 N_29 VDD mp15  l=0.13u w=0.17u m=1
M22 N_29 N_12 VDD VDD mp15  l=0.13u w=0.17u m=1
M23 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_12 N_5 VDD VDD mp15  l=0.13u w=0.52u m=1
M26 VDD N_12 QN VDD mp15  l=0.13u w=0.69u m=1
M27 VDD N_12 QN VDD mp15  l=0.13u w=0.69u m=1
.ends lachb2
* SPICE INPUT		Tue Jul 31 19:36:42 2018	lachb3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lachb3
.subckt lachb3 GND QN Q VDD RN D G
M1 N_4 G GND GND mn15  l=0.13u w=0.17u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_23 D N_5 GND mn15  l=0.13u w=0.27u m=1
M4 N_5 D N_22 GND mn15  l=0.13u w=0.27u m=1
M5 N_21 D N_5 GND mn15  l=0.13u w=0.26u m=1
M6 N_22 RN GND GND mn15  l=0.13u w=0.27u m=1
M7 N_23 RN GND GND mn15  l=0.13u w=0.27u m=1
M8 N_21 RN GND GND mn15  l=0.13u w=0.26u m=1
M9 N_24 RN GND GND mn15  l=0.13u w=0.17u m=1
M10 N_25 N_4 N_6 GND mn15  l=0.13u w=0.17u m=1
M11 N_6 N_2 N_5 GND mn15  l=0.13u w=0.27u m=1
M12 N_6 N_2 N_5 GND mn15  l=0.13u w=0.27u m=1
M13 N_25 N_18 N_24 GND mn15  l=0.13u w=0.17u m=1
M14 QN N_18 GND GND mn15  l=0.13u w=0.46u m=1
M15 QN N_18 GND GND mn15  l=0.13u w=0.46u m=1
M16 QN N_18 GND GND mn15  l=0.13u w=0.46u m=1
M17 Q N_6 GND GND mn15  l=0.13u w=0.46u m=1
M18 GND N_6 N_18 GND mn15  l=0.13u w=0.46u m=1
M19 Q N_6 GND GND mn15  l=0.13u w=0.46u m=1
M20 Q N_6 GND GND mn15  l=0.13u w=0.46u m=1
M21 N_4 G VDD VDD mp15  l=0.13u w=0.42u m=1
M22 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M23 N_5 D VDD VDD mp15  l=0.13u w=0.31u m=1
M24 N_5 D VDD VDD mp15  l=0.13u w=0.31u m=1
M25 VDD D N_5 VDD mp15  l=0.13u w=0.31u m=1
M26 N_5 D VDD VDD mp15  l=0.13u w=0.31u m=1
M27 N_6 RN VDD VDD mp15  l=0.13u w=0.31u m=1
M28 VDD RN N_6 VDD mp15  l=0.13u w=0.31u m=1
M29 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.31u m=1
M30 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.32u m=1
M31 N_97 N_2 N_6 VDD mp15  l=0.13u w=0.17u m=1
M32 QN N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M33 QN N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M34 QN N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 N_97 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M36 Q N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M37 Q N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M38 Q N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 N_18 N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends lachb3
* SPICE INPUT		Tue Jul 31 19:36:56 2018	laclb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb0
.subckt laclb0 GND QN Q VDD RN D GN
M1 N_4 GN GND GND mn15  l=0.13u w=0.17u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_7 N_4 N_5 GND mn15  l=0.13u w=0.17u m=1
M4 N_15 D N_7 GND mn15  l=0.13u w=0.26u m=1
M5 N_15 RN GND GND mn15  l=0.13u w=0.26u m=1
M6 N_16 RN GND GND mn15  l=0.13u w=0.17u m=1
M7 N_14 N_2 N_5 GND mn15  l=0.13u w=0.17u m=1
M8 N_16 N_13 N_14 GND mn15  l=0.13u w=0.17u m=1
M9 QN N_13 GND GND mn15  l=0.13u w=0.26u m=1
M10 Q N_5 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_13 N_5 GND GND mn15  l=0.13u w=0.18u m=1
M12 Q N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_13 N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
M14 N_4 GN VDD VDD mp15  l=0.13u w=0.42u m=1
M15 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M16 N_7 D VDD VDD mp15  l=0.13u w=0.38u m=1
M17 N_26 N_4 N_5 VDD mp15  l=0.13u w=0.17u m=1
M18 N_5 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M19 N_7 N_2 N_5 VDD mp15  l=0.13u w=0.17u m=1
M20 N_26 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M21 QN N_13 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends laclb0
* SPICE INPUT		Tue Jul 31 19:37:09 2018	laclb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb1
.subckt laclb1 GND QN Q RN D VDD GN
M1 N_4 GN GND GND mn15  l=0.13u w=0.17u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_7 N_4 N_5 GND mn15  l=0.13u w=0.28u m=1
M4 N_15 D N_7 GND mn15  l=0.13u w=0.37u m=1
M5 N_15 RN GND GND mn15  l=0.13u w=0.37u m=1
M6 N_16 RN GND GND mn15  l=0.13u w=0.17u m=1
M7 N_14 N_2 N_5 GND mn15  l=0.13u w=0.17u m=1
M8 N_16 N_13 N_14 GND mn15  l=0.13u w=0.17u m=1
M9 QN N_13 GND GND mn15  l=0.13u w=0.46u m=1
M10 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_13 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M12 N_4 GN VDD VDD mp15  l=0.13u w=0.42u m=1
M13 N_2 N_4 VDD VDD mp15  l=0.13u w=0.42u m=1
M14 VDD D N_7 VDD mp15  l=0.13u w=0.39u m=1
M15 N_5 RN VDD VDD mp15  l=0.13u w=0.37u m=1
M16 N_5 N_4 N_25 VDD mp15  l=0.13u w=0.17u m=1
M17 N_5 N_2 N_7 VDD mp15  l=0.13u w=0.42u m=1
M18 N_25 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 QN N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_13 N_5 VDD VDD mp15  l=0.13u w=0.37u m=1
.ends laclb1
* SPICE INPUT		Tue Jul 31 19:37:23 2018	laclb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb2
.subckt laclb2 GND QN Q VDD RN D GN
M1 N_4 GN GND GND mn15  l=0.13u w=0.2u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.17u m=1
M3 N_5 N_4 N_6 GND mn15  l=0.13u w=0.41u m=1
M4 N_16 D N_6 GND mn15  l=0.13u w=0.46u m=1
M5 N_16 RN GND GND mn15  l=0.13u w=0.46u m=1
M6 N_17 RN GND GND mn15  l=0.13u w=0.17u m=1
M7 N_15 N_2 N_5 GND mn15  l=0.13u w=0.17u m=1
M8 N_17 N_11 N_15 GND mn15  l=0.13u w=0.17u m=1
M9 GND N_5 Q GND mn15  l=0.13u w=0.46u m=1
M10 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_5 N_11 GND mn15  l=0.13u w=0.37u m=1
M12 GND N_11 QN GND mn15  l=0.13u w=0.46u m=1
M13 GND N_11 QN GND mn15  l=0.13u w=0.46u m=1
M14 N_4 GN VDD VDD mp15  l=0.13u w=0.51u m=1
M15 VDD N_4 N_2 VDD mp15  l=0.13u w=0.42u m=1
M16 N_5 N_2 N_6 VDD mp15  l=0.13u w=0.59u m=1
M17 VDD D N_6 VDD mp15  l=0.13u w=0.56u m=1
M18 N_5 RN VDD VDD mp15  l=0.13u w=0.54u m=1
M19 N_5 N_4 N_27 VDD mp15  l=0.13u w=0.17u m=1
M20 N_27 N_11 VDD VDD mp15  l=0.13u w=0.17u m=1
M21 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_11 N_5 VDD VDD mp15  l=0.13u w=0.55u m=1
M24 VDD N_11 QN VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_11 QN VDD mp15  l=0.13u w=0.69u m=1
.ends laclb2
* SPICE INPUT		Tue Jul 31 19:37:36 2018	laclb3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laclb3
.subckt laclb3 GND QN Q VDD RN D GN
M1 N_4 GN GND GND mn15  l=0.13u w=0.2u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.2u m=1
M3 N_22 D N_5 GND mn15  l=0.13u w=0.49u m=1
M4 N_5 D N_21 GND mn15  l=0.13u w=0.27u m=1
M5 N_22 RN GND GND mn15  l=0.13u w=0.49u m=1
M6 GND RN N_21 GND mn15  l=0.13u w=0.27u m=1
M7 N_23 RN GND GND mn15  l=0.13u w=0.17u m=1
M8 N_24 N_2 N_8 GND mn15  l=0.13u w=0.17u m=1
M9 N_8 N_4 N_5 GND mn15  l=0.13u w=0.26u m=1
M10 N_5 N_4 N_8 GND mn15  l=0.13u w=0.19u m=1
M11 N_24 N_18 N_23 GND mn15  l=0.13u w=0.17u m=1
M12 QN N_18 GND GND mn15  l=0.13u w=0.46u m=1
M13 QN N_18 GND GND mn15  l=0.13u w=0.46u m=1
M14 QN N_18 GND GND mn15  l=0.13u w=0.46u m=1
M15 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M16 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M17 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M18 GND N_8 N_18 GND mn15  l=0.13u w=0.41u m=1
M19 N_4 GN VDD VDD mp15  l=0.13u w=0.51u m=1
M20 N_2 N_4 VDD VDD mp15  l=0.13u w=0.51u m=1
M21 N_5 D VDD VDD mp15  l=0.13u w=0.23u m=1
M22 VDD D N_5 VDD mp15  l=0.13u w=0.23u m=1
M23 VDD D N_5 VDD mp15  l=0.13u w=0.24u m=1
M24 N_8 RN VDD VDD mp15  l=0.13u w=0.31u m=1
M25 VDD RN N_8 VDD mp15  l=0.13u w=0.31u m=1
M26 N_5 N_2 N_8 VDD mp15  l=0.13u w=0.32u m=1
M27 N_5 N_2 N_8 VDD mp15  l=0.13u w=0.32u m=1
M28 N_91 N_4 N_8 VDD mp15  l=0.13u w=0.17u m=1
M29 QN N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 QN N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 QN N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 N_91 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M33 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M34 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 N_18 N_8 VDD VDD mp15  l=0.13u w=0.63u m=1
.ends laclb3
* SPICE INPUT		Tue Jul 31 19:37:49 2018	lanhb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb0
.subckt lanhb0 VDD QN Q G GND D
M1 N_19 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_19 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 N_20 N_10 N_6 GND mn15  l=0.13u w=0.17u m=1
M4 GND N_10 N_5 GND mn15  l=0.13u w=0.17u m=1
M5 QN N_9 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_20 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M7 Q N_6 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_9 N_6 GND GND mn15  l=0.13u w=0.18u m=1
M9 GND G N_10 GND mn15  l=0.13u w=0.17u m=1
M10 N_12 D VDD VDD mp15  l=0.13u w=0.33u m=1
M11 N_13 N_5 N_6 VDD mp15  l=0.13u w=0.17u m=1
M12 N_5 N_10 VDD VDD mp15  l=0.13u w=0.42u m=1
M13 N_12 N_10 N_6 VDD mp15  l=0.13u w=0.33u m=1
M14 N_13 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M15 QN N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 Q N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_9 N_6 VDD VDD mp15  l=0.13u w=0.26u m=1
M18 VDD G N_10 VDD mp15  l=0.13u w=0.42u m=1
.ends lanhb0
* SPICE INPUT		Tue Jul 31 19:38:02 2018	lanhb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb1
.subckt lanhb1 GND QN Q VDD D G
M1 GND G N_2 GND mn15  l=0.13u w=0.2u m=1
M2 N_12 D GND GND mn15  l=0.13u w=0.28u m=1
M3 N_12 N_6 N_8 GND mn15  l=0.13u w=0.28u m=1
M4 GND N_2 N_6 GND mn15  l=0.13u w=0.2u m=1
M5 N_13 N_2 N_8 GND mn15  l=0.13u w=0.17u m=1
M6 QN N_11 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_13 N_11 GND GND mn15  l=0.13u w=0.17u m=1
M8 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M9 N_11 N_8 GND GND mn15  l=0.13u w=0.28u m=1
M10 VDD G N_2 VDD mp15  l=0.13u w=0.51u m=1
M11 N_21 D VDD VDD mp15  l=0.13u w=0.42u m=1
M12 N_22 N_6 N_8 VDD mp15  l=0.13u w=0.17u m=1
M13 N_6 N_2 VDD VDD mp15  l=0.13u w=0.51u m=1
M14 N_21 N_2 N_8 VDD mp15  l=0.13u w=0.42u m=1
M15 QN N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_22 N_11 VDD VDD mp15  l=0.13u w=0.17u m=1
M17 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_11 N_8 VDD VDD mp15  l=0.13u w=0.41u m=1
.ends lanhb1
* SPICE INPUT		Tue Jul 31 19:38:14 2018	lanhb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb2
.subckt lanhb2 VDD QN Q G D GND
M1 GND N_3 N_13 GND mn15  l=0.13u w=0.17u m=1
M2 N_64 N_3 N_6 GND mn15  l=0.13u w=0.17u m=1
M3 N_63 D GND GND mn15  l=0.13u w=0.27u m=1
M4 N_63 N_13 N_6 GND mn15  l=0.13u w=0.27u m=1
M5 N_6 N_13 N_62 GND mn15  l=0.13u w=0.27u m=1
M6 N_62 D GND GND mn15  l=0.13u w=0.27u m=1
M7 QN N_5 GND GND mn15  l=0.13u w=0.46u m=1
M8 QN N_5 GND GND mn15  l=0.13u w=0.46u m=1
M9 N_64 N_5 GND GND mn15  l=0.13u w=0.17u m=1
M10 Q N_6 GND GND mn15  l=0.13u w=0.46u m=1
M11 Q N_6 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_5 N_6 GND GND mn15  l=0.13u w=0.36u m=1
M13 GND G N_3 GND mn15  l=0.13u w=0.2u m=1
M14 N_3 G VDD VDD mp15  l=0.13u w=0.46u m=1
M15 N_15 N_13 N_6 VDD mp15  l=0.13u w=0.17u m=1
M16 QN N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 QN N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_15 N_5 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 Q N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Q N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_5 N_6 VDD VDD mp15  l=0.13u w=0.52u m=1
M22 N_13 N_3 VDD VDD mp15  l=0.13u w=0.42u m=1
M23 N_6 N_3 N_17 VDD mp15  l=0.13u w=0.405u m=1
M24 N_6 N_3 N_16 VDD mp15  l=0.13u w=0.405u m=1
M25 N_16 D VDD VDD mp15  l=0.13u w=0.405u m=1
M26 N_17 D VDD VDD mp15  l=0.13u w=0.405u m=1
.ends lanhb2
* SPICE INPUT		Tue Jul 31 19:38:28 2018	lanhb3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanhb3
.subckt lanhb3 GND Q QN VDD D G
M1 Q N_11 GND GND mn15  l=0.13u w=0.46u m=1
M2 Q N_11 GND GND mn15  l=0.13u w=0.46u m=1
M3 Q N_11 GND GND mn15  l=0.13u w=0.46u m=1
M4 GND N_11 N_4 GND mn15  l=0.13u w=0.38u m=1
M5 QN N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 QN N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 QN N_4 GND GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 N_21 GND mn15  l=0.13u w=0.17u m=1
M9 GND N_16 N_9 GND mn15  l=0.13u w=0.17u m=1
M10 N_18 D GND GND mn15  l=0.13u w=0.28u m=1
M11 N_19 D GND GND mn15  l=0.13u w=0.28u m=1
M12 N_20 D GND GND mn15  l=0.13u w=0.26u m=1
M13 N_21 N_16 N_11 GND mn15  l=0.13u w=0.17u m=1
M14 N_20 N_9 N_11 GND mn15  l=0.13u w=0.26u m=1
M15 N_11 N_9 N_18 GND mn15  l=0.13u w=0.28u m=1
M16 N_19 N_9 N_11 GND mn15  l=0.13u w=0.28u m=1
M17 GND G N_16 GND mn15  l=0.13u w=0.22u m=1
M18 N_16 G VDD VDD mp15  l=0.13u w=0.55u m=1
M19 Q N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Q N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 Q N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_4 N_11 VDD VDD mp15  l=0.13u w=0.57u m=1
M23 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_37 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_36 N_16 N_11 VDD mp15  l=0.13u w=0.41u m=1
M28 N_35 N_16 N_11 VDD mp15  l=0.13u w=0.42u m=1
M29 N_11 N_16 N_34 VDD mp15  l=0.13u w=0.42u m=1
M30 VDD N_16 N_9 VDD mp15  l=0.13u w=0.42u m=1
M31 N_34 D VDD VDD mp15  l=0.13u w=0.42u m=1
M32 N_35 D VDD VDD mp15  l=0.13u w=0.42u m=1
M33 N_36 D VDD VDD mp15  l=0.13u w=0.41u m=1
M34 N_37 N_9 N_11 VDD mp15  l=0.13u w=0.17u m=1
.ends lanhb3
* SPICE INPUT		Tue Jul 31 19:38:41 2018	lanlb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb0
.subckt lanlb0 VDD QN Q GN D GND
M1 GND N_11 N_5 GND mn15  l=0.13u w=0.17u m=1
M2 N_19 D GND GND mn15  l=0.13u w=0.18u m=1
M3 N_19 N_11 N_6 GND mn15  l=0.13u w=0.18u m=1
M4 N_20 N_5 N_6 GND mn15  l=0.13u w=0.17u m=1
M5 QN N_9 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_20 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M7 Q N_6 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_9 N_6 GND GND mn15  l=0.13u w=0.18u m=1
M9 GND GN N_11 GND mn15  l=0.13u w=0.17u m=1
M10 N_5 N_11 VDD VDD mp15  l=0.13u w=0.42u m=1
M11 N_12 D VDD VDD mp15  l=0.13u w=0.37u m=1
M12 N_12 N_5 N_6 VDD mp15  l=0.13u w=0.37u m=1
M13 N_13 N_11 N_6 VDD mp15  l=0.13u w=0.17u m=1
M14 QN N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M15 N_13 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M16 Q N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_9 N_6 VDD VDD mp15  l=0.13u w=0.26u m=1
M18 N_11 GN VDD VDD mp15  l=0.13u w=0.42u m=1
.ends lanlb0
* SPICE INPUT		Tue Jul 31 19:38:54 2018	lanlb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb1
.subckt lanlb1 GND Q QN VDD GN D
M1 Q N_11 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 N_11 GND GND mn15  l=0.13u w=0.27u m=1
M3 GND GN N_5 GND mn15  l=0.13u w=0.17u m=1
M4 GND N_5 N_9 GND mn15  l=0.13u w=0.17u m=1
M5 N_12 D GND GND mn15  l=0.13u w=0.38u m=1
M6 N_12 N_5 N_11 GND mn15  l=0.13u w=0.38u m=1
M7 QN N_4 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_13 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_13 N_9 N_11 GND mn15  l=0.13u w=0.17u m=1
M10 N_5 GN VDD VDD mp15  l=0.13u w=0.44u m=1
M11 VDD N_5 N_9 VDD mp15  l=0.13u w=0.42u m=1
M12 N_21 D VDD VDD mp15  l=0.13u w=0.57u m=1
M13 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_22 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M15 N_22 N_5 N_11 VDD mp15  l=0.13u w=0.17u m=1
M16 N_21 N_9 N_11 VDD mp15  l=0.13u w=0.57u m=1
M17 Q N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_4 N_11 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends lanlb1
* SPICE INPUT		Tue Jul 31 19:39:07 2018	lanlb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb2
.subckt lanlb2 GND QN Q VDD D GN
M1 N_3 GN GND GND mn15  l=0.13u w=0.27u m=1
M2 GND N_13 QN GND mn15  l=0.13u w=0.46u m=1
M3 GND N_13 QN GND mn15  l=0.13u w=0.46u m=1
M4 N_17 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_15 D GND GND mn15  l=0.13u w=0.33u m=1
M6 N_16 N_3 N_8 GND mn15  l=0.13u w=0.36u m=1
M7 N_8 N_3 N_15 GND mn15  l=0.13u w=0.33u m=1
M8 GND N_3 N_6 GND mn15  l=0.13u w=0.17u m=1
M9 N_16 D GND GND mn15  l=0.13u w=0.36u m=1
M10 N_17 N_6 N_8 GND mn15  l=0.13u w=0.17u m=1
M11 GND N_8 Q GND mn15  l=0.13u w=0.455u m=1
M12 GND N_8 Q GND mn15  l=0.13u w=0.455u m=1
M13 GND N_8 N_13 GND mn15  l=0.13u w=0.37u m=1
M14 N_3 GN VDD VDD mp15  l=0.13u w=0.67u m=1
M15 VDD N_13 QN VDD mp15  l=0.13u w=0.69u m=1
M16 QN N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_73 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M18 N_70 D VDD VDD mp15  l=0.13u w=0.355u m=1
M19 N_71 N_6 N_8 VDD mp15  l=0.13u w=0.355u m=1
M20 N_8 N_6 N_70 VDD mp15  l=0.13u w=0.355u m=1
M21 N_6 N_3 VDD VDD mp15  l=0.13u w=0.42u m=1
M22 N_72 D VDD VDD mp15  l=0.13u w=0.36u m=1
M23 VDD D N_71 VDD mp15  l=0.13u w=0.355u m=1
M24 N_8 N_6 N_72 VDD mp15  l=0.13u w=0.36u m=1
M25 N_73 N_3 N_8 VDD mp15  l=0.13u w=0.17u m=1
M26 VDD N_8 Q VDD mp15  l=0.13u w=0.69u m=1
M27 VDD N_8 Q VDD mp15  l=0.13u w=0.69u m=1
M28 N_13 N_8 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends lanlb2
* SPICE INPUT		Tue Jul 31 19:39:20 2018	lanlb3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=lanlb3
.subckt lanlb3 GND QN Q VDD GN D
M1 N_3 GN GND GND mn15  l=0.13u w=0.27u m=1
M2 N_18 D GND GND mn15  l=0.13u w=0.31u m=1
M3 N_19 N_3 N_8 GND mn15  l=0.13u w=0.31u m=1
M4 N_8 N_3 N_18 GND mn15  l=0.13u w=0.31u m=1
M5 GND N_3 N_6 GND mn15  l=0.13u w=0.2u m=1
M6 N_19 D GND GND mn15  l=0.13u w=0.31u m=1
M7 N_20 D GND GND mn15  l=0.13u w=0.28u m=1
M8 QN N_15 GND GND mn15  l=0.13u w=0.46u m=1
M9 QN N_15 GND GND mn15  l=0.13u w=0.46u m=1
M10 QN N_15 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_15 N_21 GND mn15  l=0.13u w=0.17u m=1
M12 N_8 N_3 N_20 GND mn15  l=0.13u w=0.28u m=1
M13 N_21 N_6 N_8 GND mn15  l=0.13u w=0.17u m=1
M14 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M15 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M16 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M17 GND N_8 N_15 GND mn15  l=0.13u w=0.45u m=1
M18 N_3 GN VDD VDD mp15  l=0.13u w=0.67u m=1
M19 N_83 D VDD VDD mp15  l=0.13u w=0.37u m=1
M20 N_84 N_6 N_8 VDD mp15  l=0.13u w=0.37u m=1
M21 N_8 N_6 N_83 VDD mp15  l=0.13u w=0.37u m=1
M22 N_6 N_3 VDD VDD mp15  l=0.13u w=0.51u m=1
M23 N_85 D VDD VDD mp15  l=0.13u w=0.6u m=1
M24 N_84 D VDD VDD mp15  l=0.13u w=0.37u m=1
M25 QN N_15 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 QN N_15 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 QN N_15 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 N_86 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_85 N_6 N_8 VDD mp15  l=0.13u w=0.6u m=1
M30 N_86 N_3 N_8 VDD mp15  l=0.13u w=0.17u m=1
M31 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M33 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M34 N_15 N_8 VDD VDD mp15  l=0.13u w=0.66u m=1
.ends lanlb3
* SPICE INPUT		Tue Jul 31 19:39:33 2018	laphb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb0
.subckt laphb0 VDD Q QN SN D GND G
M1 Q N_14 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 N_14 GND GND mn15  l=0.13u w=0.18u m=1
M3 QN N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 G GND GND mn15  l=0.13u w=0.17u m=1
M5 N_62 N_7 N_14 GND mn15  l=0.13u w=0.17u m=1
M6 GND N_7 N_10 GND mn15  l=0.13u w=0.17u m=1
M7 N_62 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_14 N_10 N_13 GND mn15  l=0.13u w=0.28u m=1
M9 N_13 D GND GND mn15  l=0.13u w=0.18u m=1
M10 GND N_9 N_14 GND mn15  l=0.13u w=0.18u m=1
M11 GND SN N_9 GND mn15  l=0.13u w=0.18u m=1
M12 Q N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_4 N_14 VDD VDD mp15  l=0.13u w=0.26u m=1
M14 VDD N_4 QN VDD mp15  l=0.13u w=0.4u m=1
M15 N_7 G VDD VDD mp15  l=0.13u w=0.42u m=1
M16 N_9 SN VDD VDD mp15  l=0.13u w=0.26u m=1
M17 VDD N_7 N_10 VDD mp15  l=0.13u w=0.42u m=1
M18 N_14 N_7 N_13 VDD mp15  l=0.13u w=0.28u m=1
M19 N_17 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M20 N_17 N_4 N_16 VDD mp15  l=0.13u w=0.17u m=1
M21 N_16 N_10 N_14 VDD mp15  l=0.13u w=0.17u m=1
M22 N_15 D N_13 VDD mp15  l=0.13u w=0.48u m=1
M23 N_15 N_9 VDD VDD mp15  l=0.13u w=0.48u m=1
.ends laphb0
* SPICE INPUT		Tue Jul 31 19:39:45 2018	laphb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb1
.subckt laphb1 GND Q QN SN D VDD G
M1 N_3 SN GND GND mn15  l=0.13u w=0.28u m=1
M2 GND N_3 N_6 GND mn15  l=0.13u w=0.28u m=1
M3 N_9 D GND GND mn15  l=0.13u w=0.28u m=1
M4 N_9 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_17 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M6 GND N_11 N_4 GND mn15  l=0.13u w=0.2u m=1
M7 N_17 N_11 N_6 GND mn15  l=0.13u w=0.17u m=1
M8 N_11 G GND GND mn15  l=0.13u w=0.2u m=1
M9 Q N_6 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_14 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M11 QN N_14 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_3 SN VDD VDD mp15  l=0.13u w=0.41u m=1
M13 N_63 N_3 VDD VDD mp15  l=0.13u w=0.7u m=1
M14 N_63 D N_9 VDD mp15  l=0.13u w=0.7u m=1
M15 N_64 N_4 N_6 VDD mp15  l=0.13u w=0.17u m=1
M16 N_65 N_14 N_64 VDD mp15  l=0.13u w=0.17u m=1
M17 N_65 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M18 VDD N_11 N_4 VDD mp15  l=0.13u w=0.51u m=1
M19 N_6 N_11 N_9 VDD mp15  l=0.13u w=0.41u m=1
M20 N_11 G VDD VDD mp15  l=0.13u w=0.51u m=1
M21 Q N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_14 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M23 QN N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends laphb1
* SPICE INPUT		Tue Jul 31 19:39:58 2018	laphb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb2
.subckt laphb2 QN GND Q D G SN VDD
M1 GND N_13 Q GND mn15  l=0.13u w=0.46u m=1
M2 Q N_13 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND N_13 N_4 GND mn15  l=0.13u w=0.37u m=1
M4 GND N_4 QN GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 QN GND mn15  l=0.13u w=0.46u m=1
M6 N_9 G GND GND mn15  l=0.13u w=0.17u m=1
M7 N_18 N_9 N_13 GND mn15  l=0.13u w=0.17u m=1
M8 GND N_9 N_10 GND mn15  l=0.13u w=0.17u m=1
M9 N_18 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M10 N_13 N_10 N_14 GND mn15  l=0.13u w=0.37u m=1
M11 N_14 D GND GND mn15  l=0.13u w=0.37u m=1
M12 N_13 N_17 GND GND mn15  l=0.13u w=0.37u m=1
M13 N_17 SN GND GND mn15  l=0.13u w=0.28u m=1
M14 Q N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 Q N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_4 N_13 VDD VDD mp15  l=0.13u w=0.55u m=1
M17 VDD N_4 QN VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_4 QN VDD mp15  l=0.13u w=0.69u m=1
M19 N_9 G VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_73 D N_14 VDD mp15  l=0.13u w=0.5u m=1
M21 N_13 N_9 N_14 VDD mp15  l=0.13u w=0.59u m=1
M22 VDD N_9 N_10 VDD mp15  l=0.13u w=0.42u m=1
M23 N_76 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 N_76 N_4 N_75 VDD mp15  l=0.13u w=0.17u m=1
M25 N_75 N_10 N_13 VDD mp15  l=0.13u w=0.17u m=1
M26 N_14 D N_74 VDD mp15  l=0.13u w=0.48u m=1
M27 N_74 N_17 VDD VDD mp15  l=0.13u w=0.48u m=1
M28 N_73 N_17 VDD VDD mp15  l=0.13u w=0.5u m=1
M29 N_17 SN VDD VDD mp15  l=0.13u w=0.42u m=1
.ends laphb2
* SPICE INPUT		Tue Jul 31 19:40:11 2018	laphb3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laphb3
.subckt laphb3 GND QN Q G VDD D SN
M1 N_3 SN GND GND mn15  l=0.13u w=0.37u m=1
M2 GND D N_7 GND mn15  l=0.13u w=0.3u m=1
M3 N_7 D GND GND mn15  l=0.13u w=0.29u m=1
M4 GND N_3 N_8 GND mn15  l=0.13u w=0.46u m=1
M5 N_7 N_4 N_8 GND mn15  l=0.13u w=0.325u m=1
M6 N_8 N_4 N_7 GND mn15  l=0.13u w=0.315u m=1
M7 N_22 N_19 GND GND mn15  l=0.13u w=0.17u m=1
M8 GND N_14 N_4 GND mn15  l=0.13u w=0.17u m=1
M9 N_22 N_14 N_8 GND mn15  l=0.13u w=0.17u m=1
M10 QN N_19 GND GND mn15  l=0.13u w=0.46u m=1
M11 QN N_19 GND GND mn15  l=0.13u w=0.46u m=1
M12 QN N_19 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND G N_14 GND mn15  l=0.13u w=0.17u m=1
M14 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M15 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M16 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M17 GND N_8 N_19 GND mn15  l=0.13u w=0.41u m=1
M18 N_3 SN VDD VDD mp15  l=0.13u w=0.55u m=1
M19 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_19 N_8 VDD VDD mp15  l=0.13u w=0.62u m=1
M23 N_82 D N_7 VDD mp15  l=0.13u w=0.62u m=1
M24 N_83 N_3 VDD VDD mp15  l=0.13u w=0.54u m=1
M25 N_82 N_3 VDD VDD mp15  l=0.13u w=0.62u m=1
M26 N_83 D N_7 VDD mp15  l=0.13u w=0.54u m=1
M27 N_84 N_4 N_8 VDD mp15  l=0.13u w=0.17u m=1
M28 N_85 N_19 N_84 VDD mp15  l=0.13u w=0.17u m=1
M29 N_85 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 VDD N_14 N_4 VDD mp15  l=0.13u w=0.42u m=1
M31 N_8 N_14 N_7 VDD mp15  l=0.13u w=0.56u m=1
M32 QN N_19 VDD VDD mp15  l=0.13u w=0.69u m=1
M33 QN N_19 VDD VDD mp15  l=0.13u w=0.69u m=1
M34 QN N_19 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 VDD G N_14 VDD mp15  l=0.13u w=0.42u m=1
.ends laphb3
* SPICE INPUT		Tue Jul 31 19:40:24 2018	laplb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb0
.subckt laplb0 VDD QN Q GND GN D SN
M1 GND SN N_3 GND mn15  l=0.13u w=0.18u m=1
M2 GND N_3 N_14 GND mn15  l=0.13u w=0.18u m=1
M3 N_14 N_6 N_13 GND mn15  l=0.13u w=0.28u m=1
M4 GND N_6 N_10 GND mn15  l=0.13u w=0.17u m=1
M5 N_62 N_10 N_14 GND mn15  l=0.13u w=0.17u m=1
M6 N_62 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M7 N_13 D GND GND mn15  l=0.13u w=0.19u m=1
M8 N_6 GN GND GND mn15  l=0.13u w=0.17u m=1
M9 QN N_9 GND GND mn15  l=0.13u w=0.26u m=1
M10 Q N_14 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_9 N_14 GND GND mn15  l=0.13u w=0.18u m=1
M12 N_3 SN VDD VDD mp15  l=0.13u w=0.26u m=1
M13 N_6 GN VDD VDD mp15  l=0.13u w=0.42u m=1
M14 VDD N_9 QN VDD mp15  l=0.13u w=0.4u m=1
M15 Q N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_9 N_14 VDD VDD mp15  l=0.13u w=0.26u m=1
M17 N_15 N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M18 N_17 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M19 VDD N_6 N_10 VDD mp15  l=0.13u w=0.42u m=1
M20 N_16 N_6 N_14 VDD mp15  l=0.13u w=0.17u m=1
M21 N_14 N_10 N_13 VDD mp15  l=0.13u w=0.42u m=1
M22 N_17 N_9 N_16 VDD mp15  l=0.13u w=0.17u m=1
M23 N_15 D N_13 VDD mp15  l=0.13u w=0.5u m=1
.ends laplb0
* SPICE INPUT		Tue Jul 31 19:40:37 2018	laplb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb1
.subckt laplb1 GND QN Q GN VDD D SN
M1 N_3 SN GND GND mn15  l=0.13u w=0.28u m=1
M2 GND N_11 N_4 GND mn15  l=0.13u w=0.17u m=1
M3 N_7 N_11 N_8 GND mn15  l=0.13u w=0.37u m=1
M4 N_7 N_3 GND GND mn15  l=0.13u w=0.28u m=1
M5 N_8 D GND GND mn15  l=0.13u w=0.33u m=1
M6 N_17 N_4 N_7 GND mn15  l=0.13u w=0.17u m=1
M7 N_17 N_16 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_11 GN GND GND mn15  l=0.13u w=0.17u m=1
M9 QN N_16 GND GND mn15  l=0.13u w=0.46u m=1
M10 Q N_7 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_16 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M12 N_3 SN VDD VDD mp15  l=0.13u w=0.42u m=1
M13 N_70 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M14 VDD N_11 N_4 VDD mp15  l=0.13u w=0.42u m=1
M15 N_69 N_11 N_7 VDD mp15  l=0.13u w=0.17u m=1
M16 N_67 D N_8 VDD mp15  l=0.13u w=0.46u m=1
M17 N_68 N_3 VDD VDD mp15  l=0.13u w=0.46u m=1
M18 N_67 N_3 VDD VDD mp15  l=0.13u w=0.46u m=1
M19 N_8 D N_68 VDD mp15  l=0.13u w=0.46u m=1
M20 N_7 N_4 N_8 VDD mp15  l=0.13u w=0.55u m=1
M21 N_70 N_16 N_69 VDD mp15  l=0.13u w=0.17u m=1
M22 N_11 GN VDD VDD mp15  l=0.13u w=0.42u m=1
M23 Q N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_16 N_7 VDD VDD mp15  l=0.13u w=0.39u m=1
M25 QN N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends laplb1
* SPICE INPUT		Tue Jul 31 19:40:49 2018	laplb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb2
.subckt laplb2 GND QN Q VDD GN D SN
M1 N_3 SN GND GND mn15  l=0.13u w=0.28u m=1
M2 N_7 N_3 GND GND mn15  l=0.13u w=0.36u m=1
M3 N_8 D GND GND mn15  l=0.13u w=0.4u m=1
M4 N_18 N_4 N_7 GND mn15  l=0.13u w=0.17u m=1
M5 N_18 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M6 GND N_11 N_4 GND mn15  l=0.13u w=0.17u m=1
M7 N_7 N_11 N_8 GND mn15  l=0.13u w=0.52u m=1
M8 N_11 GN GND GND mn15  l=0.13u w=0.17u m=1
M9 GND N_7 Q GND mn15  l=0.13u w=0.46u m=1
M10 Q N_7 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_7 N_14 GND mn15  l=0.13u w=0.37u m=1
M12 GND N_14 QN GND mn15  l=0.13u w=0.46u m=1
M13 GND N_14 QN GND mn15  l=0.13u w=0.46u m=1
M14 N_3 SN VDD VDD mp15  l=0.13u w=0.42u m=1
M15 N_73 D N_8 VDD mp15  l=0.13u w=0.535u m=1
M16 N_74 N_3 VDD VDD mp15  l=0.13u w=0.535u m=1
M17 N_73 N_3 VDD VDD mp15  l=0.13u w=0.535u m=1
M18 N_8 D N_74 VDD mp15  l=0.13u w=0.535u m=1
M19 N_7 N_4 N_8 VDD mp15  l=0.13u w=0.59u m=1
M20 N_76 N_14 N_75 VDD mp15  l=0.13u w=0.16u m=1
M21 N_76 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 VDD N_11 N_4 VDD mp15  l=0.13u w=0.42u m=1
M23 N_75 N_11 N_7 VDD mp15  l=0.13u w=0.16u m=1
M24 N_11 GN VDD VDD mp15  l=0.13u w=0.42u m=1
M25 Q N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 Q N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_14 N_7 VDD VDD mp15  l=0.13u w=0.55u m=1
M28 VDD N_14 QN VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_14 QN VDD mp15  l=0.13u w=0.69u m=1
.ends laplb2
* SPICE INPUT		Tue Jul 31 19:41:02 2018	laplb3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=laplb3
.subckt laplb3 GND Q QN SN D VDD GN
M1 Q N_16 GND GND mn15  l=0.13u w=0.46u m=1
M2 Q N_16 GND GND mn15  l=0.13u w=0.46u m=1
M3 Q N_16 GND GND mn15  l=0.13u w=0.46u m=1
M4 GND N_16 N_4 GND mn15  l=0.13u w=0.45u m=1
M5 QN N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 QN N_4 GND GND mn15  l=0.13u w=0.46u m=1
M7 QN N_4 GND GND mn15  l=0.13u w=0.46u m=1
M8 GND GN N_9 GND mn15  l=0.13u w=0.17u m=1
M9 N_14 N_9 N_16 GND mn15  l=0.13u w=0.32u m=1
M10 GND N_9 N_12 GND mn15  l=0.13u w=0.17u m=1
M11 N_16 N_9 N_14 GND mn15  l=0.13u w=0.31u m=1
M12 N_22 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M13 N_22 N_12 N_16 GND mn15  l=0.13u w=0.17u m=1
M14 GND N_21 N_16 GND mn15  l=0.13u w=0.46u m=1
M15 GND D N_14 GND mn15  l=0.13u w=0.3u m=1
M16 GND D N_14 GND mn15  l=0.13u w=0.33u m=1
M17 N_21 SN GND GND mn15  l=0.13u w=0.33u m=1
M18 Q N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 Q N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Q N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_4 N_16 VDD VDD mp15  l=0.13u w=0.67u m=1
M22 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 VDD GN N_9 VDD mp15  l=0.13u w=0.42u m=1
M26 VDD N_9 N_12 VDD mp15  l=0.13u w=0.42u m=1
M27 N_84 N_9 N_16 VDD mp15  l=0.13u w=0.17u m=1
M28 N_85 N_21 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_85 N_4 N_84 VDD mp15  l=0.13u w=0.17u m=1
M30 N_16 N_12 N_14 VDD mp15  l=0.13u w=0.59u m=1
M31 N_83 D N_14 VDD mp15  l=0.13u w=0.6u m=1
M32 N_83 N_21 VDD VDD mp15  l=0.13u w=0.6u m=1
M33 N_82 N_21 VDD VDD mp15  l=0.13u w=0.7u m=1
M34 N_82 D N_14 VDD mp15  l=0.13u w=0.7u m=1
M35 N_21 SN VDD VDD mp15  l=0.13u w=0.5u m=1
.ends laplb3
* SPICE INPUT		Tue Jul 31 19:41:16 2018	mi02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d0
.subckt mi02d0 GND Y S0 VDD B A
M1 GND B N_2 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 N_6 GND mn15  l=0.13u w=0.26u m=1
M3 Y S0 N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 A GND GND mn15  l=0.13u w=0.26u m=1
M5 GND S0 N_4 GND mn15  l=0.13u w=0.26u m=1
M6 VDD B N_2 VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 N_2 VDD mp15  l=0.13u w=0.4u m=1
M8 Y S0 N_6 VDD mp15  l=0.13u w=0.4u m=1
M9 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_4 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mi02d0
* SPICE INPUT		Tue Jul 31 19:41:29 2018	mi02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d1
.subckt mi02d1 GND Y S0 A B VDD
M1 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M2 Y S0 N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M4 Y N_4 N_6 GND mn15  l=0.13u w=0.46u m=1
M5 GND S0 N_4 GND mn15  l=0.13u w=0.28u m=1
M6 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M7 Y S0 N_6 VDD mp15  l=0.13u w=0.59u m=1
M8 N_6 A VDD VDD mp15  l=0.13u w=0.59u m=1
M9 Y N_4 N_2 VDD mp15  l=0.13u w=0.69u m=1
M10 N_4 S0 VDD VDD mp15  l=0.13u w=0.39u m=1
.ends mi02d1
* SPICE INPUT		Tue Jul 31 19:41:43 2018	mi02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d2
.subckt mi02d2 GND Y S0 B A VDD
M1 GND S0 N_4 GND mn15  l=0.13u w=0.37u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_7 N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_7 N_4 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y S0 N_2 GND mn15  l=0.13u w=0.46u m=1
M9 N_2 S0 Y GND mn15  l=0.13u w=0.46u m=1
M10 N_4 S0 VDD VDD mp15  l=0.13u w=0.55u m=1
M11 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD B N_2 VDD mp15  l=0.13u w=0.69u m=1
M13 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_7 S0 Y VDD mp15  l=0.13u w=0.595u m=1
M16 N_7 S0 Y VDD mp15  l=0.13u w=0.595u m=1
M17 N_2 N_4 Y VDD mp15  l=0.13u w=0.565u m=1
M18 N_2 N_4 Y VDD mp15  l=0.13u w=0.565u m=1
.ends mi02d2
* SPICE INPUT		Tue Jul 31 19:41:56 2018	mi02d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02d3
.subckt mi02d3 Y GND S0 A B VDD
M1 N_3 S0 Y GND mn15  l=0.13u w=0.46u m=1
M2 N_3 S0 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_3 S0 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_14 N_6 GND mn15  l=0.13u w=0.46u m=1
M5 N_6 N_14 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_6 N_14 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M10 GND S0 N_14 GND mn15  l=0.13u w=0.45u m=1
M11 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M12 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M13 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M14 N_14 S0 VDD VDD mp15  l=0.13u w=0.67u m=1
M15 N_3 B VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_3 B VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_3 B VDD VDD mp15  l=0.13u w=0.69u m=1
M18 Y S0 N_6 VDD mp15  l=0.13u w=0.59u m=1
M19 Y S0 N_6 VDD mp15  l=0.13u w=0.57u m=1
M20 N_6 S0 Y VDD mp15  l=0.13u w=0.57u m=1
M21 Y N_14 N_3 VDD mp15  l=0.13u w=0.61u m=1
M22 N_3 N_14 Y VDD mp15  l=0.13u w=0.575u m=1
M23 N_3 N_14 Y VDD mp15  l=0.13u w=0.575u m=1
M24 N_6 A VDD VDD mp15  l=0.13u w=0.65u m=1
M25 VDD A N_6 VDD mp15  l=0.13u w=0.65u m=1
M26 VDD A N_6 VDD mp15  l=0.13u w=0.66u m=1
.ends mi02d3
* SPICE INPUT		Tue Jul 31 19:42:10 2018	mi02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mi02dm
.subckt mi02dm GND Y VDD B A S0
M1 GND S0 N_4 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.36u m=1
M3 Y S0 N_2 GND mn15  l=0.13u w=0.36u m=1
M4 Y N_4 N_6 GND mn15  l=0.13u w=0.36u m=1
M5 N_6 A GND GND mn15  l=0.13u w=0.36u m=1
M6 N_4 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M7 VDD B N_2 VDD mp15  l=0.13u w=0.55u m=1
M8 Y N_4 N_2 VDD mp15  l=0.13u w=0.55u m=1
M9 Y S0 N_6 VDD mp15  l=0.13u w=0.55u m=1
M10 N_6 A VDD VDD mp15  l=0.13u w=0.55u m=1
.ends mi02dm
* SPICE INPUT		Tue Jul 31 19:42:23 2018	mx02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d0
.subckt mx02d0 VDD Y B A GND S0
M1 N_16 B GND GND mn15  l=0.13u w=0.18u m=1
M2 N_15 A GND GND mn15  l=0.13u w=0.18u m=1
M3 N_15 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M4 N_16 S0 N_6 GND mn15  l=0.13u w=0.18u m=1
M5 GND S0 N_5 GND mn15  l=0.13u w=0.18u m=1
M6 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_10 B VDD VDD mp15  l=0.13u w=0.26u m=1
M8 N_9 A VDD VDD mp15  l=0.13u w=0.26u m=1
M9 N_10 N_5 N_6 VDD mp15  l=0.13u w=0.26u m=1
M10 N_5 S0 VDD VDD mp15  l=0.13u w=0.26u m=1
M11 N_6 S0 N_9 VDD mp15  l=0.13u w=0.26u m=1
M12 Y N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mx02d0
* SPICE INPUT		Tue Jul 31 19:42:36 2018	mx02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d1
.subckt mx02d1 VDD Y GND B A S0
M1 GND S0 N_4 GND mn15  l=0.13u w=0.18u m=1
M2 N_16 S0 N_6 GND mn15  l=0.13u w=0.22u m=1
M3 N_15 A GND GND mn15  l=0.13u w=0.22u m=1
M4 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_16 B GND GND mn15  l=0.13u w=0.22u m=1
M6 N_15 N_4 N_6 GND mn15  l=0.13u w=0.22u m=1
M7 N_6 S0 N_7 VDD mp15  l=0.13u w=0.37u m=1
M8 VDD S0 N_4 VDD mp15  l=0.13u w=0.24u m=1
M9 N_7 A VDD VDD mp15  l=0.13u w=0.37u m=1
M10 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 B VDD VDD mp15  l=0.13u w=0.37u m=1
M12 N_8 N_4 N_6 VDD mp15  l=0.13u w=0.37u m=1
.ends mx02d1
* SPICE INPUT		Tue Jul 31 19:42:49 2018	mx02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d2
.subckt mx02d2 Y GND VDD B A S0
M1 N_8 N_4 N_6 GND mn15  l=0.13u w=0.32u m=1
M2 GND B N_7 GND mn15  l=0.13u w=0.3u m=1
M3 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M4 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M5 N_6 A GND GND mn15  l=0.13u w=0.3u m=1
M6 GND S0 N_4 GND mn15  l=0.13u w=0.32u m=1
M7 N_8 S0 N_7 GND mn15  l=0.13u w=0.32u m=1
M8 N_8 N_4 N_7 VDD mp15  l=0.13u w=0.5u m=1
M9 VDD B N_7 VDD mp15  l=0.13u w=0.48u m=1
M10 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M12 N_6 A VDD VDD mp15  l=0.13u w=0.48u m=1
M13 N_4 S0 VDD VDD mp15  l=0.13u w=0.46u m=1
M14 N_8 S0 N_6 VDD mp15  l=0.13u w=0.5u m=1
.ends mx02d2
* SPICE INPUT		Tue Jul 31 19:43:02 2018	mx02d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02d3
.subckt mx02d3 VDD Y GND B A S0
M1 N_16 S0 GND GND mn15  l=0.13u w=0.27u m=1
M2 N_12 A GND GND mn15  l=0.13u w=0.23u m=1
M3 GND A N_12 GND mn15  l=0.13u w=0.22u m=1
M4 N_6 S0 N_9 GND mn15  l=0.13u w=0.23u m=1
M5 N_6 S0 N_9 GND mn15  l=0.13u w=0.22u m=1
M6 N_9 N_16 N_12 GND mn15  l=0.13u w=0.23u m=1
M7 N_12 N_16 N_9 GND mn15  l=0.13u w=0.22u m=1
M8 Y N_9 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_9 GND GND mn15  l=0.13u w=0.46u m=1
M10 Y N_9 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND B N_6 GND mn15  l=0.13u w=0.23u m=1
M12 N_6 B GND GND mn15  l=0.13u w=0.22u m=1
M13 Y N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M14 Y N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M15 Y N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_6 B VDD VDD mp15  l=0.13u w=0.335u m=1
M17 N_6 B VDD VDD mp15  l=0.13u w=0.335u m=1
M18 N_12 S0 N_9 VDD mp15  l=0.13u w=0.335u m=1
M19 N_12 S0 N_9 VDD mp15  l=0.13u w=0.335u m=1
M20 N_9 N_16 N_6 VDD mp15  l=0.13u w=0.32u m=1
M21 N_9 N_16 N_6 VDD mp15  l=0.13u w=0.32u m=1
M22 N_16 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M23 N_12 A VDD VDD mp15  l=0.13u w=0.32u m=1
M24 VDD A N_12 VDD mp15  l=0.13u w=0.32u m=1
.ends mx02d3
* SPICE INPUT		Tue Jul 31 19:43:14 2018	mx02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx02dm
.subckt mx02dm GND Y VDD B A S0
M1 N_7 A GND GND mn15  l=0.13u w=0.27u m=1
M2 Y N_6 GND GND mn15  l=0.13u w=0.36u m=1
M3 N_8 B GND GND mn15  l=0.13u w=0.27u m=1
M4 N_6 N_5 N_7 GND mn15  l=0.13u w=0.27u m=1
M5 N_8 S0 N_6 GND mn15  l=0.13u w=0.27u m=1
M6 N_5 S0 GND GND mn15  l=0.13u w=0.27u m=1
M7 N_15 A VDD VDD mp15  l=0.13u w=0.41u m=1
M8 Y N_6 VDD VDD mp15  l=0.13u w=0.55u m=1
M9 N_16 B VDD VDD mp15  l=0.13u w=0.41u m=1
M10 N_5 S0 VDD VDD mp15  l=0.13u w=0.41u m=1
M11 N_6 S0 N_15 VDD mp15  l=0.13u w=0.41u m=1
M12 N_16 N_5 N_6 VDD mp15  l=0.13u w=0.41u m=1
.ends mx02dm
* SPICE INPUT		Tue Jul 31 19:43:27 2018	mx03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx03d0
.subckt mx03d0 VDD Y C S1 A GND B S0
M1 N_6 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_8 S0 N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 S0 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_8 N_5 N_7 GND mn15  l=0.13u w=0.26u m=1
M5 GND S1 N_3 GND mn15  l=0.13u w=0.26u m=1
M6 N_7 A GND GND mn15  l=0.13u w=0.26u m=1
M7 Y N_12 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_12 N_3 N_8 GND mn15  l=0.13u w=0.26u m=1
M9 N_12 S1 N_13 GND mn15  l=0.13u w=0.26u m=1
M10 N_13 C GND GND mn15  l=0.13u w=0.26u m=1
M11 N_6 B VDD VDD mp15  l=0.13u w=0.4u m=1
M12 N_8 N_5 N_6 VDD mp15  l=0.13u w=0.26u m=1
M13 N_5 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_8 S0 N_7 VDD mp15  l=0.13u w=0.26u m=1
M15 N_3 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M17 Y N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_13 N_3 N_12 VDD mp15  l=0.13u w=0.26u m=1
M19 N_12 S1 N_8 VDD mp15  l=0.13u w=0.26u m=1
M20 N_13 C VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mx03d0
* SPICE INPUT		Tue Jul 31 19:43:41 2018	mx03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx03d1
.subckt mx03d1 VDD Y GND C S1 A B S0
M1 N_12 N_3 N_7 GND mn15  l=0.13u w=0.28u m=1
M2 N_12 S1 N_13 GND mn15  l=0.13u w=0.28u m=1
M3 N_13 C GND GND mn15  l=0.13u w=0.28u m=1
M4 Y N_12 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 B GND GND mn15  l=0.13u w=0.33u m=1
M6 N_5 S0 GND GND mn15  l=0.13u w=0.28u m=1
M7 N_7 S0 N_6 GND mn15  l=0.13u w=0.28u m=1
M8 N_8 N_5 N_7 GND mn15  l=0.13u w=0.28u m=1
M9 N_8 A GND GND mn15  l=0.13u w=0.33u m=1
M10 GND S1 N_3 GND mn15  l=0.13u w=0.28u m=1
M11 N_6 B VDD VDD mp15  l=0.13u w=0.5u m=1
M12 N_7 N_5 N_6 VDD mp15  l=0.13u w=0.28u m=1
M13 N_8 S0 N_7 VDD mp15  l=0.13u w=0.28u m=1
M14 N_5 S0 VDD VDD mp15  l=0.13u w=0.39u m=1
M15 N_8 A VDD VDD mp15  l=0.13u w=0.5u m=1
M16 N_3 S1 VDD VDD mp15  l=0.13u w=0.39u m=1
M17 N_13 N_3 N_12 VDD mp15  l=0.13u w=0.28u m=1
M18 N_12 S1 N_7 VDD mp15  l=0.13u w=0.28u m=1
M19 N_13 C VDD VDD mp15  l=0.13u w=0.42u m=1
M20 Y N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends mx03d1
* SPICE INPUT		Tue Jul 31 19:43:54 2018	mx03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx03d2
.subckt mx03d2 VDD Y A S1 GND C B S0
M1 N_3 B GND GND mn15  l=0.13u w=0.23u m=1
M2 GND B N_3 GND mn15  l=0.13u w=0.23u m=1
M3 N_5 S0 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_8 S0 N_3 GND mn15  l=0.13u w=0.37u m=1
M5 N_8 N_5 N_10 GND mn15  l=0.13u w=0.37u m=1
M6 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M7 GND S1 N_7 GND mn15  l=0.13u w=0.28u m=1
M8 GND N_14 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_14 Y GND mn15  l=0.13u w=0.46u m=1
M10 N_8 N_7 N_14 GND mn15  l=0.13u w=0.37u m=1
M11 N_15 S1 N_14 GND mn15  l=0.13u w=0.37u m=1
M12 GND C N_15 GND mn15  l=0.13u w=0.41u m=1
M13 VDD B N_3 VDD mp15  l=0.13u w=0.39u m=1
M14 N_3 B VDD VDD mp15  l=0.13u w=0.3u m=1
M15 N_5 S0 VDD VDD mp15  l=0.13u w=0.39u m=1
M16 N_3 N_5 N_8 VDD mp15  l=0.13u w=0.37u m=1
M17 N_10 S0 N_8 VDD mp15  l=0.13u w=0.37u m=1
M18 N_10 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_7 S1 VDD VDD mp15  l=0.13u w=0.39u m=1
M20 VDD N_14 Y VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_14 Y VDD mp15  l=0.13u w=0.69u m=1
M22 N_15 N_7 N_14 VDD mp15  l=0.13u w=0.37u m=1
M23 N_14 S1 N_8 VDD mp15  l=0.13u w=0.37u m=1
M24 VDD C N_15 VDD mp15  l=0.13u w=0.61u m=1
.ends mx03d2
* SPICE INPUT		Tue Jul 31 19:44:07 2018	mx03d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx03d3
.subckt mx03d3 GND Y S1 VDD C B A S0
M1 N_3 B GND GND mn15  l=0.13u w=0.23u m=1
M2 GND B N_3 GND mn15  l=0.13u w=0.23u m=1
M3 N_5 S0 GND GND mn15  l=0.13u w=0.28u m=1
M4 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M6 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_9 N_13 N_8 GND mn15  l=0.13u w=0.37u m=1
M8 GND C N_10 GND mn15  l=0.13u w=0.46u m=1
M9 N_10 S1 N_8 GND mn15  l=0.13u w=0.37u m=1
M10 N_9 S0 N_3 GND mn15  l=0.13u w=0.37u m=1
M11 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M12 N_9 N_5 N_16 GND mn15  l=0.13u w=0.37u m=1
M13 GND S1 N_13 GND mn15  l=0.13u w=0.28u m=1
M14 N_3 N_5 N_9 VDD mp15  l=0.13u w=0.37u m=1
M15 N_16 S0 N_9 VDD mp15  l=0.13u w=0.37u m=1
M16 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_13 S1 VDD VDD mp15  l=0.13u w=0.39u m=1
M18 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_10 N_13 N_8 VDD mp15  l=0.13u w=0.37u m=1
M22 N_10 C VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_8 S1 N_9 VDD mp15  l=0.13u w=0.37u m=1
M24 N_3 B VDD VDD mp15  l=0.13u w=0.3u m=1
M25 VDD B N_3 VDD mp15  l=0.13u w=0.39u m=1
M26 N_5 S0 VDD VDD mp15  l=0.13u w=0.39u m=1
.ends mx03d3
* SPICE INPUT		Tue Jul 31 19:44:19 2018	mx04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d0
.subckt mx04d0 VDD Y S1 B A D S0 GND C
M1 N_68 C GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 N_4 N_68 GND mn15  l=0.13u w=0.26u m=1
M3 N_69 D GND GND mn15  l=0.13u w=0.26u m=1
M4 N_70 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_2 N_4 N_67 GND mn15  l=0.13u w=0.26u m=1
M6 N_70 S0 N_2 GND mn15  l=0.13u w=0.26u m=1
M7 N_69 S0 N_5 GND mn15  l=0.13u w=0.26u m=1
M8 N_4 S0 GND GND mn15  l=0.13u w=0.26u m=1
M9 N_67 A GND GND mn15  l=0.13u w=0.26u m=1
M10 Y N_7 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_13 S1 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_2 N_13 N_7 GND mn15  l=0.13u w=0.26u m=1
M13 N_5 S1 N_7 GND mn15  l=0.13u w=0.26u m=1
M14 N_15 C VDD VDD mp15  l=0.13u w=0.4u m=1
M15 N_15 S0 N_5 VDD mp15  l=0.13u w=0.4u m=1
M16 N_16 N_4 N_5 VDD mp15  l=0.13u w=0.4u m=1
M17 VDD D N_16 VDD mp15  l=0.13u w=0.4u m=1
M18 VDD B N_14 VDD mp15  l=0.13u w=0.4u m=1
M19 N_2 N_4 N_14 VDD mp15  l=0.13u w=0.4u m=1
M20 N_4 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_5 N_13 N_7 VDD mp15  l=0.13u w=0.26u m=1
M22 N_2 S1 N_7 VDD mp15  l=0.13u w=0.26u m=1
M23 N_17 S0 N_2 VDD mp15  l=0.13u w=0.4u m=1
M24 N_17 A VDD VDD mp15  l=0.13u w=0.4u m=1
M25 Y N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M26 N_13 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mx04d0
* SPICE INPUT		Tue Jul 31 19:44:32 2018	mx04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d1
.subckt mx04d1 VDD Y A B S1 D S0 C GND
M1 N_69 C GND GND mn15  l=0.13u w=0.32u m=1
M2 N_69 N_4 N_5 GND mn15  l=0.13u w=0.32u m=1
M3 GND D N_70 GND mn15  l=0.13u w=0.32u m=1
M4 N_71 B GND GND mn15  l=0.13u w=0.32u m=1
M5 N_2 N_4 N_68 GND mn15  l=0.13u w=0.32u m=1
M6 N_68 A GND GND mn15  l=0.13u w=0.32u m=1
M7 N_4 S0 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_2 S0 N_71 GND mn15  l=0.13u w=0.32u m=1
M9 N_70 S0 N_5 GND mn15  l=0.13u w=0.32u m=1
M10 N_2 N_14 N_9 GND mn15  l=0.13u w=0.28u m=1
M11 N_5 S1 N_9 GND mn15  l=0.13u w=0.28u m=1
M12 Y N_9 GND GND mn15  l=0.13u w=0.46u m=1
M13 N_14 S1 GND GND mn15  l=0.13u w=0.26u m=1
M14 N_16 C VDD VDD mp15  l=0.13u w=0.47u m=1
M15 N_16 S0 N_5 VDD mp15  l=0.13u w=0.47u m=1
M16 N_17 N_4 N_5 VDD mp15  l=0.13u w=0.47u m=1
M17 N_17 D VDD VDD mp15  l=0.13u w=0.47u m=1
M18 VDD B N_15 VDD mp15  l=0.13u w=0.47u m=1
M19 N_2 N_4 N_15 VDD mp15  l=0.13u w=0.47u m=1
M20 N_4 S0 VDD VDD mp15  l=0.13u w=0.42u m=1
M21 VDD A N_18 VDD mp15  l=0.13u w=0.47u m=1
M22 N_2 S0 N_18 VDD mp15  l=0.13u w=0.47u m=1
M23 N_5 N_14 N_9 VDD mp15  l=0.13u w=0.28u m=1
M24 N_2 S1 N_9 VDD mp15  l=0.13u w=0.28u m=1
M25 Y N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_14 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends mx04d1
* SPICE INPUT		Tue Jul 31 19:44:45 2018	mx04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d2
.subckt mx04d2 GND Y VDD S1 A S0 B D C
M1 N_3 S0 GND GND mn15  l=0.13u w=0.37u m=1
M2 N_21 N_3 N_4 GND mn15  l=0.13u w=0.225u m=1
M3 N_22 C GND GND mn15  l=0.13u w=0.225u m=1
M4 N_21 C GND GND mn15  l=0.13u w=0.225u m=1
M5 GND D N_20 GND mn15  l=0.13u w=0.225u m=1
M6 N_23 D GND GND mn15  l=0.13u w=0.225u m=1
M7 N_20 S0 N_4 GND mn15  l=0.13u w=0.225u m=1
M8 N_23 S0 N_4 GND mn15  l=0.13u w=0.225u m=1
M9 N_22 N_3 N_4 GND mn15  l=0.13u w=0.225u m=1
M10 N_10 S0 N_24 GND mn15  l=0.13u w=0.45u m=1
M11 N_24 B GND GND mn15  l=0.13u w=0.45u m=1
M12 N_10 N_3 N_25 GND mn15  l=0.13u w=0.45u m=1
M13 N_25 A GND GND mn15  l=0.13u w=0.45u m=1
M14 N_10 N_18 N_13 GND mn15  l=0.13u w=0.32u m=1
M15 N_4 S1 N_13 GND mn15  l=0.13u w=0.36u m=1
M16 GND S1 N_18 GND mn15  l=0.13u w=0.26u m=1
M17 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M18 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M19 N_3 S0 VDD VDD mp15  l=0.13u w=0.55u m=1
M20 N_107 C VDD VDD mp15  l=0.13u w=0.32u m=1
M21 N_106 C VDD VDD mp15  l=0.13u w=0.33u m=1
M22 N_108 D VDD VDD mp15  l=0.13u w=0.29u m=1
M23 VDD D N_105 VDD mp15  l=0.13u w=0.36u m=1
M24 N_106 S0 N_4 VDD mp15  l=0.13u w=0.33u m=1
M25 N_107 S0 N_4 VDD mp15  l=0.13u w=0.32u m=1
M26 N_108 N_3 N_4 VDD mp15  l=0.13u w=0.29u m=1
M27 N_4 N_3 N_105 VDD mp15  l=0.13u w=0.36u m=1
M28 N_110 B VDD VDD mp15  l=0.13u w=0.31u m=1
M29 VDD B N_109 VDD mp15  l=0.13u w=0.34u m=1
M30 N_10 N_3 N_110 VDD mp15  l=0.13u w=0.31u m=1
M31 N_10 N_3 N_109 VDD mp15  l=0.13u w=0.34u m=1
M32 N_111 A VDD VDD mp15  l=0.13u w=0.31u m=1
M33 N_112 A VDD VDD mp15  l=0.13u w=0.3u m=1
M34 N_111 S0 N_10 VDD mp15  l=0.13u w=0.31u m=1
M35 N_10 S0 N_112 VDD mp15  l=0.13u w=0.3u m=1
M36 N_13 N_18 N_4 VDD mp15  l=0.13u w=0.35u m=1
M37 N_10 S1 N_13 VDD mp15  l=0.13u w=0.35u m=1
M38 N_18 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
M39 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
M40 VDD N_13 Y VDD mp15  l=0.13u w=0.69u m=1
.ends mx04d2
* SPICE INPUT		Tue Jul 31 19:44:58 2018	mx04d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04d3
.subckt mx04d3 GND Y S0 S1 B D A VDD C
M1 N_3 S0 GND GND mn15  l=0.13u w=0.36u m=1
M2 N_21 S0 N_4 GND mn15  l=0.13u w=0.225u m=1
M3 N_24 S0 N_4 GND mn15  l=0.13u w=0.225u m=1
M4 N_22 N_3 N_4 GND mn15  l=0.13u w=0.225u m=1
M5 N_23 N_3 N_4 GND mn15  l=0.13u w=0.225u m=1
M6 N_23 C GND GND mn15  l=0.13u w=0.225u m=1
M7 N_22 C GND GND mn15  l=0.13u w=0.225u m=1
M8 GND D N_21 GND mn15  l=0.13u w=0.225u m=1
M9 N_24 D GND GND mn15  l=0.13u w=0.225u m=1
M10 N_10 S0 N_25 GND mn15  l=0.13u w=0.45u m=1
M11 N_25 B GND GND mn15  l=0.13u w=0.45u m=1
M12 N_10 N_3 N_26 GND mn15  l=0.13u w=0.45u m=1
M13 N_26 A GND GND mn15  l=0.13u w=0.45u m=1
M14 N_4 S1 N_13 GND mn15  l=0.13u w=0.45u m=1
M15 N_10 N_18 N_13 GND mn15  l=0.13u w=0.32u m=1
M16 GND S1 N_18 GND mn15  l=0.13u w=0.28u m=1
M17 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M18 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M19 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M20 N_3 S0 VDD VDD mp15  l=0.13u w=0.53u m=1
M21 N_50 S0 N_4 VDD mp15  l=0.13u w=0.33u m=1
M22 N_51 S0 N_4 VDD mp15  l=0.13u w=0.32u m=1
M23 N_52 N_3 N_4 VDD mp15  l=0.13u w=0.29u m=1
M24 N_4 N_3 N_49 VDD mp15  l=0.13u w=0.36u m=1
M25 N_51 C VDD VDD mp15  l=0.13u w=0.32u m=1
M26 N_50 C VDD VDD mp15  l=0.13u w=0.33u m=1
M27 VDD D N_49 VDD mp15  l=0.13u w=0.36u m=1
M28 N_52 D VDD VDD mp15  l=0.13u w=0.29u m=1
M29 N_54 N_3 N_10 VDD mp15  l=0.13u w=0.32u m=1
M30 N_10 N_3 N_53 VDD mp15  l=0.13u w=0.33u m=1
M31 N_54 B VDD VDD mp15  l=0.13u w=0.32u m=1
M32 VDD B N_53 VDD mp15  l=0.13u w=0.33u m=1
M33 N_56 A VDD VDD mp15  l=0.13u w=0.31u m=1
M34 N_55 A VDD VDD mp15  l=0.13u w=0.31u m=1
M35 N_10 S1 N_13 VDD mp15  l=0.13u w=0.53u m=1
M36 N_4 N_18 N_13 VDD mp15  l=0.13u w=0.53u m=1
M37 N_55 S0 N_10 VDD mp15  l=0.13u w=0.31u m=1
M38 N_10 S0 N_56 VDD mp15  l=0.13u w=0.31u m=1
M39 N_18 S1 VDD VDD mp15  l=0.13u w=0.42u m=1
M40 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M42 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends mx04d3
* SPICE INPUT		Tue Jul 31 19:45:11 2018	mx04dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=mx04dm
.subckt mx04dm VDD Y GND A D B S1 S0 C
M1 Y N_5 GND GND mn15  l=0.13u w=0.36u m=1
M2 N_4 S1 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_69 D GND GND mn15  l=0.13u w=0.26u m=1
M4 N_70 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 N_11 N_67 GND mn15  l=0.13u w=0.26u m=1
M6 N_11 S0 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_70 S0 N_8 GND mn15  l=0.13u w=0.26u m=1
M8 N_69 S0 N_6 GND mn15  l=0.13u w=0.26u m=1
M9 N_67 A GND GND mn15  l=0.13u w=0.26u m=1
M10 N_68 C GND GND mn15  l=0.13u w=0.26u m=1
M11 N_6 N_11 N_68 GND mn15  l=0.13u w=0.26u m=1
M12 N_8 N_4 N_5 GND mn15  l=0.13u w=0.26u m=1
M13 N_6 S1 N_5 GND mn15  l=0.13u w=0.26u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.55u m=1
M15 N_4 S1 VDD VDD mp15  l=0.13u w=0.4u m=1
M16 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.26u m=1
M17 N_14 S0 N_8 VDD mp15  l=0.13u w=0.4u m=1
M18 N_8 S1 N_5 VDD mp15  l=0.13u w=0.26u m=1
M19 N_14 A VDD VDD mp15  l=0.13u w=0.4u m=1
M20 VDD D N_17 VDD mp15  l=0.13u w=0.4u m=1
M21 N_16 S0 N_6 VDD mp15  l=0.13u w=0.4u m=1
M22 VDD B N_15 VDD mp15  l=0.13u w=0.4u m=1
M23 N_8 N_11 N_15 VDD mp15  l=0.13u w=0.4u m=1
M24 N_11 S0 VDD VDD mp15  l=0.13u w=0.4u m=1
M25 N_16 C VDD VDD mp15  l=0.13u w=0.4u m=1
M26 N_17 N_11 N_6 VDD mp15  l=0.13u w=0.4u m=1
.ends mx04dm
* SPICE INPUT		Tue Jul 31 19:45:23 2018	nd02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d0
.subckt nd02d0 VDD Y GND B A
M1 GND A N_14 GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.26u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.35u m=1
M4 Y B VDD VDD mp15  l=0.13u w=0.35u m=1
.ends nd02d0
* SPICE INPUT		Tue Jul 31 19:45:36 2018	nd02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d1
.subckt nd02d1 Y VDD A B GND
M1 GND A N_14 GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.46u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
.ends nd02d1
* SPICE INPUT		Tue Jul 31 19:45:49 2018	nd02d1p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d1p5
.subckt nd02d1p5 Y VDD A B GND
M1 GND A N_14 GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.46u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
.ends nd02d1p5
* SPICE INPUT		Tue Jul 31 19:46:02 2018	nd02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d2
.subckt nd02d2 GND Y VDD A B
M1 Y B N_5 GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M5 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M6 Y B VDD VDD mp15  l=0.13u w=0.61u m=1
M7 Y A VDD VDD mp15  l=0.13u w=0.61u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.61u m=1
.ends nd02d2
* SPICE INPUT		Tue Jul 31 19:46:15 2018	nd02d2p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d2p5
.subckt nd02d2p5 GND Y A B VDD
M1 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y B N_5 GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M5 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nd02d2p5
* SPICE INPUT		Tue Jul 31 19:46:28 2018	nd02d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d3
.subckt nd02d3 Y GND A VDD B
M1 N_3 B Y GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B Y GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B Y GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B Y GND mn15  l=0.13u w=0.46u m=1
M5 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M8 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M9 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M10 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M11 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M12 Y B VDD VDD mp15  l=0.13u w=0.61u m=1
M13 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
M14 Y A VDD VDD mp15  l=0.13u w=0.61u m=1
M15 VDD A Y VDD mp15  l=0.13u w=0.61u m=1
M16 Y A VDD VDD mp15  l=0.13u w=0.61u m=1
.ends nd02d3
* SPICE INPUT		Tue Jul 31 19:46:41 2018	nd02d3p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02d3p5
.subckt nd02d3p5 GND Y VDD A B
M1 N_8 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_9 B Y GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_8 GND mn15  l=0.13u w=0.46u m=1
M4 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_7 GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M8 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M11 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD B Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y B VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nd02d3p5
* SPICE INPUT		Tue Jul 31 19:46:54 2018	nd02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02dm
.subckt nd02dm Y VDD GND A B
M1 GND A N_14 GND mn15  l=0.13u w=0.36u m=1
M2 Y B N_14 GND mn15  l=0.13u w=0.36u m=1
M3 VDD A Y VDD mp15  l=0.13u w=0.45u m=1
M4 VDD B Y VDD mp15  l=0.13u w=0.45u m=1
.ends nd02dm
* SPICE INPUT		Tue Jul 31 19:47:07 2018	nd02od
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd02od
.subckt nd02od VDD B GND A Y
M1 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_22 B N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_3 N_5 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_22 A GND GND mn15  l=0.13u w=0.26u m=1
M5 N_5 B VDD VDD mp15  l=0.13u w=0.35u m=1
M6 N_3 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_5 A VDD VDD mp15  l=0.13u w=0.35u m=1
.ends nd02od
* SPICE INPUT		Tue Jul 31 19:47:20 2018	nd03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d0
.subckt nd03d0 VDD Y C B A GND
M1 N_19 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_19 B N_18 GND mn15  l=0.13u w=0.26u m=1
M3 Y C N_18 GND mn15  l=0.13u w=0.26u m=1
M4 Y A VDD VDD mp15  l=0.13u w=0.31u m=1
M5 Y B VDD VDD mp15  l=0.13u w=0.31u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.31u m=1
.ends nd03d0
* SPICE INPUT		Tue Jul 31 19:47:34 2018	nd03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d1
.subckt nd03d1 VDD Y C B A GND
M1 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M2 Y C N_18 GND mn15  l=0.13u w=0.46u m=1
M3 N_19 B N_18 GND mn15  l=0.13u w=0.46u m=1
M4 Y A VDD VDD mp15  l=0.13u w=0.54u m=1
M5 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M6 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
.ends nd03d1
* SPICE INPUT		Tue Jul 31 19:47:46 2018	nd03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d2
.subckt nd03d2 GND Y B C A VDD
M1 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_8 B N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_8 C Y GND mn15  l=0.13u w=0.46u m=1
M5 Y C N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M8 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
M9 VDD B Y VDD mp15  l=0.13u w=0.54u m=1
M10 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M11 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M12 Y A VDD VDD mp15  l=0.13u w=0.54u m=1
.ends nd03d2
* SPICE INPUT		Tue Jul 31 19:47:59 2018	nd03d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03d3
.subckt nd03d3 VDD Y GND C B A
M1 N_18 B N_19 GND mn15  l=0.13u w=0.46u m=1
M2 N_19 B N_18 GND mn15  l=0.13u w=0.46u m=1
M3 N_18 B N_19 GND mn15  l=0.13u w=0.46u m=1
M4 N_18 B N_19 GND mn15  l=0.13u w=0.46u m=1
M5 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_19 GND mn15  l=0.13u w=0.46u m=1
M7 N_19 A GND GND mn15  l=0.13u w=0.46u m=1
M8 GND A N_19 GND mn15  l=0.13u w=0.46u m=1
M9 Y C N_18 GND mn15  l=0.13u w=0.46u m=1
M10 Y C N_18 GND mn15  l=0.13u w=0.46u m=1
M11 N_18 C Y GND mn15  l=0.13u w=0.46u m=1
M12 N_18 C Y GND mn15  l=0.13u w=0.46u m=1
M13 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M14 VDD B Y VDD mp15  l=0.13u w=0.54u m=1
M15 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M16 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M17 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
M18 Y A VDD VDD mp15  l=0.13u w=0.54u m=1
M19 VDD A Y VDD mp15  l=0.13u w=0.54u m=1
M20 Y A VDD VDD mp15  l=0.13u w=0.54u m=1
M21 VDD C Y VDD mp15  l=0.13u w=0.54u m=1
M22 VDD C Y VDD mp15  l=0.13u w=0.54u m=1
M23 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M24 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
.ends nd03d3
* SPICE INPUT		Tue Jul 31 19:48:12 2018	nd03od
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd03od
.subckt nd03od GND Y VDD A B C
M1 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_7 C N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 N_6 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 B N_7 GND mn15  l=0.13u w=0.26u m=1
M6 N_6 C VDD VDD mp15  l=0.13u w=0.31u m=1
M7 N_5 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_6 A VDD VDD mp15  l=0.13u w=0.31u m=1
M9 N_6 B VDD VDD mp15  l=0.13u w=0.31u m=1
.ends nd03od
* SPICE INPUT		Tue Jul 31 19:48:25 2018	nd04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d0
.subckt nd04d0 VDD Y GND D C B A
M1 N_17 C N_15 GND mn15  l=0.13u w=0.26u m=1
M2 Y D N_15 GND mn15  l=0.13u w=0.26u m=1
M3 N_17 B N_16 GND mn15  l=0.13u w=0.26u m=1
M4 N_16 A GND GND mn15  l=0.13u w=0.26u m=1
M5 VDD C Y VDD mp15  l=0.13u w=0.29u m=1
M6 Y D VDD VDD mp15  l=0.13u w=0.29u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.29u m=1
M8 Y A VDD VDD mp15  l=0.13u w=0.29u m=1
.ends nd04d0
* SPICE INPUT		Tue Jul 31 19:48:38 2018	nd04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d1
.subckt nd04d1 Y VDD A D C B GND
M1 Y D N_15 GND mn15  l=0.13u w=0.46u m=1
M2 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_17 B N_16 GND mn15  l=0.13u w=0.46u m=1
M4 N_17 C N_15 GND mn15  l=0.13u w=0.46u m=1
M5 VDD D Y VDD mp15  l=0.13u w=0.52u m=1
M6 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M7 VDD B Y VDD mp15  l=0.13u w=0.52u m=1
M8 VDD C Y VDD mp15  l=0.13u w=0.52u m=1
.ends nd04d1
* SPICE INPUT		Tue Jul 31 19:48:51 2018	nd04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d2
.subckt nd04d2 VDD Y GND D C B A
M1 N_12 C N_15 GND mn15  l=0.13u w=0.46u m=1
M2 N_12 C N_15 GND mn15  l=0.13u w=0.46u m=1
M3 N_12 D Y GND mn15  l=0.13u w=0.46u m=1
M4 N_12 D Y GND mn15  l=0.13u w=0.46u m=1
M5 N_16 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_16 GND mn15  l=0.13u w=0.46u m=1
M7 N_16 B N_15 GND mn15  l=0.13u w=0.46u m=1
M8 N_16 B N_15 GND mn15  l=0.13u w=0.46u m=1
M9 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M10 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M11 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M12 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M14 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M15 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M16 VDD D Y VDD mp15  l=0.13u w=0.52u m=1
.ends nd04d2
* SPICE INPUT		Tue Jul 31 19:49:04 2018	nd04d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd04d3
.subckt nd04d3 GND VDD Y D C B A
M1 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M2 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M3 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M6 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M7 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M9 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M10 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M11 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M12 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M13 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M14 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M15 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M16 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M17 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M18 VDD B Y VDD mp15  l=0.13u w=0.52u m=1
M19 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M20 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M21 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M22 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M23 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M24 Y A VDD VDD mp15  l=0.13u w=0.52u m=1
M25 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M26 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M27 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M28 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M29 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M30 VDD D Y VDD mp15  l=0.13u w=0.52u m=1
M31 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M32 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
.ends nd04d3
* SPICE INPUT		Tue Jul 31 19:49:18 2018	nd12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d0
.subckt nd12d0 Y GND B VDD AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 GND N_3 N_5 GND mn15  l=0.13u w=0.26u m=1
M3 Y B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_3 AN VDD VDD mp15  l=0.13u w=0.4u m=1
M5 VDD N_3 Y VDD mp15  l=0.13u w=0.35u m=1
M6 Y B VDD VDD mp15  l=0.13u w=0.35u m=1
.ends nd12d0
* SPICE INPUT		Tue Jul 31 19:49:31 2018	nd12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d1
.subckt nd12d1 Y GND VDD B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.3u m=1
M2 GND N_3 N_5 GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_5 GND mn15  l=0.13u w=0.46u m=1
M4 VDD AN N_3 VDD mp15  l=0.13u w=0.45u m=1
M5 VDD N_3 Y VDD mp15  l=0.13u w=0.63u m=1
M6 VDD B Y VDD mp15  l=0.13u w=0.63u m=1
.ends nd12d1
* SPICE INPUT		Tue Jul 31 19:49:43 2018	nd12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d2
.subckt nd12d2 GND Y VDD B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.46u m=1
M2 N_7 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y B N_6 GND mn15  l=0.13u w=0.46u m=1
M4 Y B N_7 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_3 N_6 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M7 Y N_3 VDD VDD mp15  l=0.13u w=0.63u m=1
M8 VDD B Y VDD mp15  l=0.13u w=0.63u m=1
M9 Y B VDD VDD mp15  l=0.13u w=0.63u m=1
M10 Y N_3 VDD VDD mp15  l=0.13u w=0.63u m=1
.ends nd12d2
* SPICE INPUT		Tue Jul 31 19:49:56 2018	nd12d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12d3
.subckt nd12d3 GND Y VDD B AN
M1 GND AN N_4 GND mn15  l=0.13u w=0.4u m=1
M2 N_4 AN GND GND mn15  l=0.13u w=0.4u m=1
M3 N_10 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_11 B Y GND mn15  l=0.13u w=0.46u m=1
M5 Y B N_10 GND mn15  l=0.13u w=0.46u m=1
M6 Y B N_9 GND mn15  l=0.13u w=0.46u m=1
M7 Y B N_12 GND mn15  l=0.13u w=0.46u m=1
M8 GND N_4 N_9 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_11 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M11 VDD AN N_4 VDD mp15  l=0.13u w=0.55u m=1
M12 N_4 AN VDD VDD mp15  l=0.13u w=0.55u m=1
M13 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M14 Y B VDD VDD mp15  l=0.13u w=0.61u m=1
M15 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M16 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M17 VDD B Y VDD mp15  l=0.13u w=0.61u m=1
M18 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
M19 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M20 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
.ends nd12d3
* SPICE INPUT		Tue Jul 31 19:50:08 2018	nd12dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd12dm
.subckt nd12dm Y GND AN VDD B
M1 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y B N_5 GND mn15  l=0.13u w=0.36u m=1
M3 GND N_3 N_5 GND mn15  l=0.13u w=0.36u m=1
M4 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
M5 VDD B Y VDD mp15  l=0.13u w=0.45u m=1
M6 VDD N_3 Y VDD mp15  l=0.13u w=0.45u m=1
.ends nd12dm
* SPICE INPUT		Tue Jul 31 19:50:21 2018	nd13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d0
.subckt nd13d0 Y GND AN C B VDD
M1 N_6 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M2 Y C N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_6 B N_5 GND mn15  l=0.13u w=0.26u m=1
M4 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M5 Y N_3 VDD VDD mp15  l=0.13u w=0.31u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.31u m=1
M7 Y B VDD VDD mp15  l=0.13u w=0.31u m=1
M8 N_3 AN VDD VDD mp15  l=0.13u w=0.4u m=1
.ends nd13d0
* SPICE INPUT		Tue Jul 31 19:50:34 2018	nd13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d1
.subckt nd13d1 Y GND C VDD B AN
M1 N_6 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M2 Y C N_5 GND mn15  l=0.13u w=0.46u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.3u m=1
M4 N_6 B N_5 GND mn15  l=0.13u w=0.46u m=1
M5 Y N_3 VDD VDD mp15  l=0.13u w=0.56u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.56u m=1
M7 VDD AN N_3 VDD mp15  l=0.13u w=0.45u m=1
M8 Y B VDD VDD mp15  l=0.13u w=0.56u m=1
.ends nd13d1
* SPICE INPUT		Tue Jul 31 19:50:47 2018	nd13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d2
.subckt nd13d2 GND Y VDD B C AN
M1 N_9 B N_6 GND mn15  l=0.13u w=0.46u m=1
M2 GND N_4 N_6 GND mn15  l=0.13u w=0.46u m=1
M3 N_4 AN GND GND mn15  l=0.13u w=0.36u m=1
M4 N_8 B N_7 GND mn15  l=0.13u w=0.46u m=1
M5 N_7 N_4 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_9 C Y GND mn15  l=0.13u w=0.46u m=1
M7 N_8 C Y GND mn15  l=0.13u w=0.46u m=1
M8 VDD B Y VDD mp15  l=0.13u w=0.56u m=1
M9 VDD N_4 Y VDD mp15  l=0.13u w=0.56u m=1
M10 N_4 AN VDD VDD mp15  l=0.13u w=0.55u m=1
M11 Y B VDD VDD mp15  l=0.13u w=0.56u m=1
M12 Y N_4 VDD VDD mp15  l=0.13u w=0.56u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.56u m=1
M14 Y C VDD VDD mp15  l=0.13u w=0.56u m=1
.ends nd13d2
* SPICE INPUT		Tue Jul 31 19:51:00 2018	nd13d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd13d3
.subckt nd13d3 Y VDD AN B GND C
M1 N_5 AN GND GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 N_18 GND mn15  l=0.13u w=0.46u m=1
M3 GND N_5 N_18 GND mn15  l=0.13u w=0.46u m=1
M4 GND N_5 N_18 GND mn15  l=0.13u w=0.46u m=1
M5 N_18 N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_21 B N_18 GND mn15  l=0.13u w=0.46u m=1
M7 N_21 B N_18 GND mn15  l=0.13u w=0.46u m=1
M8 N_21 B N_18 GND mn15  l=0.13u w=0.46u m=1
M9 N_21 B N_18 GND mn15  l=0.13u w=0.46u m=1
M10 N_21 C Y GND mn15  l=0.13u w=0.46u m=1
M11 N_21 C Y GND mn15  l=0.13u w=0.46u m=1
M12 N_21 C Y GND mn15  l=0.13u w=0.46u m=1
M13 N_21 C Y GND mn15  l=0.13u w=0.46u m=1
M14 N_5 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_5 Y VDD mp15  l=0.13u w=0.54u m=1
M16 VDD N_5 Y VDD mp15  l=0.13u w=0.54u m=1
M17 VDD N_5 Y VDD mp15  l=0.13u w=0.54u m=1
M18 Y N_5 VDD VDD mp15  l=0.13u w=0.54u m=1
M19 VDD B Y VDD mp15  l=0.13u w=0.54u m=1
M20 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M21 VDD B Y VDD mp15  l=0.13u w=0.54u m=1
M22 Y B VDD VDD mp15  l=0.13u w=0.54u m=1
M23 VDD C Y VDD mp15  l=0.13u w=0.54u m=1
M24 VDD C Y VDD mp15  l=0.13u w=0.54u m=1
M25 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
M26 Y C VDD VDD mp15  l=0.13u w=0.54u m=1
.ends nd13d3
* SPICE INPUT		Tue Jul 31 19:51:13 2018	nd14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d0
.subckt nd14d0 Y GND VDD D C B AN
M1 N_7 C N_5 GND mn15  l=0.13u w=0.26u m=1
M2 Y D N_5 GND mn15  l=0.13u w=0.26u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 B N_6 GND mn15  l=0.13u w=0.26u m=1
M5 N_6 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M6 VDD C Y VDD mp15  l=0.13u w=0.29u m=1
M7 Y D VDD VDD mp15  l=0.13u w=0.29u m=1
M8 N_3 AN VDD VDD mp15  l=0.13u w=0.4u m=1
M9 Y B VDD VDD mp15  l=0.13u w=0.29u m=1
M10 Y N_3 VDD VDD mp15  l=0.13u w=0.29u m=1
.ends nd14d0
* SPICE INPUT		Tue Jul 31 19:51:27 2018	nd14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d1
.subckt nd14d1 Y GND VDD D C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.3u m=1
M2 N_7 C N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_7 B N_6 GND mn15  l=0.13u w=0.46u m=1
M4 Y D N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_6 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 AN VDD VDD mp15  l=0.13u w=0.45u m=1
M7 VDD C Y VDD mp15  l=0.13u w=0.52u m=1
M8 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M9 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M10 Y N_3 VDD VDD mp15  l=0.13u w=0.52u m=1
.ends nd14d1
* SPICE INPUT		Tue Jul 31 19:51:39 2018	nd14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d2
.subckt nd14d2 VDD Y GND D C B AN
M1 N_3 AN GND GND mn15  l=0.13u w=0.4u m=1
M2 N_18 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND N_3 N_18 GND mn15  l=0.13u w=0.46u m=1
M4 N_18 B N_17 GND mn15  l=0.13u w=0.46u m=1
M5 N_18 B N_17 GND mn15  l=0.13u w=0.46u m=1
M6 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M7 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_14 C N_17 GND mn15  l=0.13u w=0.46u m=1
M9 N_14 C N_17 GND mn15  l=0.13u w=0.46u m=1
M10 N_3 AN VDD VDD mp15  l=0.13u w=0.6u m=1
M11 Y D VDD VDD mp15  l=0.13u w=0.52u m=1
M12 VDD D Y VDD mp15  l=0.13u w=0.52u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M14 Y C VDD VDD mp15  l=0.13u w=0.52u m=1
M15 Y N_3 VDD VDD mp15  l=0.13u w=0.52u m=1
M16 Y N_3 VDD VDD mp15  l=0.13u w=0.52u m=1
M17 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
M18 Y B VDD VDD mp15  l=0.13u w=0.52u m=1
.ends nd14d2
* SPICE INPUT		Tue Jul 31 19:51:53 2018	nd14d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd14d3
.subckt nd14d3 GND VDD Y D C B AN
M1 GND AN N_12 GND mn15  l=0.13u w=0.4u m=1
M2 GND AN N_12 GND mn15  l=0.13u w=0.4u m=1
M3 N_11 N_12 GND GND mn15  l=0.13u w=0.46u m=1
M4 GND N_12 N_11 GND mn15  l=0.13u w=0.46u m=1
M5 N_11 N_12 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_12 N_11 GND mn15  l=0.13u w=0.46u m=1
M7 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M8 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M9 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M10 N_11 B N_10 GND mn15  l=0.13u w=0.46u m=1
M11 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M12 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M13 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M14 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M15 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M16 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M17 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M18 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M19 VDD AN N_12 VDD mp15  l=0.13u w=0.58u m=1
M20 VDD AN N_12 VDD mp15  l=0.13u w=0.58u m=1
M21 VDD N_12 Y VDD mp15  l=0.13u w=0.5u m=1
M22 Y N_12 VDD VDD mp15  l=0.13u w=0.5u m=1
M23 VDD N_12 Y VDD mp15  l=0.13u w=0.5u m=1
M24 Y N_12 VDD VDD mp15  l=0.13u w=0.5u m=1
M25 Y B VDD VDD mp15  l=0.13u w=0.5u m=1
M26 Y B VDD VDD mp15  l=0.13u w=0.5u m=1
M27 Y B VDD VDD mp15  l=0.13u w=0.5u m=1
M28 Y B VDD VDD mp15  l=0.13u w=0.5u m=1
M29 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M30 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M31 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M32 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M33 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M34 VDD D Y VDD mp15  l=0.13u w=0.5u m=1
M35 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M36 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
.ends nd14d3
* SPICE INPUT		Tue Jul 31 19:52:07 2018	nd24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d0
.subckt nd24d0 Y GND BN D AN VDD C
M1 N_9 N_5 N_8 GND mn15  l=0.13u w=0.26u m=1
M2 N_9 C N_7 GND mn15  l=0.13u w=0.26u m=1
M3 N_8 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 D Y GND mn15  l=0.13u w=0.26u m=1
M5 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M6 GND BN N_5 GND mn15  l=0.13u w=0.26u m=1
M7 N_5 BN VDD VDD mp15  l=0.13u w=0.4u m=1
M8 VDD N_5 Y VDD mp15  l=0.13u w=0.29u m=1
M9 Y C VDD VDD mp15  l=0.13u w=0.29u m=1
M10 Y N_3 VDD VDD mp15  l=0.13u w=0.29u m=1
M11 Y D VDD VDD mp15  l=0.13u w=0.29u m=1
M12 N_3 AN VDD VDD mp15  l=0.13u w=0.4u m=1
.ends nd24d0
* SPICE INPUT		Tue Jul 31 19:52:20 2018	nd24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d1
.subckt nd24d1 GND Y BN AN D C VDD
M1 GND BN N_2 GND mn15  l=0.13u w=0.3u m=1
M2 GND AN N_5 GND mn15  l=0.13u w=0.3u m=1
M3 N_8 N_5 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_9 N_2 N_8 GND mn15  l=0.13u w=0.46u m=1
M5 N_9 C N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_7 D Y GND mn15  l=0.13u w=0.46u m=1
M7 N_2 BN VDD VDD mp15  l=0.13u w=0.43u m=1
M8 VDD AN N_5 VDD mp15  l=0.13u w=0.43u m=1
M9 Y N_5 VDD VDD mp15  l=0.13u w=0.5u m=1
M10 Y N_2 VDD VDD mp15  l=0.13u w=0.5u m=1
M11 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M12 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
.ends nd24d1
* SPICE INPUT		Tue Jul 31 19:52:33 2018	nd24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d2
.subckt nd24d2 GND Y BN AN VDD D C
M1 N_3 AN GND GND mn15  l=0.13u w=0.4u m=1
M2 N_4 BN GND GND mn15  l=0.13u w=0.4u m=1
M3 N_6 N_4 N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_6 N_4 N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_6 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_3 N_6 GND mn15  l=0.13u w=0.46u m=1
M7 N_11 C N_5 GND mn15  l=0.13u w=0.46u m=1
M8 N_11 C N_5 GND mn15  l=0.13u w=0.46u m=1
M9 N_11 D Y GND mn15  l=0.13u w=0.46u m=1
M10 N_11 D Y GND mn15  l=0.13u w=0.46u m=1
M11 N_3 AN VDD VDD mp15  l=0.13u w=0.58u m=1
M12 N_4 BN VDD VDD mp15  l=0.13u w=0.58u m=1
M13 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M14 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M15 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M16 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M17 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M18 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M19 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M20 VDD D Y VDD mp15  l=0.13u w=0.5u m=1
.ends nd24d2
* SPICE INPUT		Tue Jul 31 19:52:46 2018	nd24d3
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nd24d3
.subckt nd24d3 VDD Y GND D C AN BN
M1 N_4 BN GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.46u m=1
M3 N_27 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_27 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_27 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_27 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_27 N_4 N_26 GND mn15  l=0.13u w=0.46u m=1
M8 N_27 N_4 N_26 GND mn15  l=0.13u w=0.46u m=1
M9 N_27 N_4 N_26 GND mn15  l=0.13u w=0.46u m=1
M10 N_27 N_4 N_26 GND mn15  l=0.13u w=0.46u m=1
M11 N_23 C N_26 GND mn15  l=0.13u w=0.46u m=1
M12 N_23 C N_26 GND mn15  l=0.13u w=0.46u m=1
M13 N_23 C N_26 GND mn15  l=0.13u w=0.46u m=1
M14 N_23 C N_26 GND mn15  l=0.13u w=0.46u m=1
M15 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M16 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M17 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M18 N_23 D Y GND mn15  l=0.13u w=0.46u m=1
M19 N_4 BN VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_3 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M21 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M22 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M23 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M24 Y N_3 VDD VDD mp15  l=0.13u w=0.5u m=1
M25 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M26 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M27 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M28 Y N_4 VDD VDD mp15  l=0.13u w=0.5u m=1
M29 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M30 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M31 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M32 Y C VDD VDD mp15  l=0.13u w=0.5u m=1
M33 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M34 VDD D Y VDD mp15  l=0.13u w=0.5u m=1
M35 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
M36 Y D VDD VDD mp15  l=0.13u w=0.5u m=1
.ends nd24d3
* SPICE INPUT		Tue Jul 31 19:52:58 2018	nr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d0
.subckt nr02d0 Y GND VDD B A
M1 GND B Y GND mn15  l=0.13u w=0.26u m=1
M2 GND A Y GND mn15  l=0.13u w=0.26u m=1
M3 Y B N_8 VDD mp15  l=0.13u w=0.4u m=1
M4 VDD A N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends nr02d0
* SPICE INPUT		Tue Jul 31 19:53:11 2018	nr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d1
.subckt nr02d1 Y GND VDD B A
M1 GND B Y GND mn15  l=0.13u w=0.34u m=1
M2 GND A Y GND mn15  l=0.13u w=0.34u m=1
M3 Y B N_8 VDD mp15  l=0.13u w=0.69u m=1
M4 VDD A N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends nr02d1
* SPICE INPUT		Tue Jul 31 19:53:24 2018	nr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d2
.subckt nr02d2 VDD Y GND A B
M1 GND B Y GND mn15  l=0.13u w=0.34u m=1
M2 Y B GND GND mn15  l=0.13u w=0.34u m=1
M3 Y A GND GND mn15  l=0.13u w=0.34u m=1
M4 GND A Y GND mn15  l=0.13u w=0.34u m=1
M5 Y B N_5 VDD mp15  l=0.13u w=0.69u m=1
M6 Y B N_6 VDD mp15  l=0.13u w=0.69u m=1
M7 N_6 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 VDD A N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends nr02d2
* SPICE INPUT		Tue Jul 31 19:53:38 2018	nr02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02d4
.subckt nr02d4 Y GND VDD B A
M1 GND A Y GND mn15  l=0.13u w=0.34u m=1
M2 Y A GND GND mn15  l=0.13u w=0.34u m=1
M3 GND A Y GND mn15  l=0.13u w=0.34u m=1
M4 Y A GND GND mn15  l=0.13u w=0.34u m=1
M5 GND B Y GND mn15  l=0.13u w=0.34u m=1
M6 GND B Y GND mn15  l=0.13u w=0.34u m=1
M7 GND B Y GND mn15  l=0.13u w=0.34u m=1
M8 Y B GND GND mn15  l=0.13u w=0.34u m=1
M9 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M13 Y B N_13 VDD mp15  l=0.13u w=0.69u m=1
M14 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M16 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
.ends nr02d4
* SPICE INPUT		Tue Jul 31 19:53:50 2018	nr02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr02dm
.subckt nr02dm Y GND VDD B A
M1 GND B Y GND mn15  l=0.13u w=0.27u m=1
M2 GND A Y GND mn15  l=0.13u w=0.27u m=1
M3 Y B N_8 VDD mp15  l=0.13u w=0.55u m=1
M4 VDD A N_8 VDD mp15  l=0.13u w=0.55u m=1
.ends nr02dm
* SPICE INPUT		Tue Jul 31 19:54:03 2018	nr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d0
.subckt nr03d0 GND Y VDD C B A
M1 Y C GND GND mn15  l=0.13u w=0.26u m=1
M2 Y B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y A GND GND mn15  l=0.13u w=0.26u m=1
M4 Y C N_16 VDD mp15  l=0.13u w=0.4u m=1
M5 N_17 B N_16 VDD mp15  l=0.13u w=0.4u m=1
M6 N_17 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends nr03d0
* SPICE INPUT		Tue Jul 31 19:54:17 2018	nr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d1
.subckt nr03d1 Y VDD GND C B A
M1 Y C GND GND mn15  l=0.13u w=0.29u m=1
M2 Y B GND GND mn15  l=0.13u w=0.29u m=1
M3 Y A GND GND mn15  l=0.13u w=0.29u m=1
M4 Y C N_4 VDD mp15  l=0.13u w=0.69u m=1
M5 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M6 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nr03d1
* SPICE INPUT		Tue Jul 31 19:54:29 2018	nr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d2
.subckt nr03d2 Y VDD GND C B A
M1 Y A GND GND mn15  l=0.13u w=0.29u m=1
M2 Y A GND GND mn15  l=0.13u w=0.29u m=1
M3 GND B Y GND mn15  l=0.13u w=0.29u m=1
M4 Y C GND GND mn15  l=0.13u w=0.29u m=1
M5 Y B GND GND mn15  l=0.13u w=0.29u m=1
M6 GND C Y GND mn15  l=0.13u w=0.29u m=1
M7 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_12 B N_9 VDD mp15  l=0.13u w=0.69u m=1
M10 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M12 Y C N_9 VDD mp15  l=0.13u w=0.69u m=1
.ends nr03d2
* SPICE INPUT		Tue Jul 31 19:54:42 2018	nr03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr03d4
.subckt nr03d4 Y GND VDD C B A
M1 GND A Y GND mn15  l=0.13u w=0.29u m=1
M2 GND A Y GND mn15  l=0.13u w=0.29u m=1
M3 GND A Y GND mn15  l=0.13u w=0.29u m=1
M4 Y A GND GND mn15  l=0.13u w=0.29u m=1
M5 GND C Y GND mn15  l=0.13u w=0.29u m=1
M6 GND C Y GND mn15  l=0.13u w=0.29u m=1
M7 GND C Y GND mn15  l=0.13u w=0.29u m=1
M8 Y C GND GND mn15  l=0.13u w=0.29u m=1
M9 GND B Y GND mn15  l=0.13u w=0.29u m=1
M10 Y B GND GND mn15  l=0.13u w=0.29u m=1
M11 GND B Y GND mn15  l=0.13u w=0.29u m=1
M12 Y B GND GND mn15  l=0.13u w=0.29u m=1
M13 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_18 C Y VDD mp15  l=0.13u w=0.69u m=1
M18 N_18 C Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_18 C Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y C N_18 VDD mp15  l=0.13u w=0.69u m=1
M21 N_18 B N_20 VDD mp15  l=0.13u w=0.69u m=1
M22 N_20 B N_18 VDD mp15  l=0.13u w=0.69u m=1
M23 N_18 B N_20 VDD mp15  l=0.13u w=0.69u m=1
M24 N_20 B N_18 VDD mp15  l=0.13u w=0.69u m=1
.ends nr03d4
* SPICE INPUT		Tue Jul 31 19:54:55 2018	nr04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d0
.subckt nr04d0 GND Y VDD D C B A
M1 Y A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y D GND GND mn15  l=0.13u w=0.26u m=1
M4 Y C GND GND mn15  l=0.13u w=0.26u m=1
M5 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_14 B N_13 VDD mp15  l=0.13u w=0.4u m=1
M7 Y D N_12 VDD mp15  l=0.13u w=0.4u m=1
M8 N_14 C N_12 VDD mp15  l=0.13u w=0.4u m=1
.ends nr04d0
* SPICE INPUT		Tue Jul 31 19:55:08 2018	nr04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d1
.subckt nr04d1 Y VDD GND D C B A
M1 GND D Y GND mn15  l=0.13u w=0.28u m=1
M2 Y A GND GND mn15  l=0.13u w=0.28u m=1
M3 GND B Y GND mn15  l=0.13u w=0.28u m=1
M4 GND C Y GND mn15  l=0.13u w=0.28u m=1
M5 Y D N_4 VDD mp15  l=0.13u w=0.69u m=1
M6 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_6 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M8 N_6 C N_4 VDD mp15  l=0.13u w=0.69u m=1
.ends nr04d1
* SPICE INPUT		Tue Jul 31 19:55:21 2018	nr04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d2
.subckt nr04d2 GND Y VDD D C B A
M1 Y D GND GND mn15  l=0.13u w=0.28u m=1
M2 GND D Y GND mn15  l=0.13u w=0.28u m=1
M3 Y C GND GND mn15  l=0.13u w=0.28u m=1
M4 Y C GND GND mn15  l=0.13u w=0.28u m=1
M5 Y B GND GND mn15  l=0.13u w=0.28u m=1
M6 Y B GND GND mn15  l=0.13u w=0.28u m=1
M7 Y A GND GND mn15  l=0.13u w=0.28u m=1
M8 Y A GND GND mn15  l=0.13u w=0.28u m=1
M9 N_16 B N_15 VDD mp15  l=0.13u w=0.69u m=1
M10 N_16 B N_15 VDD mp15  l=0.13u w=0.69u m=1
M11 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_16 VDD mp15  l=0.13u w=0.69u m=1
M13 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_12 C N_15 VDD mp15  l=0.13u w=0.69u m=1
M16 N_15 C N_12 VDD mp15  l=0.13u w=0.69u m=1
.ends nr04d2
* SPICE INPUT		Tue Jul 31 19:55:34 2018	nr04d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr04d4
.subckt nr04d4 VDD Y GND D C B A
M1 Y B GND GND mn15  l=0.13u w=0.28u m=1
M2 Y B GND GND mn15  l=0.13u w=0.28u m=1
M3 Y B GND GND mn15  l=0.13u w=0.28u m=1
M4 Y B GND GND mn15  l=0.13u w=0.28u m=1
M5 Y C GND GND mn15  l=0.13u w=0.28u m=1
M6 Y C GND GND mn15  l=0.13u w=0.28u m=1
M7 Y C GND GND mn15  l=0.13u w=0.28u m=1
M8 Y C GND GND mn15  l=0.13u w=0.28u m=1
M9 Y D GND GND mn15  l=0.13u w=0.28u m=1
M10 GND D Y GND mn15  l=0.13u w=0.28u m=1
M11 Y D GND GND mn15  l=0.13u w=0.28u m=1
M12 Y D GND GND mn15  l=0.13u w=0.28u m=1
M13 Y A GND GND mn15  l=0.13u w=0.28u m=1
M14 Y A GND GND mn15  l=0.13u w=0.28u m=1
M15 Y A GND GND mn15  l=0.13u w=0.28u m=1
M16 Y A GND GND mn15  l=0.13u w=0.28u m=1
M17 N_3 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M18 N_3 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M19 N_3 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M20 N_2 B N_3 VDD mp15  l=0.13u w=0.69u m=1
M21 N_3 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD A N_3 VDD mp15  l=0.13u w=0.69u m=1
M23 N_3 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 VDD A N_3 VDD mp15  l=0.13u w=0.69u m=1
M25 N_12 C N_2 VDD mp15  l=0.13u w=0.69u m=1
M26 N_2 C N_12 VDD mp15  l=0.13u w=0.69u m=1
M27 N_12 C N_2 VDD mp15  l=0.13u w=0.69u m=1
M28 N_2 C N_12 VDD mp15  l=0.13u w=0.69u m=1
M29 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M31 N_12 D Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y D N_12 VDD mp15  l=0.13u w=0.69u m=1
.ends nr04d4
* SPICE INPUT		Tue Jul 31 19:55:46 2018	nr12d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d0
.subckt nr12d0 Y VDD GND B AN
M1 GND N_3 Y GND mn15  l=0.13u w=0.26u m=1
M2 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M3 GND B Y GND mn15  l=0.13u w=0.26u m=1
M4 VDD N_3 N_5 VDD mp15  l=0.13u w=0.4u m=1
M5 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
M6 Y B N_5 VDD mp15  l=0.13u w=0.4u m=1
.ends nr12d0
* SPICE INPUT		Tue Jul 31 19:55:59 2018	nr12d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d1
.subckt nr12d1 Y VDD GND B AN
M1 GND N_3 Y GND mn15  l=0.13u w=0.34u m=1
M2 GND B Y GND mn15  l=0.13u w=0.34u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.28u m=1
M4 VDD N_3 N_5 VDD mp15  l=0.13u w=0.69u m=1
M5 Y B N_5 VDD mp15  l=0.13u w=0.69u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.42u m=1
.ends nr12d1
* SPICE INPUT		Tue Jul 31 19:56:11 2018	nr12d1p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d1p5
.subckt nr12d1p5 Y VDD GND B AN
M1 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND B Y GND mn15  l=0.13u w=0.46u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.42u m=1
M4 VDD N_3 N_5 VDD mp15  l=0.13u w=0.69u m=1
M5 Y B N_5 VDD mp15  l=0.13u w=0.69u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.52u m=1
.ends nr12d1p5
* SPICE INPUT		Tue Jul 31 19:56:24 2018	nr12d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d2
.subckt nr12d2 VDD Y GND B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.34u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.34u m=1
M3 GND B Y GND mn15  l=0.13u w=0.34u m=1
M4 Y B GND GND mn15  l=0.13u w=0.34u m=1
M5 Y N_3 GND GND mn15  l=0.13u w=0.34u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.52u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y B N_6 VDD mp15  l=0.13u w=0.69u m=1
M9 Y B N_7 VDD mp15  l=0.13u w=0.69u m=1
M10 N_6 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nr12d2
* SPICE INPUT		Tue Jul 31 19:56:37 2018	nr12d2p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d2p5
.subckt nr12d2p5 VDD Y GND B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.46u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND B Y GND mn15  l=0.13u w=0.46u m=1
M4 Y B GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.69u m=1
M7 N_7 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y B N_6 VDD mp15  l=0.13u w=0.69u m=1
M9 Y B N_7 VDD mp15  l=0.13u w=0.69u m=1
M10 N_6 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends nr12d2p5
* SPICE INPUT		Tue Jul 31 19:56:51 2018	nr12d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12d4
.subckt nr12d4 Y GND VDD B AN
M1 GND B Y GND mn15  l=0.13u w=0.34u m=1
M2 GND B Y GND mn15  l=0.13u w=0.34u m=1
M3 GND B Y GND mn15  l=0.13u w=0.34u m=1
M4 Y B GND GND mn15  l=0.13u w=0.34u m=1
M5 N_5 AN GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.34u m=1
M7 Y N_5 GND GND mn15  l=0.13u w=0.34u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.34u m=1
M9 Y N_5 GND GND mn15  l=0.13u w=0.34u m=1
M10 VDD AN N_5 VDD mp15  l=0.13u w=0.69u m=1
M11 Y B N_14 VDD mp15  l=0.13u w=0.69u m=1
M12 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M13 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M15 N_14 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
M17 N_14 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
.ends nr12d4
* SPICE INPUT		Tue Jul 31 19:57:05 2018	nr12dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr12dm
.subckt nr12dm Y VDD GND B AN
M1 GND N_3 Y GND mn15  l=0.13u w=0.27u m=1
M2 GND B Y GND mn15  l=0.13u w=0.27u m=1
M3 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M4 VDD N_3 N_5 VDD mp15  l=0.13u w=0.55u m=1
M5 Y B N_5 VDD mp15  l=0.13u w=0.55u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
.ends nr12dm
* SPICE INPUT		Tue Jul 31 19:57:18 2018	nr13d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d0
.subckt nr13d0 Y VDD GND C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 Y B GND GND mn15  l=0.13u w=0.26u m=1
M4 Y C GND GND mn15  l=0.13u w=0.26u m=1
M5 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
M6 N_8 N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_8 B N_7 VDD mp15  l=0.13u w=0.4u m=1
M8 Y C N_7 VDD mp15  l=0.13u w=0.4u m=1
.ends nr13d0
* SPICE INPUT		Tue Jul 31 19:57:31 2018	nr13d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d1
.subckt nr13d1 Y VDD GND C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.28u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.29u m=1
M3 Y B GND GND mn15  l=0.13u w=0.29u m=1
M4 Y C GND GND mn15  l=0.13u w=0.29u m=1
M5 VDD AN N_3 VDD mp15  l=0.13u w=0.42u m=1
M6 N_8 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_8 B N_7 VDD mp15  l=0.13u w=0.69u m=1
M8 Y C N_7 VDD mp15  l=0.13u w=0.69u m=1
.ends nr13d1
* SPICE INPUT		Tue Jul 31 19:57:44 2018	nr13d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d2
.subckt nr13d2 Y GND VDD C B AN
M1 Y B GND GND mn15  l=0.13u w=0.29u m=1
M2 Y B GND GND mn15  l=0.13u w=0.29u m=1
M3 Y N_5 GND GND mn15  l=0.13u w=0.29u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.29u m=1
M5 N_5 AN GND GND mn15  l=0.13u w=0.33u m=1
M6 GND C Y GND mn15  l=0.13u w=0.29u m=1
M7 GND C Y GND mn15  l=0.13u w=0.29u m=1
M8 N_12 B N_14 VDD mp15  l=0.13u w=0.69u m=1
M9 N_14 B N_12 VDD mp15  l=0.13u w=0.69u m=1
M10 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_12 C Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 N_14 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD AN N_5 VDD mp15  l=0.13u w=0.5u m=1
.ends nr13d2
* SPICE INPUT		Tue Jul 31 19:57:57 2018	nr13d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr13d4
.subckt nr13d4 Y GND VDD C B AN
M1 N_5 AN GND GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.29u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.29u m=1
M4 GND N_5 Y GND mn15  l=0.13u w=0.29u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.29u m=1
M6 GND C Y GND mn15  l=0.13u w=0.29u m=1
M7 GND C Y GND mn15  l=0.13u w=0.29u m=1
M8 GND C Y GND mn15  l=0.13u w=0.29u m=1
M9 Y C GND GND mn15  l=0.13u w=0.29u m=1
M10 GND B Y GND mn15  l=0.13u w=0.29u m=1
M11 Y B GND GND mn15  l=0.13u w=0.29u m=1
M12 GND B Y GND mn15  l=0.13u w=0.29u m=1
M13 Y B GND GND mn15  l=0.13u w=0.29u m=1
M14 VDD AN N_5 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_5 N_21 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_5 N_21 VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_5 N_21 VDD mp15  l=0.13u w=0.69u m=1
M18 N_21 N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 Y C N_19 VDD mp15  l=0.13u w=0.69u m=1
M20 N_19 C Y VDD mp15  l=0.13u w=0.69u m=1
M21 N_19 C Y VDD mp15  l=0.13u w=0.69u m=1
M22 N_19 C Y VDD mp15  l=0.13u w=0.69u m=1
M23 N_19 B N_21 VDD mp15  l=0.13u w=0.69u m=1
M24 N_21 B N_19 VDD mp15  l=0.13u w=0.69u m=1
M25 N_19 B N_21 VDD mp15  l=0.13u w=0.69u m=1
M26 N_21 B N_19 VDD mp15  l=0.13u w=0.69u m=1
.ends nr13d4
* SPICE INPUT		Tue Jul 31 19:58:10 2018	nr14d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d0
.subckt nr14d0 Y VDD GND D C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND B Y GND mn15  l=0.13u w=0.26u m=1
M4 GND D Y GND mn15  l=0.13u w=0.26u m=1
M5 GND C Y GND mn15  l=0.13u w=0.26u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.4u m=1
M7 N_9 N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_10 B N_9 VDD mp15  l=0.13u w=0.4u m=1
M9 Y D N_8 VDD mp15  l=0.13u w=0.4u m=1
M10 N_10 C N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends nr14d0
* SPICE INPUT		Tue Jul 31 19:58:23 2018	nr14d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d1
.subckt nr14d1 Y VDD GND D C B AN
M1 GND AN N_3 GND mn15  l=0.13u w=0.28u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M3 GND B Y GND mn15  l=0.13u w=0.28u m=1
M4 GND D Y GND mn15  l=0.13u w=0.28u m=1
M5 GND C Y GND mn15  l=0.13u w=0.28u m=1
M6 VDD AN N_3 VDD mp15  l=0.13u w=0.42u m=1
M7 N_9 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_10 B N_9 VDD mp15  l=0.13u w=0.69u m=1
M9 Y D N_8 VDD mp15  l=0.13u w=0.69u m=1
M10 N_10 C N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends nr14d1
* SPICE INPUT		Tue Jul 31 19:58:36 2018	nr14d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d2
.subckt nr14d2 GND Y VDD D C B AN
M1 Y D GND GND mn15  l=0.13u w=0.28u m=1
M2 GND D Y GND mn15  l=0.13u w=0.28u m=1
M3 Y C GND GND mn15  l=0.13u w=0.28u m=1
M4 Y C GND GND mn15  l=0.13u w=0.28u m=1
M5 Y N_12 GND GND mn15  l=0.13u w=0.28u m=1
M6 Y N_12 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y B GND GND mn15  l=0.13u w=0.28u m=1
M8 Y B GND GND mn15  l=0.13u w=0.28u m=1
M9 N_12 AN GND GND mn15  l=0.13u w=0.33u m=1
M10 N_12 AN VDD VDD mp15  l=0.13u w=0.5u m=1
M11 N_18 N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_12 N_18 VDD mp15  l=0.13u w=0.69u m=1
M13 N_18 B N_17 VDD mp15  l=0.13u w=0.69u m=1
M14 N_18 B N_17 VDD mp15  l=0.13u w=0.69u m=1
M15 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M16 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M17 N_14 C N_17 VDD mp15  l=0.13u w=0.69u m=1
M18 N_17 C N_14 VDD mp15  l=0.13u w=0.69u m=1
.ends nr14d2
* SPICE INPUT		Tue Jul 31 19:58:49 2018	nr14d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr14d4
.subckt nr14d4 VDD Y GND D C B AN
M1 N_2 AN GND GND mn15  l=0.13u w=0.46u m=1
M2 Y N_2 GND GND mn15  l=0.13u w=0.28u m=1
M3 Y N_2 GND GND mn15  l=0.13u w=0.28u m=1
M4 Y N_2 GND GND mn15  l=0.13u w=0.28u m=1
M5 Y N_2 GND GND mn15  l=0.13u w=0.28u m=1
M6 Y B GND GND mn15  l=0.13u w=0.28u m=1
M7 Y B GND GND mn15  l=0.13u w=0.28u m=1
M8 Y B GND GND mn15  l=0.13u w=0.28u m=1
M9 Y B GND GND mn15  l=0.13u w=0.28u m=1
M10 Y C GND GND mn15  l=0.13u w=0.28u m=1
M11 Y C GND GND mn15  l=0.13u w=0.28u m=1
M12 Y C GND GND mn15  l=0.13u w=0.28u m=1
M13 Y C GND GND mn15  l=0.13u w=0.28u m=1
M14 Y D GND GND mn15  l=0.13u w=0.28u m=1
M15 GND D Y GND mn15  l=0.13u w=0.28u m=1
M16 Y D GND GND mn15  l=0.13u w=0.28u m=1
M17 Y D GND GND mn15  l=0.13u w=0.28u m=1
M18 VDD AN N_2 VDD mp15  l=0.13u w=0.69u m=1
M19 N_5 N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_2 N_5 VDD mp15  l=0.13u w=0.69u m=1
M21 N_5 N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_2 N_5 VDD mp15  l=0.13u w=0.69u m=1
M23 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M24 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M25 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M26 N_4 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M27 N_14 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M28 N_4 C N_14 VDD mp15  l=0.13u w=0.69u m=1
M29 N_14 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M30 N_4 C N_14 VDD mp15  l=0.13u w=0.69u m=1
M31 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M32 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M33 N_14 D Y VDD mp15  l=0.13u w=0.69u m=1
M34 Y D N_14 VDD mp15  l=0.13u w=0.69u m=1
.ends nr14d4
* SPICE INPUT		Tue Jul 31 19:59:02 2018	nr24d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d0
.subckt nr24d0 GND Y VDD AN C D BN
M1 N_5 AN GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND N_3 Y GND mn15  l=0.13u w=0.26u m=1
M4 Y C GND GND mn15  l=0.13u w=0.26u m=1
M5 Y D GND GND mn15  l=0.13u w=0.26u m=1
M6 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M7 VDD AN N_5 VDD mp15  l=0.13u w=0.4u m=1
M8 N_15 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_16 N_3 N_15 VDD mp15  l=0.13u w=0.4u m=1
M10 N_16 C N_14 VDD mp15  l=0.13u w=0.4u m=1
M11 N_14 D Y VDD mp15  l=0.13u w=0.4u m=1
M12 VDD BN N_3 VDD mp15  l=0.13u w=0.4u m=1
.ends nr24d0
* SPICE INPUT		Tue Jul 31 19:59:14 2018	nr24d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d1
.subckt nr24d1 GND Y VDD AN C D BN
M1 N_5 AN GND GND mn15  l=0.13u w=0.28u m=1
M2 Y N_5 GND GND mn15  l=0.13u w=0.28u m=1
M3 GND N_3 Y GND mn15  l=0.13u w=0.28u m=1
M4 Y C GND GND mn15  l=0.13u w=0.28u m=1
M5 Y D GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 BN GND GND mn15  l=0.13u w=0.28u m=1
M7 VDD AN N_5 VDD mp15  l=0.13u w=0.42u m=1
M8 N_15 N_5 VDD VDD mp15  l=0.13u w=0.7u m=1
M9 N_16 N_3 N_15 VDD mp15  l=0.13u w=0.7u m=1
M10 N_16 C N_14 VDD mp15  l=0.13u w=0.7u m=1
M11 N_14 D Y VDD mp15  l=0.13u w=0.7u m=1
M12 VDD BN N_3 VDD mp15  l=0.13u w=0.42u m=1
.ends nr24d1
* SPICE INPUT		Tue Jul 31 19:59:27 2018	nr24d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d2
.subckt nr24d2 GND Y VDD C BN AN D
M1 N_4 BN GND GND mn15  l=0.13u w=0.4u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.4u m=1
M3 Y D GND GND mn15  l=0.13u w=0.28u m=1
M4 GND D Y GND mn15  l=0.13u w=0.28u m=1
M5 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M8 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M9 Y C GND GND mn15  l=0.13u w=0.28u m=1
M10 Y C GND GND mn15  l=0.13u w=0.28u m=1
M11 N_4 BN VDD VDD mp15  l=0.13u w=0.6u m=1
M12 N_3 AN VDD VDD mp15  l=0.13u w=0.6u m=1
M13 N_21 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_3 N_21 VDD mp15  l=0.13u w=0.69u m=1
M15 N_21 N_4 N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_21 N_4 N_20 VDD mp15  l=0.13u w=0.69u m=1
M17 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M18 N_19 D Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_19 C N_20 VDD mp15  l=0.13u w=0.69u m=1
M20 N_20 C N_19 VDD mp15  l=0.13u w=0.69u m=1
.ends nr24d2
* SPICE INPUT		Tue Jul 31 19:59:40 2018	nr24d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=nr24d4
.subckt nr24d4 VDD Y GND D C AN BN
M1 N_4 BN GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 AN GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M4 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M5 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M8 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M9 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M10 Y N_4 GND GND mn15  l=0.13u w=0.28u m=1
M11 Y C GND GND mn15  l=0.13u w=0.28u m=1
M12 Y C GND GND mn15  l=0.13u w=0.28u m=1
M13 Y C GND GND mn15  l=0.13u w=0.28u m=1
M14 Y C GND GND mn15  l=0.13u w=0.28u m=1
M15 Y D GND GND mn15  l=0.13u w=0.28u m=1
M16 GND D Y GND mn15  l=0.13u w=0.28u m=1
M17 Y D GND GND mn15  l=0.13u w=0.28u m=1
M18 Y D GND GND mn15  l=0.13u w=0.28u m=1
M19 N_4 BN VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_3 AN VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_6 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_3 N_6 VDD mp15  l=0.13u w=0.69u m=1
M23 N_6 N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_3 N_6 VDD mp15  l=0.13u w=0.69u m=1
M25 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.69u m=1
M26 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.69u m=1
M27 N_6 N_4 N_5 VDD mp15  l=0.13u w=0.69u m=1
M28 N_5 N_4 N_6 VDD mp15  l=0.13u w=0.69u m=1
M29 N_15 C N_5 VDD mp15  l=0.13u w=0.69u m=1
M30 N_5 C N_15 VDD mp15  l=0.13u w=0.69u m=1
M31 N_15 C N_5 VDD mp15  l=0.13u w=0.69u m=1
M32 N_5 C N_15 VDD mp15  l=0.13u w=0.69u m=1
M33 N_15 D Y VDD mp15  l=0.13u w=0.69u m=1
M34 N_15 D Y VDD mp15  l=0.13u w=0.69u m=1
M35 N_15 D Y VDD mp15  l=0.13u w=0.69u m=1
M36 Y D N_15 VDD mp15  l=0.13u w=0.69u m=1
.ends nr24d4
* SPICE INPUT		Tue Jul 31 19:59:53 2018	oai211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d0
.subckt oai211d0 Y GND VDD D C B A
M1 N_4 C N_6 GND mn15  l=0.13u w=0.26u m=1
M2 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M3 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_6 D Y GND mn15  l=0.13u w=0.26u m=1
M5 Y C VDD VDD mp15  l=0.13u w=0.27u m=1
M6 N_13 B Y VDD mp15  l=0.13u w=0.4u m=1
M7 N_13 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 Y D VDD VDD mp15  l=0.13u w=0.27u m=1
.ends oai211d0
* SPICE INPUT		Tue Jul 31 20:00:06 2018	oai211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d1
.subckt oai211d1 Y GND VDD D C B A
M1 N_4 C N_6 GND mn15  l=0.13u w=0.46u m=1
M2 N_4 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M4 Y D N_6 GND mn15  l=0.13u w=0.46u m=1
M5 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M6 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M7 N_14 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oai211d1
* SPICE INPUT		Tue Jul 31 20:00:19 2018	oai211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d2
.subckt oai211d2 GND Y B A D C VDD
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_2 C N_9 GND mn15  l=0.13u w=0.46u m=1
M6 Y D N_9 GND mn15  l=0.13u w=0.46u m=1
M7 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_10 C N_2 GND mn15  l=0.13u w=0.46u m=1
M9 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_21 B Y VDD mp15  l=0.13u w=0.69u m=1
M11 Y B N_20 VDD mp15  l=0.13u w=0.69u m=1
M12 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M14 VDD D Y VDD mp15  l=0.13u w=0.48u m=1
M15 VDD D Y VDD mp15  l=0.13u w=0.48u m=1
M16 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
.ends oai211d2
* SPICE INPUT		Tue Jul 31 20:00:33 2018	oai211d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai211d4
.subckt oai211d4 GND VDD D Y C A B
M1 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_10 B GND GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_10 GND mn15  l=0.13u w=0.46u m=1
M4 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND A N_10 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_10 GND mn15  l=0.13u w=0.46u m=1
M7 GND B N_10 GND mn15  l=0.13u w=0.46u m=1
M8 GND B N_10 GND mn15  l=0.13u w=0.46u m=1
M9 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M10 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M11 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M12 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M13 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M14 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M15 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M16 N_9 C N_10 GND mn15  l=0.13u w=0.46u m=1
M17 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_16 B Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_15 B Y VDD mp15  l=0.13u w=0.69u m=1
M20 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M22 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M23 VDD D Y VDD mp15  l=0.13u w=0.46u m=1
M24 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M25 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M26 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M28 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M29 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M30 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M31 N_18 B Y VDD mp15  l=0.13u w=0.69u m=1
M32 N_17 B Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai211d4
* SPICE INPUT		Tue Jul 31 20:00:46 2018	oai21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d0
.subckt oai21d0 Y GND VDD C B A
M1 GND A N_2 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.26u m=1
M3 Y C N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_20 A VDD VDD mp15  l=0.13u w=0.4u m=1
M5 N_20 B Y VDD mp15  l=0.13u w=0.4u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.27u m=1
.ends oai21d0
* SPICE INPUT		Tue Jul 31 20:00:59 2018	oai21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d1
.subckt oai21d1 Y GND VDD C B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 Y C N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M5 N_20 B Y VDD mp15  l=0.13u w=0.69u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oai21d1
* SPICE INPUT		Tue Jul 31 20:01:12 2018	oai21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d2
.subckt oai21d2 Y VDD GND C A B
M1 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 C Y GND mn15  l=0.13u w=0.46u m=1
M3 N_12 C Y GND mn15  l=0.13u w=0.46u m=1
M4 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND B N_12 GND mn15  l=0.13u w=0.46u m=1
M6 N_12 B GND GND mn15  l=0.13u w=0.46u m=1
M7 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 VDD C Y VDD mp15  l=0.13u w=0.46u m=1
M9 VDD C Y VDD mp15  l=0.13u w=0.46u m=1
M10 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 B Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y B N_7 VDD mp15  l=0.13u w=0.69u m=1
.ends oai21d2
* SPICE INPUT		Tue Jul 31 20:01:25 2018	oai21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21d4
.subckt oai21d4 Y VDD GND C A B
M1 GND A N_20 GND mn15  l=0.13u w=0.46u m=1
M2 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M7 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M8 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M10 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M11 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M12 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M13 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_14 B Y VDD mp15  l=0.13u w=0.69u m=1
M17 Y B N_13 VDD mp15  l=0.13u w=0.69u m=1
M18 N_12 B Y VDD mp15  l=0.13u w=0.69u m=1
M19 Y B N_11 VDD mp15  l=0.13u w=0.69u m=1
M20 N_14 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD C Y VDD mp15  l=0.13u w=0.46u m=1
M22 VDD C Y VDD mp15  l=0.13u w=0.46u m=1
M23 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
M24 Y C VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oai21d4
* SPICE INPUT		Tue Jul 31 20:01:38 2018	oai21dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21dm
.subckt oai21dm Y GND VDD C B A
M1 GND B N_2 GND mn15  l=0.13u w=0.36u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.36u m=1
M3 Y C N_2 GND mn15  l=0.13u w=0.36u m=1
M4 N_20 B Y VDD mp15  l=0.13u w=0.55u m=1
M5 N_20 A VDD VDD mp15  l=0.13u w=0.55u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.37u m=1
.ends oai21dm
* SPICE INPUT		Tue Jul 31 20:01:51 2018	oai21md0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21md0
.subckt oai21md0 VDD Y B CN GND A
M1 N_3 CN GND GND mn15  l=0.13u w=0.26u m=1
M2 GND A N_9 GND mn15  l=0.13u w=0.26u m=1
M3 GND B N_9 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_3 N_9 GND mn15  l=0.13u w=0.26u m=1
M5 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_6 B Y VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_3 VDD VDD mp15  l=0.13u w=0.27u m=1
M8 N_3 CN VDD VDD mp15  l=0.13u w=0.4u m=1
.ends oai21md0
* SPICE INPUT		Tue Jul 31 20:02:04 2018	oai21md1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21md1
.subckt oai21md1 Y VDD GND CN B A
M1 GND A N_11 GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M3 Y N_5 N_11 GND mn15  l=0.13u w=0.46u m=1
M4 GND CN N_5 GND mn15  l=0.13u w=0.26u m=1
M5 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 N_7 B Y VDD mp15  l=0.13u w=0.69u m=1
M7 VDD N_5 Y VDD mp15  l=0.13u w=0.46u m=1
M8 VDD CN N_5 VDD mp15  l=0.13u w=0.4u m=1
.ends oai21md1
* SPICE INPUT		Tue Jul 31 20:02:18 2018	oai21md2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21md2
.subckt oai21md2 Y GND VDD CN B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M5 Y N_9 N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_2 N_9 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND CN N_9 GND mn15  l=0.13u w=0.3u m=1
M8 VDD A N_13 VDD mp15  l=0.13u w=0.69u m=1
M9 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M12 Y N_9 VDD VDD mp15  l=0.13u w=0.46u m=1
M13 Y N_9 VDD VDD mp15  l=0.13u w=0.46u m=1
M14 N_9 CN VDD VDD mp15  l=0.13u w=0.43u m=1
.ends oai21md2
* SPICE INPUT		Tue Jul 31 20:02:31 2018	oai21md4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai21md4
.subckt oai21md4 Y GND VDD CN B A
M1 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 N_15 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_3 N_15 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_3 N_15 Y GND mn15  l=0.13u w=0.46u m=1
M8 N_3 N_15 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M10 GND B N_3 GND mn15  l=0.13u w=0.46u m=1
M11 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M12 GND B N_3 GND mn15  l=0.13u w=0.46u m=1
M13 GND CN N_15 GND mn15  l=0.13u w=0.46u m=1
M14 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M15 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M16 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD A N_20 VDD mp15  l=0.13u w=0.69u m=1
M18 Y N_15 VDD VDD mp15  l=0.13u w=0.46u m=1
M19 VDD N_15 Y VDD mp15  l=0.13u w=0.46u m=1
M20 Y N_15 VDD VDD mp15  l=0.13u w=0.46u m=1
M21 Y N_15 VDD VDD mp15  l=0.13u w=0.46u m=1
M22 Y B N_20 VDD mp15  l=0.13u w=0.55u m=1
M23 N_20 B Y VDD mp15  l=0.13u w=0.55u m=1
M24 Y B N_20 VDD mp15  l=0.13u w=0.55u m=1
M25 Y B N_20 VDD mp15  l=0.13u w=0.55u m=1
M26 Y B N_20 VDD mp15  l=0.13u w=0.56u m=1
M27 VDD CN N_15 VDD mp15  l=0.13u w=0.69u m=1
.ends oai21md4
* SPICE INPUT		Tue Jul 31 20:02:44 2018	oai221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d0
.subckt oai221d0 VDD Y GND E C D B A
M1 GND B N_14 GND mn15  l=0.13u w=0.26u m=1
M2 GND A N_14 GND mn15  l=0.13u w=0.26u m=1
M3 N_13 D N_14 GND mn15  l=0.13u w=0.26u m=1
M4 N_14 C N_13 GND mn15  l=0.13u w=0.26u m=1
M5 Y E N_13 GND mn15  l=0.13u w=0.26u m=1
M6 Y B N_8 VDD mp15  l=0.13u w=0.4u m=1
M7 Y D N_7 VDD mp15  l=0.13u w=0.4u m=1
M8 N_7 C VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y E VDD VDD mp15  l=0.13u w=0.27u m=1
.ends oai221d0
* SPICE INPUT		Tue Jul 31 20:02:57 2018	oai221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d1
.subckt oai221d1 GND Y VDD E C D B A
M1 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 Y E N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 C N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_5 D N_2 GND mn15  l=0.13u w=0.46u m=1
M6 Y B N_18 VDD mp15  l=0.13u w=0.69u m=1
M7 N_17 C VDD VDD mp15  l=0.13u w=0.69u m=1
M8 Y D N_17 VDD mp15  l=0.13u w=0.69u m=1
M9 N_18 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 Y E VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oai221d1
* SPICE INPUT		Tue Jul 31 20:03:10 2018	oai221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d2
.subckt oai221d2 Y VDD GND E C D A B
M1 N_20 C N_22 GND mn15  l=0.13u w=0.46u m=1
M2 N_20 D N_22 GND mn15  l=0.13u w=0.46u m=1
M3 N_20 D N_22 GND mn15  l=0.13u w=0.46u m=1
M4 N_20 C N_22 GND mn15  l=0.13u w=0.46u m=1
M5 N_20 E Y GND mn15  l=0.13u w=0.46u m=1
M6 N_20 E Y GND mn15  l=0.13u w=0.46u m=1
M7 GND B N_22 GND mn15  l=0.13u w=0.46u m=1
M8 N_22 B GND GND mn15  l=0.13u w=0.46u m=1
M9 GND A N_22 GND mn15  l=0.13u w=0.46u m=1
M10 N_22 A GND GND mn15  l=0.13u w=0.46u m=1
M11 N_11 C VDD VDD mp15  l=0.13u w=0.595u m=1
M12 N_11 D Y VDD mp15  l=0.13u w=0.595u m=1
M13 Y D N_10 VDD mp15  l=0.13u w=0.595u m=1
M14 N_10 C VDD VDD mp15  l=0.13u w=0.595u m=1
M15 VDD E Y VDD mp15  l=0.13u w=0.46u m=1
M16 VDD E Y VDD mp15  l=0.13u w=0.46u m=1
M17 Y B N_12 VDD mp15  l=0.13u w=0.69u m=1
M18 Y B N_13 VDD mp15  l=0.13u w=0.69u m=1
M19 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends oai221d2
* SPICE INPUT		Tue Jul 31 20:03:23 2018	oai221d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai221d4
.subckt oai221d4 Y D C A B GND VDD E
M1 N_10 C N_11 GND mn15  l=0.13u w=0.46u m=1
M2 N_10 C N_11 GND mn15  l=0.13u w=0.46u m=1
M3 N_10 C N_11 GND mn15  l=0.13u w=0.46u m=1
M4 N_10 D N_11 GND mn15  l=0.13u w=0.46u m=1
M5 N_10 D N_11 GND mn15  l=0.13u w=0.46u m=1
M6 N_10 D N_11 GND mn15  l=0.13u w=0.46u m=1
M7 N_10 D N_11 GND mn15  l=0.13u w=0.46u m=1
M8 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M9 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M10 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M11 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M12 N_10 C N_11 GND mn15  l=0.13u w=0.46u m=1
M13 N_11 B GND GND mn15  l=0.13u w=0.46u m=1
M14 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M15 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M16 GND A N_11 GND mn15  l=0.13u w=0.46u m=1
M17 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M18 GND B N_11 GND mn15  l=0.13u w=0.46u m=1
M19 N_11 A GND GND mn15  l=0.13u w=0.46u m=1
M20 GND A N_11 GND mn15  l=0.13u w=0.46u m=1
M21 N_21 B Y VDD mp15  l=0.13u w=0.69u m=1
M22 N_20 B Y VDD mp15  l=0.13u w=0.69u m=1
M23 N_22 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_22 B Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_23 B Y VDD mp15  l=0.13u w=0.69u m=1
M28 N_24 C VDD VDD mp15  l=0.13u w=0.595u m=1
M29 N_24 D Y VDD mp15  l=0.13u w=0.595u m=1
M30 N_23 A VDD VDD mp15  l=0.13u w=0.69u m=1
M31 N_26 C VDD VDD mp15  l=0.13u w=0.595u m=1
M32 N_25 C VDD VDD mp15  l=0.13u w=0.595u m=1
M33 N_25 D Y VDD mp15  l=0.13u w=0.595u m=1
M34 N_26 D Y VDD mp15  l=0.13u w=0.595u m=1
M35 N_27 D Y VDD mp15  l=0.13u w=0.595u m=1
M36 VDD E Y VDD mp15  l=0.13u w=0.46u m=1
M37 VDD E Y VDD mp15  l=0.13u w=0.46u m=1
M38 Y E VDD VDD mp15  l=0.13u w=0.46u m=1
M39 Y E VDD VDD mp15  l=0.13u w=0.46u m=1
M40 N_27 C VDD VDD mp15  l=0.13u w=0.595u m=1
.ends oai221d4
* SPICE INPUT		Tue Jul 31 20:03:37 2018	oai222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d0
.subckt oai222d0 Y VDD GND F E C D B A
M1 N_14 E Y GND mn15  l=0.13u w=0.26u m=1
M2 N_14 F Y GND mn15  l=0.13u w=0.26u m=1
M3 N_14 C N_16 GND mn15  l=0.13u w=0.26u m=1
M4 GND A N_16 GND mn15  l=0.13u w=0.26u m=1
M5 N_16 B GND GND mn15  l=0.13u w=0.26u m=1
M6 N_16 D N_14 GND mn15  l=0.13u w=0.26u m=1
M7 VDD C N_11 VDD mp15  l=0.13u w=0.4u m=1
M8 VDD E N_9 VDD mp15  l=0.13u w=0.4u m=1
M9 Y F N_9 VDD mp15  l=0.13u w=0.4u m=1
M10 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M11 Y B N_10 VDD mp15  l=0.13u w=0.4u m=1
M12 N_11 D Y VDD mp15  l=0.13u w=0.4u m=1
.ends oai222d0
* SPICE INPUT		Tue Jul 31 20:03:50 2018	oai222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d1
.subckt oai222d1 GND Y VDD E F C D B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 D N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M5 Y E N_3 GND mn15  l=0.13u w=0.46u m=1
M6 Y F N_3 GND mn15  l=0.13u w=0.46u m=1
M7 VDD E N_21 VDD mp15  l=0.13u w=0.69u m=1
M8 Y F N_21 VDD mp15  l=0.13u w=0.69u m=1
M9 N_23 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_23 B Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_24 D Y VDD mp15  l=0.13u w=0.36u m=1
M12 VDD C N_24 VDD mp15  l=0.13u w=0.36u m=1
M13 VDD C N_22 VDD mp15  l=0.13u w=0.35u m=1
M14 Y D N_22 VDD mp15  l=0.13u w=0.35u m=1
.ends oai222d1
* SPICE INPUT		Tue Jul 31 20:04:02 2018	oai222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d2
.subckt oai222d2 Y GND VDD A B D F E C
M1 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M2 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M3 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M4 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_7 C N_3 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 D N_7 GND mn15  l=0.13u w=0.46u m=1
M8 N_3 D N_7 GND mn15  l=0.13u w=0.46u m=1
M9 N_7 B GND GND mn15  l=0.13u w=0.46u m=1
M10 GND A N_7 GND mn15  l=0.13u w=0.46u m=1
M11 N_7 A GND GND mn15  l=0.13u w=0.46u m=1
M12 N_7 B GND GND mn15  l=0.13u w=0.46u m=1
M13 N_21 E VDD VDD mp15  l=0.13u w=0.46u m=1
M14 N_21 E VDD VDD mp15  l=0.13u w=0.46u m=1
M15 N_21 E VDD VDD mp15  l=0.13u w=0.46u m=1
M16 N_20 C VDD VDD mp15  l=0.13u w=0.46u m=1
M17 VDD C N_20 VDD mp15  l=0.13u w=0.46u m=1
M18 N_20 C VDD VDD mp15  l=0.13u w=0.46u m=1
M19 N_20 D Y VDD mp15  l=0.13u w=0.46u m=1
M20 N_20 D Y VDD mp15  l=0.13u w=0.46u m=1
M21 N_20 D Y VDD mp15  l=0.13u w=0.46u m=1
M22 N_28 B Y VDD mp15  l=0.13u w=0.69u m=1
M23 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_27 B Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_21 F Y VDD mp15  l=0.13u w=0.46u m=1
M27 Y F N_21 VDD mp15  l=0.13u w=0.46u m=1
M28 Y F N_21 VDD mp15  l=0.13u w=0.46u m=1
.ends oai222d2
* SPICE INPUT		Tue Jul 31 20:04:15 2018	oai222d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai222d4
.subckt oai222d4 GND Y F C VDD E A D B
M1 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M4 N_2 C N_3 GND mn15  l=0.13u w=0.46u m=1
M5 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M7 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M8 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M9 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M10 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M11 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M12 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M13 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M14 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M15 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M16 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M17 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M18 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M19 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M20 N_3 F Y GND mn15  l=0.13u w=0.46u m=1
M21 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M22 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M23 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M24 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M25 N_37 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD A N_37 VDD mp15  l=0.13u w=0.69u m=1
M27 N_37 A VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD A N_37 VDD mp15  l=0.13u w=0.69u m=1
M29 N_37 B Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y B N_37 VDD mp15  l=0.13u w=0.69u m=1
M31 N_37 B Y VDD mp15  l=0.13u w=0.69u m=1
M32 N_37 B Y VDD mp15  l=0.13u w=0.69u m=1
M33 Y F N_31 VDD mp15  l=0.13u w=0.565u m=1
M34 Y F N_31 VDD mp15  l=0.13u w=0.565u m=1
M35 Y F N_31 VDD mp15  l=0.13u w=0.565u m=1
M36 N_31 F Y VDD mp15  l=0.13u w=0.565u m=1
M37 Y F N_31 VDD mp15  l=0.13u w=0.5u m=1
M38 VDD C N_33 VDD mp15  l=0.13u w=0.56u m=1
M39 N_33 C VDD VDD mp15  l=0.13u w=0.55u m=1
M40 N_33 C VDD VDD mp15  l=0.13u w=0.55u m=1
M41 VDD C N_33 VDD mp15  l=0.13u w=0.55u m=1
M42 N_33 C VDD VDD mp15  l=0.13u w=0.55u m=1
M43 Y D N_33 VDD mp15  l=0.13u w=0.565u m=1
M44 Y D N_33 VDD mp15  l=0.13u w=0.565u m=1
M45 Y D N_33 VDD mp15  l=0.13u w=0.565u m=1
M46 N_33 D Y VDD mp15  l=0.13u w=0.565u m=1
M47 N_33 D Y VDD mp15  l=0.13u w=0.5u m=1
M48 N_31 E VDD VDD mp15  l=0.13u w=0.56u m=1
M49 VDD E N_31 VDD mp15  l=0.13u w=0.55u m=1
M50 N_31 E VDD VDD mp15  l=0.13u w=0.55u m=1
M51 N_31 E VDD VDD mp15  l=0.13u w=0.55u m=1
M52 N_31 E VDD VDD mp15  l=0.13u w=0.55u m=1
.ends oai222d4
* SPICE INPUT		Tue Jul 31 20:04:28 2018	oai22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d0
.subckt oai22d0 VDD Y GND A C B D
M1 N_12 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_12 D Y GND mn15  l=0.13u w=0.26u m=1
M3 N_12 B GND GND mn15  l=0.13u w=0.26u m=1
M4 N_12 C Y GND mn15  l=0.13u w=0.26u m=1
M5 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y D N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 Y B N_8 VDD mp15  l=0.13u w=0.4u m=1
M8 VDD C N_7 VDD mp15  l=0.13u w=0.4u m=1
.ends oai22d0
* SPICE INPUT		Tue Jul 31 20:04:41 2018	oai22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d1
.subckt oai22d1 VDD Y GND A C B D
M1 N_12 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_12 D Y GND mn15  l=0.13u w=0.46u m=1
M3 N_12 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_12 C Y GND mn15  l=0.13u w=0.46u m=1
M5 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y D N_7 VDD mp15  l=0.13u w=0.595u m=1
M7 N_8 B Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD C N_7 VDD mp15  l=0.13u w=0.595u m=1
.ends oai22d1
* SPICE INPUT		Tue Jul 31 20:04:54 2018	oai22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d2
.subckt oai22d2 VDD Y GND D A B C
M1 GND B N_20 GND mn15  l=0.13u w=0.46u m=1
M2 N_20 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M5 N_20 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_20 C Y GND mn15  l=0.13u w=0.46u m=1
M7 N_20 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_20 D Y GND mn15  l=0.13u w=0.46u m=1
M9 N_9 B Y VDD mp15  l=0.13u w=0.69u m=1
M10 Y B N_8 VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 VDD C N_7 VDD mp15  l=0.13u w=0.595u m=1
M13 N_9 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_10 C VDD VDD mp15  l=0.13u w=0.595u m=1
M15 Y D N_7 VDD mp15  l=0.13u w=0.595u m=1
M16 Y D N_10 VDD mp15  l=0.13u w=0.595u m=1
.ends oai22d2
* SPICE INPUT		Tue Jul 31 20:05:07 2018	oai22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22d4
.subckt oai22d4 VDD Y A B D GND C
M1 GND B N_30 GND mn15  l=0.13u w=0.46u m=1
M2 N_30 B GND GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_30 GND mn15  l=0.13u w=0.46u m=1
M4 N_30 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_30 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_30 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_30 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_30 C Y GND mn15  l=0.13u w=0.46u m=1
M9 N_30 A GND GND mn15  l=0.13u w=0.46u m=1
M10 N_30 C Y GND mn15  l=0.13u w=0.46u m=1
M11 N_30 D Y GND mn15  l=0.13u w=0.46u m=1
M12 N_30 D Y GND mn15  l=0.13u w=0.46u m=1
M13 N_30 C Y GND mn15  l=0.13u w=0.46u m=1
M14 N_30 C Y GND mn15  l=0.13u w=0.46u m=1
M15 N_30 D Y GND mn15  l=0.13u w=0.46u m=1
M16 N_30 D Y GND mn15  l=0.13u w=0.46u m=1
M17 N_15 B Y VDD mp15  l=0.13u w=0.69u m=1
M18 Y B N_14 VDD mp15  l=0.13u w=0.69u m=1
M19 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_13 B Y VDD mp15  l=0.13u w=0.69u m=1
M21 Y B N_12 VDD mp15  l=0.13u w=0.69u m=1
M22 N_14 A VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_13 A VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_16 C VDD VDD mp15  l=0.13u w=0.595u m=1
M25 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD C N_11 VDD mp15  l=0.13u w=0.595u m=1
M27 Y D N_11 VDD mp15  l=0.13u w=0.595u m=1
M28 Y D N_18 VDD mp15  l=0.13u w=0.595u m=1
M29 N_18 C VDD VDD mp15  l=0.13u w=0.595u m=1
M30 N_17 C VDD VDD mp15  l=0.13u w=0.595u m=1
M31 N_17 D Y VDD mp15  l=0.13u w=0.595u m=1
M32 Y D N_16 VDD mp15  l=0.13u w=0.595u m=1
.ends oai22d4
* SPICE INPUT		Tue Jul 31 20:05:20 2018	oai22dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai22dm
.subckt oai22dm VDD Y GND A C B D
M1 N_12 A GND GND mn15  l=0.13u w=0.36u m=1
M2 N_12 D Y GND mn15  l=0.13u w=0.36u m=1
M3 N_12 B GND GND mn15  l=0.13u w=0.36u m=1
M4 N_12 C Y GND mn15  l=0.13u w=0.36u m=1
M5 N_8 A VDD VDD mp15  l=0.13u w=0.55u m=1
M6 Y D N_7 VDD mp15  l=0.13u w=0.55u m=1
M7 Y B N_8 VDD mp15  l=0.13u w=0.55u m=1
M8 VDD C N_7 VDD mp15  l=0.13u w=0.55u m=1
.ends oai22dm
* SPICE INPUT		Tue Jul 31 20:05:32 2018	oai2m1d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai2m1d0
.subckt oai2m1d0 VDD Y GND C A BN
M1 Y C N_11 GND mn15  l=0.13u w=0.26u m=1
M2 N_11 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 GND A N_11 GND mn15  l=0.13u w=0.26u m=1
M4 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M5 N_3 BN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.27u m=1
M7 N_7 N_3 Y VDD mp15  l=0.13u w=0.4u m=1
M8 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends oai2m1d0
* SPICE INPUT		Tue Jul 31 20:05:45 2018	oai2m1d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai2m1d1
.subckt oai2m1d1 GND Y VDD C A BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.26u m=1
M2 Y C N_4 GND mn15  l=0.13u w=0.46u m=1
M3 N_4 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_4 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 BN VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M7 N_26 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M8 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends oai2m1d1
* SPICE INPUT		Tue Jul 31 20:05:57 2018	oai2m1d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai2m1d2
.subckt oai2m1d2 GND Y VDD C A BN
M1 N_3 BN GND GND mn15  l=0.13u w=0.46u m=1
M2 N_5 C Y GND mn15  l=0.13u w=0.46u m=1
M3 N_5 C Y GND mn15  l=0.13u w=0.46u m=1
M4 N_5 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_5 N_3 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_3 BN VDD VDD mp15  l=0.13u w=0.69u m=1
M9 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M10 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M11 N_39 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M12 N_39 A VDD VDD mp15  l=0.13u w=0.69u m=1
M13 N_38 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_38 N_3 Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai2m1d2
* SPICE INPUT		Tue Jul 31 20:06:10 2018	oai2m1d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai2m1d4
.subckt oai2m1d4 GND Y VDD C A BN
M1 GND BN N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND BN N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M6 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M7 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M8 N_6 C Y GND mn15  l=0.13u w=0.46u m=1
M9 N_6 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_6 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_6 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M13 N_6 A GND GND mn15  l=0.13u w=0.46u m=1
M14 N_6 N_2 GND GND mn15  l=0.13u w=0.46u m=1
M15 VDD BN N_2 VDD mp15  l=0.13u w=0.69u m=1
M16 VDD BN N_2 VDD mp15  l=0.13u w=0.69u m=1
M17 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_29 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M20 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M21 Y C VDD VDD mp15  l=0.13u w=0.48u m=1
M22 VDD C Y VDD mp15  l=0.13u w=0.48u m=1
M23 N_29 N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M24 N_28 N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M25 N_27 N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M26 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M28 N_26 N_2 Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai2m1d4
* SPICE INPUT		Tue Jul 31 20:06:23 2018	oai31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d0
.subckt oai31d0 VDD Y GND D A B C
M1 N_11 C GND GND mn15  l=0.13u w=0.26u m=1
M2 N_11 B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y D N_11 GND mn15  l=0.13u w=0.26u m=1
M4 GND A N_11 GND mn15  l=0.13u w=0.26u m=1
M5 N_7 C Y VDD mp15  l=0.13u w=0.4u m=1
M6 N_8 B N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 Y D VDD VDD mp15  l=0.13u w=0.27u m=1
M8 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends oai31d0
* SPICE INPUT		Tue Jul 31 20:06:36 2018	oai31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d1
.subckt oai31d1 Y GND VDD D A B C
M1 Y D N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 C GND GND mn15  l=0.13u w=0.46u m=1
M5 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M6 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_15 B N_14 VDD mp15  l=0.13u w=0.69u m=1
M8 N_14 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai31d1
* SPICE INPUT		Tue Jul 31 20:06:50 2018	oai31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d2
.subckt oai31d2 Y VDD GND D A B C
M1 GND A N_17 GND mn15  l=0.13u w=0.46u m=1
M2 N_17 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_17 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_17 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_17 D Y GND mn15  l=0.13u w=0.46u m=1
M7 N_17 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_17 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_9 B N_8 VDD mp15  l=0.13u w=0.69u m=1
M11 N_9 C Y VDD mp15  l=0.13u w=0.69u m=1
M12 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
M13 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD D Y VDD mp15  l=0.13u w=0.46u m=1
M15 VDD D Y VDD mp15  l=0.13u w=0.46u m=1
M16 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends oai31d2
* SPICE INPUT		Tue Jul 31 20:07:03 2018	oai31d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai31d4
.subckt oai31d4 GND VDD Y D C B A
M1 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M2 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M3 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M4 N_9 D Y GND mn15  l=0.13u w=0.46u m=1
M5 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_9 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_9 B GND GND mn15  l=0.13u w=0.46u m=1
M10 N_9 B GND GND mn15  l=0.13u w=0.46u m=1
M11 N_9 B GND GND mn15  l=0.13u w=0.46u m=1
M12 N_9 B GND GND mn15  l=0.13u w=0.46u m=1
M13 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M14 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M15 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M16 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M17 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 VDD A N_11 VDD mp15  l=0.13u w=0.69u m=1
M19 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_11 VDD mp15  l=0.13u w=0.69u m=1
M21 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M22 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M23 N_11 B N_10 VDD mp15  l=0.13u w=0.69u m=1
M24 N_10 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M25 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M26 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M27 Y D VDD VDD mp15  l=0.13u w=0.46u m=1
M28 VDD D Y VDD mp15  l=0.13u w=0.46u m=1
M29 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
M30 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
M31 Y C N_10 VDD mp15  l=0.13u w=0.69u m=1
M32 N_10 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai31d4
* SPICE INPUT		Tue Jul 31 20:07:16 2018	oai32d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d0
.subckt oai32d0 Y VDD GND E D A B C
M1 N_12 D Y GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_12 GND mn15  l=0.13u w=0.26u m=1
M3 N_12 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_12 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y E N_12 GND mn15  l=0.13u w=0.26u m=1
M6 VDD D N_8 VDD mp15  l=0.13u w=0.4u m=1
M7 N_10 B N_9 VDD mp15  l=0.13u w=0.4u m=1
M8 N_9 C Y VDD mp15  l=0.13u w=0.4u m=1
M9 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 Y E N_8 VDD mp15  l=0.13u w=0.4u m=1
.ends oai32d0
* SPICE INPUT		Tue Jul 31 20:07:29 2018	oai32d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d1
.subckt oai32d1 Y GND VDD D E A B C
M1 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M2 N_3 D Y GND mn15  l=0.13u w=0.46u m=1
M3 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_14 D VDD VDD mp15  l=0.13u w=0.345u m=1
M7 Y E N_14 VDD mp15  l=0.13u w=0.345u m=1
M8 Y E N_17 VDD mp15  l=0.13u w=0.345u m=1
M9 N_17 D VDD VDD mp15  l=0.13u w=0.345u m=1
M10 N_16 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_16 B N_15 VDD mp15  l=0.13u w=0.69u m=1
M12 N_15 C Y VDD mp15  l=0.13u w=0.69u m=1
.ends oai32d1
* SPICE INPUT		Tue Jul 31 20:07:42 2018	oai32d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d2
.subckt oai32d2 Y GND VDD E D A B C
M1 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 D Y GND mn15  l=0.13u w=0.46u m=1
M6 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M7 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_3 D Y GND mn15  l=0.13u w=0.46u m=1
M9 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M10 N_3 E Y GND mn15  l=0.13u w=0.46u m=1
M11 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_27 B N_26 VDD mp15  l=0.13u w=0.69u m=1
M13 N_27 C Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_29 C Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD D N_28 VDD mp15  l=0.13u w=0.455u m=1
M16 N_32 D VDD VDD mp15  l=0.13u w=0.455u m=1
M17 N_30 B N_29 VDD mp15  l=0.13u w=0.69u m=1
M18 Y E N_28 VDD mp15  l=0.13u w=0.455u m=1
M19 N_30 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_31 D VDD VDD mp15  l=0.13u w=0.455u m=1
M21 N_32 E Y VDD mp15  l=0.13u w=0.455u m=1
M22 Y E N_31 VDD mp15  l=0.13u w=0.455u m=1
.ends oai32d2
* SPICE INPUT		Tue Jul 31 20:07:55 2018	oai32d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai32d4
.subckt oai32d4 D GND VDD Y E C B A
M1 N_10 B GND GND mn15  l=0.13u w=0.46u m=1
M2 N_10 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_10 B GND GND mn15  l=0.13u w=0.46u m=1
M4 GND B N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M6 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M7 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M8 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M9 N_10 D Y GND mn15  l=0.13u w=0.46u m=1
M10 N_10 C GND GND mn15  l=0.13u w=0.46u m=1
M11 N_10 C GND GND mn15  l=0.13u w=0.46u m=1
M12 N_10 C GND GND mn15  l=0.13u w=0.46u m=1
M13 GND C N_10 GND mn15  l=0.13u w=0.46u m=1
M14 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M15 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M16 N_10 E Y GND mn15  l=0.13u w=0.46u m=1
M17 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M18 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M19 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M20 N_10 A GND GND mn15  l=0.13u w=0.46u m=1
M21 N_12 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M22 N_12 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M23 N_12 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M24 N_11 B N_12 VDD mp15  l=0.13u w=0.69u m=1
M25 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M27 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M29 N_37 D VDD VDD mp15  l=0.13u w=0.47u m=1
M30 N_38 E Y VDD mp15  l=0.13u w=0.47u m=1
M31 N_39 D VDD VDD mp15  l=0.13u w=0.47u m=1
M32 VDD D N_38 VDD mp15  l=0.13u w=0.47u m=1
M33 N_41 D VDD VDD mp15  l=0.13u w=0.47u m=1
M34 VDD D N_40 VDD mp15  l=0.13u w=0.47u m=1
M35 N_11 C Y VDD mp15  l=0.13u w=0.69u m=1
M36 N_11 C Y VDD mp15  l=0.13u w=0.69u m=1
M37 Y C N_11 VDD mp15  l=0.13u w=0.69u m=1
M38 N_11 C Y VDD mp15  l=0.13u w=0.69u m=1
M39 N_40 E Y VDD mp15  l=0.13u w=0.47u m=1
M40 Y E N_39 VDD mp15  l=0.13u w=0.47u m=1
M41 Y E N_37 VDD mp15  l=0.13u w=0.47u m=1
M42 Y E N_41 VDD mp15  l=0.13u w=0.47u m=1
.ends oai32d4
* SPICE INPUT		Tue Jul 31 20:08:09 2018	oai33d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d0
.subckt oai33d0 VDD Y GND D E F C B A
M1 Y D N_15 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_15 GND mn15  l=0.13u w=0.26u m=1
M3 Y E N_15 GND mn15  l=0.13u w=0.26u m=1
M4 N_15 F Y GND mn15  l=0.13u w=0.26u m=1
M5 N_15 C GND GND mn15  l=0.13u w=0.26u m=1
M6 N_15 A GND GND mn15  l=0.13u w=0.26u m=1
M7 VDD D N_9 VDD mp15  l=0.13u w=0.4u m=1
M8 N_11 B N_10 VDD mp15  l=0.13u w=0.4u m=1
M9 N_12 E N_9 VDD mp15  l=0.13u w=0.4u m=1
M10 N_12 F Y VDD mp15  l=0.13u w=0.4u m=1
M11 Y C N_11 VDD mp15  l=0.13u w=0.4u m=1
M12 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends oai33d0
* SPICE INPUT		Tue Jul 31 20:08:22 2018	oai33d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d1
.subckt oai33d1 Y GND VDD D E F C B A
M1 GND C N_2 GND mn15  l=0.13u w=0.46u m=1
M2 Y F N_2 GND mn15  l=0.13u w=0.46u m=1
M3 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M5 Y D N_2 GND mn15  l=0.13u w=0.46u m=1
M6 Y E N_2 GND mn15  l=0.13u w=0.46u m=1
M7 Y C N_42 VDD mp15  l=0.13u w=0.69u m=1
M8 Y F N_13 VDD mp15  l=0.13u w=0.69u m=1
M9 N_42 B N_41 VDD mp15  l=0.13u w=0.69u m=1
M10 N_41 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_13 E N_12 VDD mp15  l=0.13u w=0.35u m=1
M12 N_12 E N_13 VDD mp15  l=0.13u w=0.34u m=1
M13 VDD D N_12 VDD mp15  l=0.13u w=0.69u m=1
.ends oai33d1
* SPICE INPUT		Tue Jul 31 20:08:35 2018	oai33d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d2
.subckt oai33d2 Y GND VDD E F D B C A
M1 GND A N_3 GND mn15  l=0.13u w=0.35u m=1
M2 GND B N_3 GND mn15  l=0.13u w=0.34u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.35u m=1
M4 N_3 A GND GND mn15  l=0.13u w=0.34u m=1
M5 N_3 C GND GND mn15  l=0.13u w=0.35u m=1
M6 N_3 C GND GND mn15  l=0.13u w=0.34u m=1
M7 N_3 E Y GND mn15  l=0.13u w=0.35u m=1
M8 N_3 E Y GND mn15  l=0.13u w=0.34u m=1
M9 N_3 D Y GND mn15  l=0.13u w=0.34u m=1
M10 N_3 D Y GND mn15  l=0.13u w=0.35u m=1
M11 N_3 F Y GND mn15  l=0.13u w=0.34u m=1
M12 N_3 F Y GND mn15  l=0.13u w=0.35u m=1
M13 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_15 B N_27 VDD mp15  l=0.13u w=0.69u m=1
M15 N_15 B N_28 VDD mp15  l=0.13u w=0.69u m=1
M16 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_15 C Y VDD mp15  l=0.13u w=0.69u m=1
M18 N_15 C Y VDD mp15  l=0.13u w=0.69u m=1
M19 N_23 E N_20 VDD mp15  l=0.13u w=0.46u m=1
M20 N_20 E N_23 VDD mp15  l=0.13u w=0.46u m=1
M21 N_23 E N_20 VDD mp15  l=0.13u w=0.46u m=1
M22 N_23 D VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_23 D VDD VDD mp15  l=0.13u w=0.69u m=1
M24 N_20 F Y VDD mp15  l=0.13u w=0.46u m=1
M25 N_20 F Y VDD mp15  l=0.13u w=0.46u m=1
M26 Y F N_20 VDD mp15  l=0.13u w=0.46u m=1
.ends oai33d2
* SPICE INPUT		Tue Jul 31 20:08:48 2018	oai33d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oai33d4
.subckt oai33d4 GND F Y D C E VDD B A
M1 N_14 F Y GND mn15  l=0.13u w=0.56u m=1
M2 Y F N_14 GND mn15  l=0.13u w=0.56u m=1
M3 Y F N_14 GND mn15  l=0.13u w=0.56u m=1
M4 Y F N_14 GND mn15  l=0.13u w=0.16u m=1
M5 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M6 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M7 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M8 N_14 A GND GND mn15  l=0.13u w=0.46u m=1
M9 N_14 B GND GND mn15  l=0.13u w=0.46u m=1
M10 N_14 B GND GND mn15  l=0.13u w=0.46u m=1
M11 N_14 B GND GND mn15  l=0.13u w=0.46u m=1
M12 N_14 B GND GND mn15  l=0.13u w=0.46u m=1
M13 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M14 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M15 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M16 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M17 N_14 E Y GND mn15  l=0.13u w=0.46u m=1
M18 N_14 E Y GND mn15  l=0.13u w=0.46u m=1
M19 N_14 E Y GND mn15  l=0.13u w=0.46u m=1
M20 Y E N_14 GND mn15  l=0.13u w=0.46u m=1
M21 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M22 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M23 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M24 N_14 D Y GND mn15  l=0.13u w=0.46u m=1
M25 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M27 N_12 A VDD VDD mp15  l=0.13u w=0.69u m=1
M28 VDD A N_12 VDD mp15  l=0.13u w=0.69u m=1
M29 N_13 B N_12 VDD mp15  l=0.13u w=0.69u m=1
M30 N_12 B N_13 VDD mp15  l=0.13u w=0.69u m=1
M31 N_12 B N_13 VDD mp15  l=0.13u w=0.69u m=1
M32 N_12 B N_13 VDD mp15  l=0.13u w=0.69u m=1
M33 Y F N_15 VDD mp15  l=0.13u w=0.6u m=1
M34 Y F N_15 VDD mp15  l=0.13u w=0.6u m=1
M35 Y F N_15 VDD mp15  l=0.13u w=0.6u m=1
M36 N_15 F Y VDD mp15  l=0.13u w=0.6u m=1
M37 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
M38 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
M39 Y C N_13 VDD mp15  l=0.13u w=0.69u m=1
M40 N_13 C Y VDD mp15  l=0.13u w=0.69u m=1
M41 N_11 E N_15 VDD mp15  l=0.13u w=0.6u m=1
M42 N_15 E N_11 VDD mp15  l=0.13u w=0.6u m=1
M43 N_11 E N_15 VDD mp15  l=0.13u w=0.6u m=1
M44 N_15 E N_11 VDD mp15  l=0.13u w=0.6u m=1
M45 N_11 D VDD VDD mp15  l=0.13u w=0.6u m=1
M46 N_11 D VDD VDD mp15  l=0.13u w=0.6u m=1
M47 N_11 D VDD VDD mp15  l=0.13u w=0.6u m=1
M48 VDD D N_11 VDD mp15  l=0.13u w=0.6u m=1
.ends oai33d4
* SPICE INPUT		Tue Jul 31 20:09:01 2018	oaim21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d0
.subckt oaim21d0 Y GND VDD C AN BN
M1 N_6 BN N_3 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 N_5 GND mn15  l=0.13u w=0.26u m=1
M3 GND C N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 AN GND GND mn15  l=0.13u w=0.26u m=1
M5 N_3 BN VDD VDD mp15  l=0.13u w=0.35u m=1
M6 Y N_3 VDD VDD mp15  l=0.13u w=0.35u m=1
M7 VDD C Y VDD mp15  l=0.13u w=0.35u m=1
M8 N_3 AN VDD VDD mp15  l=0.13u w=0.35u m=1
.ends oaim21d0
* SPICE INPUT		Tue Jul 31 20:09:14 2018	oaim21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d1
.subckt oaim21d1 Y GND VDD C AN BN
M1 Y N_3 N_5 GND mn15  l=0.13u w=0.46u m=1
M2 GND C N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 AN GND GND mn15  l=0.13u w=0.29u m=1
M4 N_6 BN N_3 GND mn15  l=0.13u w=0.29u m=1
M5 VDD N_3 Y VDD mp15  l=0.13u w=0.61u m=1
M6 VDD C Y VDD mp15  l=0.13u w=0.61u m=1
M7 N_3 AN VDD VDD mp15  l=0.13u w=0.35u m=1
M8 N_3 BN VDD VDD mp15  l=0.13u w=0.35u m=1
.ends oaim21d1
* SPICE INPUT		Tue Jul 31 20:09:27 2018	oaim21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d2
.subckt oaim21d2 GND Y VDD C AN BN
M1 Y N_3 N_6 GND mn15  l=0.13u w=0.46u m=1
M2 Y N_3 N_8 GND mn15  l=0.13u w=0.46u m=1
M3 N_6 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_8 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_7 AN GND GND mn15  l=0.13u w=0.37u m=1
M6 N_7 BN N_3 GND mn15  l=0.13u w=0.37u m=1
M7 VDD N_3 Y VDD mp15  l=0.13u w=0.61u m=1
M8 VDD N_3 Y VDD mp15  l=0.13u w=0.61u m=1
M9 VDD C Y VDD mp15  l=0.13u w=0.61u m=1
M10 Y C VDD VDD mp15  l=0.13u w=0.61u m=1
M11 VDD AN N_3 VDD mp15  l=0.13u w=0.46u m=1
M12 N_3 BN VDD VDD mp15  l=0.13u w=0.46u m=1
.ends oaim21d2
* SPICE INPUT		Tue Jul 31 20:09:40 2018	oaim21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21d4
.subckt oaim21d4 GND Y C VDD AN BN
M1 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 C GND GND mn15  l=0.13u w=0.46u m=1
M3 N_13 N_4 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_4 N_12 GND mn15  l=0.13u w=0.46u m=1
M5 N_12 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_11 AN GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_4 N_9 GND mn15  l=0.13u w=0.46u m=1
M8 Y N_4 N_14 GND mn15  l=0.13u w=0.46u m=1
M9 N_11 BN N_4 GND mn15  l=0.13u w=0.46u m=1
M10 N_4 BN N_10 GND mn15  l=0.13u w=0.46u m=1
M11 N_9 C GND GND mn15  l=0.13u w=0.46u m=1
M12 N_10 AN GND GND mn15  l=0.13u w=0.46u m=1
M13 Y C VDD VDD mp15  l=0.13u w=0.61u m=1
M14 Y C VDD VDD mp15  l=0.13u w=0.61u m=1
M15 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M16 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M17 Y C VDD VDD mp15  l=0.13u w=0.61u m=1
M18 VDD AN N_4 VDD mp15  l=0.13u w=0.57u m=1
M19 VDD N_4 Y VDD mp15  l=0.13u w=0.61u m=1
M20 Y N_4 VDD VDD mp15  l=0.13u w=0.61u m=1
M21 N_4 BN VDD VDD mp15  l=0.13u w=0.57u m=1
M22 N_4 BN VDD VDD mp15  l=0.13u w=0.57u m=1
M23 VDD C Y VDD mp15  l=0.13u w=0.61u m=1
M24 N_4 AN VDD VDD mp15  l=0.13u w=0.57u m=1
.ends oaim21d4
* SPICE INPUT		Tue Jul 31 20:09:53 2018	oaim21dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim21dm
.subckt oaim21dm Y GND VDD C AN BN
M1 Y N_3 N_5 GND mn15  l=0.13u w=0.36u m=1
M2 N_6 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 N_6 BN N_3 GND mn15  l=0.13u w=0.26u m=1
M4 GND C N_5 GND mn15  l=0.13u w=0.36u m=1
M5 VDD N_3 Y VDD mp15  l=0.13u w=0.45u m=1
M6 N_3 AN VDD VDD mp15  l=0.13u w=0.35u m=1
M7 N_3 BN VDD VDD mp15  l=0.13u w=0.35u m=1
M8 VDD C Y VDD mp15  l=0.13u w=0.45u m=1
.ends oaim21dm
* SPICE INPUT		Tue Jul 31 20:10:06 2018	oaim22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d0
.subckt oaim22d0 VDD Y GND D C AN BN
M1 Y N_6 N_10 GND mn15  l=0.13u w=0.26u m=1
M2 N_15 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 N_10 D GND GND mn15  l=0.13u w=0.26u m=1
M4 GND C N_10 GND mn15  l=0.13u w=0.26u m=1
M5 N_15 BN N_6 GND mn15  l=0.13u w=0.26u m=1
M6 N_6 AN VDD VDD mp15  l=0.13u w=0.35u m=1
M7 Y N_6 VDD VDD mp15  l=0.13u w=0.27u m=1
M8 N_7 D Y VDD mp15  l=0.13u w=0.4u m=1
M9 N_7 C VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_6 BN VDD VDD mp15  l=0.13u w=0.35u m=1
.ends oaim22d0
* SPICE INPUT		Tue Jul 31 20:10:19 2018	oaim22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d1
.subckt oaim22d1 VDD Y GND D C AN BN
M1 Y N_6 N_10 GND mn15  l=0.13u w=0.46u m=1
M2 N_15 AN GND GND mn15  l=0.13u w=0.29u m=1
M3 N_10 D GND GND mn15  l=0.13u w=0.46u m=1
M4 GND C N_10 GND mn15  l=0.13u w=0.46u m=1
M5 N_15 BN N_6 GND mn15  l=0.13u w=0.29u m=1
M6 N_6 AN VDD VDD mp15  l=0.13u w=0.37u m=1
M7 Y N_6 VDD VDD mp15  l=0.13u w=0.48u m=1
M8 N_7 D Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_7 C VDD VDD mp15  l=0.13u w=0.69u m=1
M10 N_6 BN VDD VDD mp15  l=0.13u w=0.37u m=1
.ends oaim22d1
* SPICE INPUT		Tue Jul 31 20:10:32 2018	oaim22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d2
.subckt oaim22d2 VDD Y GND C D BN AN
M1 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M2 N_14 D GND GND mn15  l=0.13u w=0.46u m=1
M3 N_14 D GND GND mn15  l=0.13u w=0.46u m=1
M4 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_14 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_14 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_5 BN N_19 GND mn15  l=0.13u w=0.46u m=1
M8 GND AN N_19 GND mn15  l=0.13u w=0.46u m=1
M9 VDD C N_9 VDD mp15  l=0.13u w=0.69u m=1
M10 Y D N_9 VDD mp15  l=0.13u w=0.69u m=1
M11 Y D N_10 VDD mp15  l=0.13u w=0.69u m=1
M12 N_10 C VDD VDD mp15  l=0.13u w=0.69u m=1
M13 Y N_5 VDD VDD mp15  l=0.13u w=0.47u m=1
M14 Y N_5 VDD VDD mp15  l=0.13u w=0.46u m=1
M15 N_5 BN VDD VDD mp15  l=0.13u w=0.6u m=1
M16 N_5 AN VDD VDD mp15  l=0.13u w=0.6u m=1
.ends oaim22d2
* SPICE INPUT		Tue Jul 31 20:10:45 2018	oaim22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22d4
.subckt oaim22d4 VDD Y AN BN D GND C
M1 N_27 D GND GND mn15  l=0.13u w=0.46u m=1
M2 N_27 D GND GND mn15  l=0.13u w=0.46u m=1
M3 N_27 C GND GND mn15  l=0.13u w=0.46u m=1
M4 N_27 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M5 N_27 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_27 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_27 N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 N_27 C GND GND mn15  l=0.13u w=0.46u m=1
M9 N_27 C GND GND mn15  l=0.13u w=0.46u m=1
M10 N_27 D GND GND mn15  l=0.13u w=0.46u m=1
M11 N_27 D GND GND mn15  l=0.13u w=0.46u m=1
M12 N_27 C GND GND mn15  l=0.13u w=0.46u m=1
M13 N_5 BN N_29 GND mn15  l=0.13u w=0.46u m=1
M14 N_5 BN N_30 GND mn15  l=0.13u w=0.46u m=1
M15 N_30 AN GND GND mn15  l=0.13u w=0.46u m=1
M16 GND AN N_29 GND mn15  l=0.13u w=0.46u m=1
M17 N_5 BN VDD VDD mp15  l=0.13u w=0.55u m=1
M18 N_5 BN VDD VDD mp15  l=0.13u w=0.55u m=1
M19 N_5 AN VDD VDD mp15  l=0.13u w=0.55u m=1
M20 N_17 D Y VDD mp15  l=0.13u w=0.69u m=1
M21 Y D N_16 VDD mp15  l=0.13u w=0.69u m=1
M22 N_16 C VDD VDD mp15  l=0.13u w=0.69u m=1
M23 Y N_5 VDD VDD mp15  l=0.13u w=0.46u m=1
M24 Y N_5 VDD VDD mp15  l=0.13u w=0.46u m=1
M25 VDD N_5 Y VDD mp15  l=0.13u w=0.46u m=1
M26 Y N_5 VDD VDD mp15  l=0.13u w=0.46u m=1
M27 N_5 AN VDD VDD mp15  l=0.13u w=0.55u m=1
M28 N_18 C VDD VDD mp15  l=0.13u w=0.69u m=1
M29 N_17 C VDD VDD mp15  l=0.13u w=0.69u m=1
M30 Y D N_15 VDD mp15  l=0.13u w=0.69u m=1
M31 Y D N_18 VDD mp15  l=0.13u w=0.69u m=1
M32 VDD C N_15 VDD mp15  l=0.13u w=0.69u m=1
.ends oaim22d4
* SPICE INPUT		Tue Jul 31 20:10:58 2018	oaim22dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=oaim22dm
.subckt oaim22dm VDD Y GND D C AN BN
M1 GND C N_10 GND mn15  l=0.13u w=0.36u m=1
M2 N_15 AN GND GND mn15  l=0.13u w=0.26u m=1
M3 N_15 BN N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_10 D GND GND mn15  l=0.13u w=0.36u m=1
M5 Y N_6 N_10 GND mn15  l=0.13u w=0.36u m=1
M6 Y N_6 VDD VDD mp15  l=0.13u w=0.38u m=1
M7 N_7 C VDD VDD mp15  l=0.13u w=0.55u m=1
M8 N_6 AN VDD VDD mp15  l=0.13u w=0.35u m=1
M9 N_6 BN VDD VDD mp15  l=0.13u w=0.35u m=1
M10 N_7 D Y VDD mp15  l=0.13u w=0.55u m=1
.ends oaim22dm
* SPICE INPUT		Tue Jul 31 20:11:11 2018	or02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d0
.subckt or02d0 VDD Y GND A B
M1 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_5 B N_4 VDD mp15  l=0.13u w=0.4u m=1
M5 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends or02d0
* SPICE INPUT		Tue Jul 31 20:11:24 2018	or02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d1
.subckt or02d1 VDD Y GND A B
M1 N_4 B GND GND mn15  l=0.13u w=0.29u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.29u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 B N_4 VDD mp15  l=0.13u w=0.58u m=1
M5 N_5 A VDD VDD mp15  l=0.13u w=0.58u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or02d1
* SPICE INPUT		Tue Jul 31 20:11:37 2018	or02d1p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d1p5
.subckt or02d1p5 VDD Y A B GND
M1 N_4 B GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 B N_4 VDD mp15  l=0.13u w=0.69u m=1
M5 N_5 A VDD VDD mp15  l=0.13u w=0.69u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or02d1p5
* SPICE INPUT		Tue Jul 31 20:11:50 2018	or02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d2
.subckt or02d2 Y GND VDD A B
M1 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.35u m=1
M4 N_5 B GND GND mn15  l=0.13u w=0.35u m=1
M5 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M6 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M7 N_11 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_11 B N_5 VDD mp15  l=0.13u w=0.69u m=1
.ends or02d2
* SPICE INPUT		Tue Jul 31 20:12:04 2018	or02d2p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d2p5
.subckt or02d2p5 Y VDD GND A B
M1 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_7 A VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_8 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M9 N_5 B N_7 VDD mp15  l=0.13u w=0.69u m=1
M10 N_8 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
.ends or02d2p5
* SPICE INPUT		Tue Jul 31 20:12:17 2018	or02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d4
.subckt or02d4 Y GND VDD A B
M1 N_6 A GND GND mn15  l=0.13u w=0.29u m=1
M2 N_6 B GND GND mn15  l=0.13u w=0.29u m=1
M3 N_6 B GND GND mn15  l=0.13u w=0.29u m=1
M4 N_6 A GND GND mn15  l=0.13u w=0.29u m=1
M5 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M6 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_16 A VDD VDD mp15  l=0.13u w=0.67u m=1
M10 N_17 B N_6 VDD mp15  l=0.13u w=0.67u m=1
M11 N_6 B N_16 VDD mp15  l=0.13u w=0.67u m=1
M12 N_17 A VDD VDD mp15  l=0.13u w=0.67u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or02d4
* SPICE INPUT		Tue Jul 31 20:12:31 2018	or02d4p5
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02d4p5
.subckt or02d4p5 Y GND VDD A B
M1 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_5 GND mn15  l=0.13u w=0.46u m=1
M3 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_5 A GND GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M7 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M9 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M11 N_15 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M12 N_5 B N_15 VDD mp15  l=0.13u w=0.69u m=1
M13 N_15 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD A N_15 VDD mp15  l=0.13u w=0.69u m=1
M15 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_15 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or02d4p5
* SPICE INPUT		Tue Jul 31 20:12:44 2018	or02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02dm
.subckt or02dm VDD Y GND A B
M1 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M4 N_5 B N_4 VDD mp15  l=0.13u w=0.4u m=1
M5 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends or02dm
* SPICE INPUT		Tue Jul 31 20:12:57 2018	or02od
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or02od
.subckt or02od B A GND VDD Y
M1 N_2 A GND GND mn15  l=0.13u w=0.3u m=1
M2 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M3 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M4 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M5 GND B N_2 GND mn15  l=0.13u w=0.3u m=1
M6 VDD A N_18 VDD mp15  l=0.13u w=0.6u m=1
M7 N_2 B N_18 VDD mp15  l=0.13u w=0.6u m=1
.ends or02od
* SPICE INPUT		Tue Jul 31 20:13:10 2018	or03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d0
.subckt or03d0 VDD Y GND A B C
M1 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_4 C GND GND mn15  l=0.13u w=0.26u m=1
M5 N_8 B N_7 VDD mp15  l=0.13u w=0.4u m=1
M6 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_7 C N_4 VDD mp15  l=0.13u w=0.4u m=1
.ends or03d0
* SPICE INPUT		Tue Jul 31 20:13:24 2018	or03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d1
.subckt or03d1 VDD Y GND A B C
M1 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.28u m=1
M3 N_4 B GND GND mn15  l=0.13u w=0.28u m=1
M4 N_4 C GND GND mn15  l=0.13u w=0.28u m=1
M5 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M6 N_6 A VDD VDD mp15  l=0.13u w=0.66u m=1
M7 N_6 B N_5 VDD mp15  l=0.13u w=0.66u m=1
M8 N_5 C N_4 VDD mp15  l=0.13u w=0.66u m=1
.ends or03d1
* SPICE INPUT		Tue Jul 31 20:13:37 2018	or03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d2
.subckt or03d2 Y VDD GND A B C
M1 N_4 A GND GND mn15  l=0.13u w=0.34u m=1
M2 N_4 C GND GND mn15  l=0.13u w=0.34u m=1
M3 N_4 B GND GND mn15  l=0.13u w=0.34u m=1
M4 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 VDD A N_7 VDD mp15  l=0.13u w=0.69u m=1
M7 N_6 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M8 N_7 B N_6 VDD mp15  l=0.13u w=0.69u m=1
M9 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends or03d2
* SPICE INPUT		Tue Jul 31 20:13:50 2018	or03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03d4
.subckt or03d4 Y VDD B C A GND
M1 N_5 A GND GND mn15  l=0.13u w=0.32u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND C N_5 GND mn15  l=0.13u w=0.33u m=1
M7 N_5 C GND GND mn15  l=0.13u w=0.33u m=1
M8 GND A N_5 GND mn15  l=0.13u w=0.34u m=1
M9 N_5 B GND GND mn15  l=0.13u w=0.32u m=1
M10 N_5 B GND GND mn15  l=0.13u w=0.34u m=1
M11 VDD A N_9 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M15 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M16 N_12 C N_5 VDD mp15  l=0.13u w=0.77u m=1
M17 N_5 C N_10 VDD mp15  l=0.13u w=0.61u m=1
M18 VDD A N_11 VDD mp15  l=0.13u w=0.69u m=1
M19 N_10 B N_9 VDD mp15  l=0.13u w=0.61u m=1
M20 N_12 B N_11 VDD mp15  l=0.13u w=0.77u m=1
.ends or03d4
* SPICE INPUT		Tue Jul 31 20:14:03 2018	or03dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or03dm
.subckt or03dm VDD Y GND A B C
M1 N_4 C GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.36u m=1
M4 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_7 C N_4 VDD mp15  l=0.13u w=0.4u m=1
M6 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
M8 N_8 B N_7 VDD mp15  l=0.13u w=0.4u m=1
.ends or03dm
* SPICE INPUT		Tue Jul 31 20:14:16 2018	or04d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d0
.subckt or04d0 VDD Y GND A B C D
M1 GND C N_4 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_4 D GND GND mn15  l=0.13u w=0.26u m=1
M5 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M6 N_9 C N_8 VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_8 D N_4 VDD mp15  l=0.13u w=0.4u m=1
M10 N_10 B N_9 VDD mp15  l=0.13u w=0.4u m=1
.ends or04d0
* SPICE INPUT		Tue Jul 31 20:14:28 2018	or04d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d1
.subckt or04d1 VDD Y GND A B C D
M1 N_4 D GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND C N_4 GND mn15  l=0.13u w=0.26u m=1
M4 N_4 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_4 A GND GND mn15  l=0.13u w=0.26u m=1
M6 N_8 D N_4 VDD mp15  l=0.13u w=0.4u m=1
M7 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M8 N_9 C N_8 VDD mp15  l=0.13u w=0.4u m=1
M9 N_10 B N_9 VDD mp15  l=0.13u w=0.4u m=1
M10 N_10 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends or04d1
* SPICE INPUT		Tue Jul 31 20:14:41 2018	or04d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d2
.subckt or04d2 Y VDD GND A B C D
M1 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_4 D GND GND mn15  l=0.13u w=0.28u m=1
M4 GND C N_4 GND mn15  l=0.13u w=0.28u m=1
M5 N_4 B GND GND mn15  l=0.13u w=0.28u m=1
M6 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M7 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_6 D N_4 VDD mp15  l=0.13u w=0.69u m=1
M10 N_7 C N_6 VDD mp15  l=0.13u w=0.69u m=1
M11 N_8 B N_7 VDD mp15  l=0.13u w=0.69u m=1
M12 VDD A N_8 VDD mp15  l=0.13u w=0.69u m=1
.ends or04d2
* SPICE INPUT		Tue Jul 31 20:14:54 2018	or04d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=or04d4
.subckt or04d4 Y GND VDD A B C D
M1 N_6 D GND GND mn15  l=0.13u w=0.29u m=1
M2 N_6 D GND GND mn15  l=0.13u w=0.29u m=1
M3 N_6 C GND GND mn15  l=0.13u w=0.29u m=1
M4 N_6 C GND GND mn15  l=0.13u w=0.29u m=1
M5 N_6 A GND GND mn15  l=0.13u w=0.29u m=1
M6 N_6 B GND GND mn15  l=0.13u w=0.29u m=1
M7 N_6 B GND GND mn15  l=0.13u w=0.29u m=1
M8 N_6 A GND GND mn15  l=0.13u w=0.29u m=1
M9 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M13 N_19 D N_6 VDD mp15  l=0.13u w=0.69u m=1
M14 N_6 D N_19 VDD mp15  l=0.13u w=0.69u m=1
M15 N_19 C N_18 VDD mp15  l=0.13u w=0.69u m=1
M16 N_19 C N_18 VDD mp15  l=0.13u w=0.69u m=1
M17 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_25 B N_18 VDD mp15  l=0.13u w=0.69u m=1
M19 N_18 B N_24 VDD mp15  l=0.13u w=0.69u m=1
M20 VDD A N_25 VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends or04d4
* SPICE INPUT		Tue Jul 31 20:15:07 2018	ora211d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d0
.subckt ora211d0 VDD Y GND A B C D
M1 N_11 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_11 B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_11 C N_15 GND mn15  l=0.13u w=0.26u m=1
M5 N_15 D N_4 GND mn15  l=0.13u w=0.26u m=1
M6 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_7 B N_4 VDD mp15  l=0.13u w=0.4u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_4 C VDD VDD mp15  l=0.13u w=0.27u m=1
M10 VDD D N_4 VDD mp15  l=0.13u w=0.27u m=1
.ends ora211d0
* SPICE INPUT		Tue Jul 31 20:15:20 2018	ora211d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d1
.subckt ora211d1 VDD Y GND A B C D
M1 N_11 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_11 B GND GND mn15  l=0.13u w=0.26u m=1
M3 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_11 C N_15 GND mn15  l=0.13u w=0.26u m=1
M5 N_15 D N_4 GND mn15  l=0.13u w=0.26u m=1
M6 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_7 B N_4 VDD mp15  l=0.13u w=0.4u m=1
M8 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_4 C VDD VDD mp15  l=0.13u w=0.27u m=1
M10 VDD D N_4 VDD mp15  l=0.13u w=0.27u m=1
.ends ora211d1
* SPICE INPUT		Tue Jul 31 20:15:33 2018	ora211d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d2
.subckt ora211d2 Y GND VDD D C B A
M1 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_6 C N_9 GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_6 GND mn15  l=0.13u w=0.46u m=1
M5 N_6 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_5 D N_9 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 C VDD VDD mp15  l=0.13u w=0.48u m=1
M8 N_36 A VDD VDD mp15  l=0.13u w=0.69u m=1
M9 N_36 B N_5 VDD mp15  l=0.13u w=0.69u m=1
M10 N_5 D VDD VDD mp15  l=0.13u w=0.48u m=1
M11 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ora211d2
* SPICE INPUT		Tue Jul 31 20:15:46 2018	ora211d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora211d4
.subckt ora211d4 GND Y VDD C D A B
M1 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_15 D N_8 GND mn15  l=0.13u w=0.46u m=1
M6 N_8 D N_14 GND mn15  l=0.13u w=0.46u m=1
M7 N_15 C N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_2 C N_14 GND mn15  l=0.13u w=0.46u m=1
M9 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_8 Y GND mn15  l=0.13u w=0.46u m=1
M13 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M15 VDD N_8 Y VDD mp15  l=0.13u w=0.69u m=1
M16 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_25 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_26 B N_8 VDD mp15  l=0.13u w=0.69u m=1
M19 N_8 B N_25 VDD mp15  l=0.13u w=0.69u m=1
M20 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M21 N_8 D VDD VDD mp15  l=0.13u w=0.46u m=1
M22 N_8 D VDD VDD mp15  l=0.13u w=0.46u m=1
M23 VDD C N_8 VDD mp15  l=0.13u w=0.46u m=1
M24 N_8 C VDD VDD mp15  l=0.13u w=0.46u m=1
.ends ora211d4
* SPICE INPUT		Tue Jul 31 20:15:58 2018	ora21d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d0
.subckt ora21d0 VDD Y GND C B A
M1 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_10 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C N_10 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_6 B N_5 VDD mp15  l=0.13u w=0.4u m=1
M8 N_5 C VDD VDD mp15  l=0.13u w=0.27u m=1
.ends ora21d0
* SPICE INPUT		Tue Jul 31 20:16:12 2018	ora21d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d1
.subckt ora21d1 VDD Y GND C B A
M1 N_10 A GND GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_10 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 C N_10 GND mn15  l=0.13u w=0.26u m=1
M4 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 A VDD VDD mp15  l=0.13u w=0.4u m=1
M6 N_6 B N_5 VDD mp15  l=0.13u w=0.4u m=1
M7 N_5 C VDD VDD mp15  l=0.13u w=0.27u m=1
M8 Y N_5 VDD VDD mp15  l=0.13u w=0.34u m=1
M9 Y N_5 VDD VDD mp15  l=0.13u w=0.34u m=1
.ends ora21d1
* SPICE INPUT		Tue Jul 31 20:16:24 2018	ora21d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d2
.subckt ora21d2 GND Y VDD C B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M4 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M5 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M6 N_30 A VDD VDD mp15  l=0.13u w=0.69u m=1
M7 N_30 B N_3 VDD mp15  l=0.13u w=0.69u m=1
M8 VDD C N_3 VDD mp15  l=0.13u w=0.48u m=1
M9 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ora21d2
* SPICE INPUT		Tue Jul 31 20:16:38 2018	ora21d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora21d4
.subckt ora21d4 GND Y VDD C A B
M1 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M7 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M10 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M11 N_20 A VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_21 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M13 N_2 B N_20 VDD mp15  l=0.13u w=0.69u m=1
M14 N_21 A VDD VDD mp15  l=0.13u w=0.69u m=1
M15 VDD C N_2 VDD mp15  l=0.13u w=0.48u m=1
M16 VDD C N_2 VDD mp15  l=0.13u w=0.48u m=1
M17 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M18 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M19 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M20 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora21d4
* SPICE INPUT		Tue Jul 31 20:16:51 2018	ora221d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora221d0
.subckt ora221d0 VDD Y GND E D C A B
M1 GND A N_16 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_16 GND mn15  l=0.13u w=0.26u m=1
M3 N_14 C N_16 GND mn15  l=0.13u w=0.26u m=1
M4 N_14 D N_16 GND mn15  l=0.13u w=0.26u m=1
M5 N_3 E N_14 GND mn15  l=0.13u w=0.26u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_8 B N_3 VDD mp15  l=0.13u w=0.4u m=1
M9 N_9 C VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_9 D N_3 VDD mp15  l=0.13u w=0.4u m=1
M11 N_3 E VDD VDD mp15  l=0.13u w=0.27u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ora221d0
* SPICE INPUT		Tue Jul 31 20:17:05 2018	ora221d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora221d1
.subckt ora221d1 VDD Y GND E D C A B
M1 GND B N_16 GND mn15  l=0.13u w=0.26u m=1
M2 GND A N_16 GND mn15  l=0.13u w=0.26u m=1
M3 N_14 C N_16 GND mn15  l=0.13u w=0.26u m=1
M4 N_14 D N_16 GND mn15  l=0.13u w=0.26u m=1
M5 N_3 E N_14 GND mn15  l=0.13u w=0.26u m=1
M6 Y N_3 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_8 B N_3 VDD mp15  l=0.13u w=0.4u m=1
M8 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_9 C VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_9 D N_3 VDD mp15  l=0.13u w=0.4u m=1
M11 N_3 E VDD VDD mp15  l=0.13u w=0.27u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora221d1
* SPICE INPUT		Tue Jul 31 20:17:18 2018	ora221d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora221d2
.subckt ora221d2 Y GND VDD E D C A B
M1 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_6 C N_5 GND mn15  l=0.13u w=0.46u m=1
M5 N_5 B GND GND mn15  l=0.13u w=0.46u m=1
M6 N_10 E N_6 GND mn15  l=0.13u w=0.46u m=1
M7 N_5 D N_6 GND mn15  l=0.13u w=0.46u m=1
M8 VDD E N_10 VDD mp15  l=0.13u w=0.48u m=1
M9 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M10 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M11 N_15 D N_10 VDD mp15  l=0.13u w=0.35u m=1
M12 N_15 D N_10 VDD mp15  l=0.13u w=0.34u m=1
M13 VDD A N_44 VDD mp15  l=0.13u w=0.69u m=1
M14 VDD C N_15 VDD mp15  l=0.13u w=0.69u m=1
M15 N_44 B N_10 VDD mp15  l=0.13u w=0.69u m=1
.ends ora221d2
* SPICE INPUT		Tue Jul 31 20:17:32 2018	ora221d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora221d4
.subckt ora221d4 GND Y VDD E D C A B
M1 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M2 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_2 C N_3 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M7 N_2 D N_3 GND mn15  l=0.13u w=0.565u m=1
M8 N_3 D N_2 GND mn15  l=0.13u w=0.355u m=1
M9 GND N_16 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_16 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_16 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_16 Y GND mn15  l=0.13u w=0.46u m=1
M13 N_3 E N_16 GND mn15  l=0.13u w=0.565u m=1
M14 N_3 E N_16 GND mn15  l=0.13u w=0.355u m=1
M15 N_16 B N_28 VDD mp15  l=0.13u w=0.69u m=1
M16 N_16 B N_24 VDD mp15  l=0.13u w=0.69u m=1
M17 N_28 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_24 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_19 C VDD VDD mp15  l=0.13u w=0.46u m=1
M20 VDD C N_19 VDD mp15  l=0.13u w=0.46u m=1
M21 N_19 C VDD VDD mp15  l=0.13u w=0.46u m=1
M22 N_16 D N_19 VDD mp15  l=0.13u w=0.56u m=1
M23 N_16 D N_19 VDD mp15  l=0.13u w=0.56u m=1
M24 N_16 D N_19 VDD mp15  l=0.13u w=0.26u m=1
M25 N_16 E VDD VDD mp15  l=0.13u w=0.6u m=1
M26 N_16 E VDD VDD mp15  l=0.13u w=0.36u m=1
M27 VDD N_16 Y VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_16 Y VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_16 Y VDD mp15  l=0.13u w=0.69u m=1
M30 Y N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora221d4
* SPICE INPUT		Tue Jul 31 20:17:45 2018	ora222d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora222d0
.subckt ora222d0 VDD Y GND F E C D B A
M1 GND A N_19 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_19 GND mn15  l=0.13u w=0.26u m=1
M3 N_17 D N_19 GND mn15  l=0.13u w=0.26u m=1
M4 N_19 C N_17 GND mn15  l=0.13u w=0.26u m=1
M5 N_2 E N_17 GND mn15  l=0.13u w=0.26u m=1
M6 N_2 F N_17 GND mn15  l=0.13u w=0.26u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_2 B N_12 VDD mp15  l=0.13u w=0.4u m=1
M10 N_13 D N_2 VDD mp15  l=0.13u w=0.4u m=1
M11 N_13 C VDD VDD mp15  l=0.13u w=0.4u m=1
M12 VDD E N_11 VDD mp15  l=0.13u w=0.4u m=1
M13 N_2 F N_11 VDD mp15  l=0.13u w=0.4u m=1
M14 Y N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ora222d0
* SPICE INPUT		Tue Jul 31 20:17:58 2018	ora222d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora222d1
.subckt ora222d1 VDD Y GND F E C D B A
M1 GND A N_19 GND mn15  l=0.13u w=0.26u m=1
M2 GND B N_19 GND mn15  l=0.13u w=0.26u m=1
M3 N_17 D N_19 GND mn15  l=0.13u w=0.26u m=1
M4 N_19 C N_17 GND mn15  l=0.13u w=0.26u m=1
M5 N_2 E N_17 GND mn15  l=0.13u w=0.26u m=1
M6 N_2 F N_17 GND mn15  l=0.13u w=0.26u m=1
M7 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_12 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_2 B N_12 VDD mp15  l=0.13u w=0.4u m=1
M10 N_13 D N_2 VDD mp15  l=0.13u w=0.4u m=1
M11 N_13 C VDD VDD mp15  l=0.13u w=0.4u m=1
M12 VDD E N_11 VDD mp15  l=0.13u w=0.4u m=1
M13 N_2 F N_11 VDD mp15  l=0.13u w=0.4u m=1
M14 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora222d1
* SPICE INPUT		Tue Jul 31 20:18:11 2018	ora222d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora222d2
.subckt ora222d2 GND Y VDD E F C D B A
M1 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_2 D N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 E N_7 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 F N_7 GND mn15  l=0.13u w=0.46u m=1
M7 GND N_7 Y GND mn15  l=0.13u w=0.46u m=1
M8 GND N_7 Y GND mn15  l=0.13u w=0.46u m=1
M9 N_7 D N_24 VDD mp15  l=0.13u w=0.34u m=1
M10 N_25 A VDD VDD mp15  l=0.13u w=0.69u m=1
M11 N_25 B N_7 VDD mp15  l=0.13u w=0.69u m=1
M12 N_26 D N_7 VDD mp15  l=0.13u w=0.35u m=1
M13 N_26 C VDD VDD mp15  l=0.13u w=0.35u m=1
M14 VDD C N_24 VDD mp15  l=0.13u w=0.34u m=1
M15 VDD N_7 Y VDD mp15  l=0.13u w=0.69u m=1
M16 VDD N_7 Y VDD mp15  l=0.13u w=0.69u m=1
M17 VDD E N_27 VDD mp15  l=0.13u w=0.69u m=1
M18 N_27 F N_7 VDD mp15  l=0.13u w=0.69u m=1
.ends ora222d2
* SPICE INPUT		Tue Jul 31 20:18:24 2018	ora222d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora222d4
.subckt ora222d4 GND Y F VDD E C D B A
M1 N_2 B GND GND mn15  l=0.13u w=0.46u m=1
M2 GND A N_2 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 A GND GND mn15  l=0.13u w=0.46u m=1
M4 GND B N_2 GND mn15  l=0.13u w=0.46u m=1
M5 N_3 D N_2 GND mn15  l=0.13u w=0.45u m=1
M6 N_2 C N_3 GND mn15  l=0.13u w=0.56u m=1
M7 N_2 C N_3 GND mn15  l=0.13u w=0.36u m=1
M8 N_3 D N_2 GND mn15  l=0.13u w=0.47u m=1
M9 N_3 F N_11 GND mn15  l=0.13u w=0.565u m=1
M10 N_3 F N_11 GND mn15  l=0.13u w=0.355u m=1
M11 N_3 E N_11 GND mn15  l=0.13u w=0.565u m=1
M12 N_3 E N_11 GND mn15  l=0.13u w=0.355u m=1
M13 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M14 Y N_11 GND GND mn15  l=0.13u w=0.46u m=1
M15 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M16 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M17 N_37 B N_11 VDD mp15  l=0.13u w=0.69u m=1
M18 N_38 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_37 A VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_11 B N_38 VDD mp15  l=0.13u w=0.69u m=1
M21 N_11 F N_36 VDD mp15  l=0.13u w=0.55u m=1
M22 N_42 E VDD VDD mp15  l=0.13u w=0.42u m=1
M23 VDD E N_36 VDD mp15  l=0.13u w=0.55u m=1
M24 VDD E N_43 VDD mp15  l=0.13u w=0.41u m=1
M25 N_11 D N_39 VDD mp15  l=0.13u w=0.69u m=1
M26 N_40 C VDD VDD mp15  l=0.13u w=0.27u m=1
M27 VDD C N_39 VDD mp15  l=0.13u w=0.605u m=1
M28 N_40 D N_11 VDD mp15  l=0.13u w=0.27u m=1
M29 N_41 D N_11 VDD mp15  l=0.13u w=0.42u m=1
M30 N_41 C VDD VDD mp15  l=0.13u w=0.505u m=1
M31 N_43 F N_11 VDD mp15  l=0.13u w=0.41u m=1
M32 N_11 F N_42 VDD mp15  l=0.13u w=0.42u m=1
M33 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
M34 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
M36 Y N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora222d4
* SPICE INPUT		Tue Jul 31 20:18:37 2018	ora22d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora22d0
.subckt ora22d0 VDD Y GND C D B A
M1 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_13 D N_4 GND mn15  l=0.13u w=0.26u m=1
M3 N_13 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_13 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_13 C N_4 GND mn15  l=0.13u w=0.26u m=1
M6 N_4 D N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_4 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M9 VDD C N_7 VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ora22d0
* SPICE INPUT		Tue Jul 31 20:18:51 2018	ora22d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora22d1
.subckt ora22d1 VDD Y GND C D B A
M1 Y N_4 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_13 D N_4 GND mn15  l=0.13u w=0.26u m=1
M3 N_13 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_13 B GND GND mn15  l=0.13u w=0.26u m=1
M5 N_13 C N_4 GND mn15  l=0.13u w=0.26u m=1
M6 N_4 D N_7 VDD mp15  l=0.13u w=0.4u m=1
M7 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M8 N_4 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M9 VDD C N_7 VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora22d1
* SPICE INPUT		Tue Jul 31 20:19:03 2018	ora22d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora22d2
.subckt ora22d2 Y GND VDD C D B A
M1 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_5 Y GND mn15  l=0.13u w=0.46u m=1
M3 N_6 C N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_6 B GND GND mn15  l=0.13u w=0.46u m=1
M5 N_6 D N_5 GND mn15  l=0.13u w=0.46u m=1
M6 GND A N_6 GND mn15  l=0.13u w=0.46u m=1
M7 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M8 VDD N_5 Y VDD mp15  l=0.13u w=0.69u m=1
M9 N_12 C VDD VDD mp15  l=0.13u w=0.345u m=1
M10 N_12 C VDD VDD mp15  l=0.13u w=0.345u m=1
M11 N_5 B N_17 VDD mp15  l=0.13u w=0.69u m=1
M12 N_5 D N_12 VDD mp15  l=0.13u w=0.69u m=1
M13 N_17 A VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora22d2
* SPICE INPUT		Tue Jul 31 20:19:16 2018	ora22d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora22d4
.subckt ora22d4 GND Y VDD C D A B
M1 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M2 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M4 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M6 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M7 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M8 N_3 C N_2 GND mn15  l=0.13u w=0.46u m=1
M9 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M13 N_26 A VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_27 B N_2 VDD mp15  l=0.13u w=0.69u m=1
M15 N_2 B N_26 VDD mp15  l=0.13u w=0.69u m=1
M16 N_27 A VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_2 D N_25 VDD mp15  l=0.13u w=0.6u m=1
M18 N_2 D N_28 VDD mp15  l=0.13u w=0.6u m=1
M19 N_25 C VDD VDD mp15  l=0.13u w=0.6u m=1
M20 N_28 C VDD VDD mp15  l=0.13u w=0.6u m=1
M21 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora22d4
* SPICE INPUT		Tue Jul 31 20:19:29 2018	ora31d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d0
.subckt ora31d0 VDD Y A B C GND D
M1 N_11 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_11 B GND GND mn15  l=0.13u w=0.26u m=1
M3 N_11 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_11 D N_5 GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_9 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_9 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M8 N_8 C N_5 VDD mp15  l=0.13u w=0.4u m=1
M9 N_5 D VDD VDD mp15  l=0.13u w=0.27u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends ora31d0
* SPICE INPUT		Tue Jul 31 20:19:42 2018	ora31d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d1
.subckt ora31d1 VDD Y GND A B C D
M1 N_12 A GND GND mn15  l=0.13u w=0.26u m=1
M2 N_12 D N_5 GND mn15  l=0.13u w=0.26u m=1
M3 N_12 C GND GND mn15  l=0.13u w=0.26u m=1
M4 N_12 B GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_5 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_9 A VDD VDD mp15  l=0.13u w=0.4u m=1
M7 N_5 D VDD VDD mp15  l=0.13u w=0.27u m=1
M8 N_8 C N_5 VDD mp15  l=0.13u w=0.4u m=1
M9 N_9 B N_8 VDD mp15  l=0.13u w=0.4u m=1
M10 Y N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora31d1
* SPICE INPUT		Tue Jul 31 20:19:55 2018	ora31d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d2
.subckt ora31d2 Y GND VDD A B C D
M1 N_6 D N_4 GND mn15  l=0.13u w=0.46u m=1
M2 N_6 C GND GND mn15  l=0.13u w=0.46u m=1
M3 N_6 B GND GND mn15  l=0.13u w=0.46u m=1
M4 GND A N_6 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M6 GND N_4 Y GND mn15  l=0.13u w=0.46u m=1
M7 N_4 D VDD VDD mp15  l=0.13u w=0.48u m=1
M8 N_31 C N_4 VDD mp15  l=0.13u w=0.69u m=1
M9 N_32 B N_31 VDD mp15  l=0.13u w=0.69u m=1
M10 VDD A N_32 VDD mp15  l=0.13u w=0.69u m=1
M11 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
M12 VDD N_4 Y VDD mp15  l=0.13u w=0.69u m=1
.ends ora31d2
* SPICE INPUT		Tue Jul 31 20:20:08 2018	ora31d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=ora31d4
.subckt ora31d4 GND Y D VDD C B A
M1 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M2 N_3 D N_2 GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_3 GND mn15  l=0.13u w=0.46u m=1
M4 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M5 N_3 C GND GND mn15  l=0.13u w=0.46u m=1
M6 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M7 N_3 B GND GND mn15  l=0.13u w=0.46u m=1
M8 N_3 A GND GND mn15  l=0.13u w=0.46u m=1
M9 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M10 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M13 VDD D N_2 VDD mp15  l=0.13u w=0.48u m=1
M14 VDD D N_2 VDD mp15  l=0.13u w=0.48u m=1
M15 N_60 C N_2 VDD mp15  l=0.13u w=0.69u m=1
M16 N_61 B N_60 VDD mp15  l=0.13u w=0.69u m=1
M17 N_61 A VDD VDD mp15  l=0.13u w=0.69u m=1
M18 N_62 A VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_63 C N_2 VDD mp15  l=0.13u w=0.69u m=1
M20 N_63 B N_62 VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends ora31d4
* SPICE INPUT		Tue Jul 31 20:20:21 2018	pulld
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=pulld
.subckt pulld GND Y VDD EN
M1 N_4 EN GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 GND GND mn15  l=0.13u w=0.26u m=1
M3 VDD EN N_4 VDD mp15  l=0.13u w=0.4u m=1
.ends pulld
* SPICE INPUT		Tue Jul 31 20:20:34 2018	pullu
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=pullu
.subckt pullu VDD Y GND E
M1 GND E N_4 GND mn15  l=0.13u w=0.26u m=1
M2 Y N_4 VDD VDD mp15  l=0.13u w=0.26u m=1
M3 N_4 E VDD VDD mp15  l=0.13u w=0.4u m=1
.ends pullu
* SPICE INPUT		Tue Jul 31 20:20:46 2018	sdanrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdanrq0
.subckt sdanrq0 GND Q VDD CK SE SI D1 D0
M1 N_18 D0 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 D1 N_18 GND mn15  l=0.13u w=0.26u m=1
M3 N_19 SE N_6 GND mn15  l=0.13u w=0.24u m=1
M4 N_6 N_2 N_5 GND mn15  l=0.13u w=0.28u m=1
M5 N_19 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND SE N_2 GND mn15  l=0.13u w=0.18u m=1
M7 GND CK N_8 GND mn15  l=0.13u w=0.17u m=1
M8 N_20 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M9 N_20 N_8 N_10 GND mn15  l=0.13u w=0.28u m=1
M10 N_21 N_7 N_10 GND mn15  l=0.13u w=0.17u m=1
M11 GND N_13 N_21 GND mn15  l=0.13u w=0.17u m=1
M12 N_13 N_10 GND GND mn15  l=0.13u w=0.28u m=1
M13 N_13 N_7 N_12 GND mn15  l=0.13u w=0.28u m=1
M14 N_22 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M15 N_22 N_8 N_12 GND mn15  l=0.13u w=0.17u m=1
M16 GND N_8 N_7 GND mn15  l=0.13u w=0.17u m=1
M17 Q N_12 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_17 N_12 GND GND mn15  l=0.13u w=0.18u m=1
M19 VDD D0 N_5 VDD mp15  l=0.13u w=0.35u m=1
M20 N_5 D1 VDD VDD mp15  l=0.13u w=0.35u m=1
M21 N_38 N_2 N_6 VDD mp15  l=0.13u w=0.37u m=1
M22 N_38 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M23 N_6 SE N_5 VDD mp15  l=0.13u w=0.42u m=1
M24 N_2 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M25 N_8 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M26 N_39 N_6 VDD VDD mp15  l=0.13u w=0.42u m=1
M27 N_10 N_7 N_39 VDD mp15  l=0.13u w=0.42u m=1
M28 N_40 N_8 N_10 VDD mp15  l=0.13u w=0.17u m=1
M29 VDD N_13 N_40 VDD mp15  l=0.13u w=0.17u m=1
M30 N_13 N_10 VDD VDD mp15  l=0.13u w=0.42u m=1
M31 N_41 N_7 N_12 VDD mp15  l=0.13u w=0.17u m=1
M32 N_41 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M33 N_7 N_8 VDD VDD mp15  l=0.13u w=0.42u m=1
M34 N_12 N_8 N_13 VDD mp15  l=0.13u w=0.42u m=1
M35 Q N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M36 N_17 N_12 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends sdanrq0
* SPICE INPUT		Tue Jul 31 20:20:59 2018	sdanrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdanrq1
.subckt sdanrq1 GND Q CK SE D1 SI D0 VDD
M1 N_18 D0 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 D1 N_18 GND mn15  l=0.13u w=0.26u m=1
M3 N_6 N_2 N_5 GND mn15  l=0.13u w=0.28u m=1
M4 N_19 SE N_6 GND mn15  l=0.13u w=0.24u m=1
M5 N_19 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND SE N_2 GND mn15  l=0.13u w=0.18u m=1
M7 GND CK N_9 GND mn15  l=0.13u w=0.2u m=1
M8 N_20 N_9 N_11 GND mn15  l=0.13u w=0.28u m=1
M9 N_21 N_7 N_11 GND mn15  l=0.13u w=0.17u m=1
M10 N_20 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M11 GND N_9 N_7 GND mn15  l=0.13u w=0.2u m=1
M12 N_22 N_9 N_14 GND mn15  l=0.13u w=0.17u m=1
M13 N_22 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M14 GND N_13 N_21 GND mn15  l=0.13u w=0.17u m=1
M15 N_13 N_11 GND GND mn15  l=0.13u w=0.36u m=1
M16 N_14 N_7 N_13 GND mn15  l=0.13u w=0.36u m=1
M17 Q N_14 GND GND mn15  l=0.13u w=0.46u m=1
M18 N_17 N_14 GND GND mn15  l=0.13u w=0.28u m=1
M19 VDD D0 N_5 VDD mp15  l=0.13u w=0.35u m=1
M20 N_5 D1 VDD VDD mp15  l=0.13u w=0.35u m=1
M21 N_38 N_2 N_6 VDD mp15  l=0.13u w=0.37u m=1
M22 N_38 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M23 N_6 SE N_5 VDD mp15  l=0.13u w=0.42u m=1
M24 VDD SE N_2 VDD mp15  l=0.13u w=0.28u m=1
M25 N_9 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M26 N_11 N_7 N_39 VDD mp15  l=0.13u w=0.42u m=1
M27 N_39 N_6 VDD VDD mp15  l=0.13u w=0.42u m=1
M28 N_13 N_9 N_14 VDD mp15  l=0.13u w=0.52u m=1
M29 N_7 N_9 VDD VDD mp15  l=0.13u w=0.51u m=1
M30 N_41 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M31 N_41 N_7 N_14 VDD mp15  l=0.13u w=0.17u m=1
M32 N_40 N_9 N_11 VDD mp15  l=0.13u w=0.17u m=1
M33 VDD N_13 N_40 VDD mp15  l=0.13u w=0.17u m=1
M34 N_13 N_11 VDD VDD mp15  l=0.13u w=0.52u m=1
M35 Q N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 N_17 N_14 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends sdanrq1
* SPICE INPUT		Tue Jul 31 20:21:12 2018	sdanrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdanrq2
.subckt sdanrq2 GND Q CK SE SI VDD D1 D0
M1 N_2 D1 N_20 GND mn15  l=0.13u w=0.46u m=1
M2 GND D0 N_20 GND mn15  l=0.13u w=0.46u m=1
M3 GND N_14 Q GND mn15  l=0.13u w=0.46u m=1
M4 GND N_14 Q GND mn15  l=0.13u w=0.46u m=1
M5 GND N_14 N_6 GND mn15  l=0.13u w=0.37u m=1
M6 N_23 N_9 N_14 GND mn15  l=0.13u w=0.17u m=1
M7 GND N_9 N_8 GND mn15  l=0.13u w=0.23u m=1
M8 N_14 N_8 N_13 GND mn15  l=0.13u w=0.41u m=1
M9 GND N_13 N_22 GND mn15  l=0.13u w=0.17u m=1
M10 N_23 N_6 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_13 N_11 GND GND mn15  l=0.13u w=0.41u m=1
M12 N_22 N_8 N_11 GND mn15  l=0.13u w=0.17u m=1
M13 GND CK N_9 GND mn15  l=0.13u w=0.28u m=1
M14 N_21 N_9 N_11 GND mn15  l=0.13u w=0.41u m=1
M15 N_21 N_18 GND GND mn15  l=0.13u w=0.41u m=1
M16 N_24 SE N_18 GND mn15  l=0.13u w=0.28u m=1
M17 GND SE N_16 GND mn15  l=0.13u w=0.24u m=1
M18 N_2 N_16 N_18 GND mn15  l=0.13u w=0.41u m=1
M19 N_24 SI GND GND mn15  l=0.13u w=0.28u m=1
M20 Q N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_14 Q VDD mp15  l=0.13u w=0.69u m=1
M22 N_6 N_14 VDD VDD mp15  l=0.13u w=0.55u m=1
M23 N_14 N_9 N_13 VDD mp15  l=0.13u w=0.63u m=1
M24 VDD N_9 N_8 VDD mp15  l=0.13u w=0.55u m=1
M25 N_98 N_8 N_14 VDD mp15  l=0.13u w=0.17u m=1
M26 N_98 N_6 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_100 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 N_13 N_11 VDD VDD mp15  l=0.13u w=0.315u m=1
M29 N_13 N_11 VDD VDD mp15  l=0.13u w=0.315u m=1
M30 N_99 N_8 N_11 VDD mp15  l=0.13u w=0.62u m=1
M31 N_100 N_9 N_11 VDD mp15  l=0.13u w=0.17u m=1
M32 N_9 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M33 N_99 N_18 VDD VDD mp15  l=0.13u w=0.62u m=1
M34 VDD SE N_16 VDD mp15  l=0.13u w=0.37u m=1
M35 N_2 D1 VDD VDD mp15  l=0.13u w=0.61u m=1
M36 N_101 N_16 N_18 VDD mp15  l=0.13u w=0.42u m=1
M37 VDD D0 N_2 VDD mp15  l=0.13u w=0.61u m=1
M38 N_101 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M39 N_18 SE N_2 VDD mp15  l=0.13u w=0.63u m=1
.ends sdanrq2
* SPICE INPUT		Tue Jul 31 20:21:25 2018	sdbfb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb0
.subckt sdbfb0 VDD Q QN SN RN GND CKN SI D SE
M1 N_110 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_110 N_5 N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_111 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_5 GND mn15  l=0.13u w=0.18u m=1
M5 N_111 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CKN N_3 GND mn15  l=0.13u w=0.18u m=1
M7 N_112 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M8 GND N_3 N_7 GND mn15  l=0.13u w=0.17u m=1
M9 N_112 N_3 N_10 GND mn15  l=0.13u w=0.17u m=1
M10 N_10 N_7 N_6 GND mn15  l=0.13u w=0.18u m=1
M11 N_12 N_10 N_36 GND mn15  l=0.13u w=0.14u m=1
M12 N_36 N_10 N_12 GND mn15  l=0.13u w=0.14u m=1
M13 N_14 N_3 N_12 GND mn15  l=0.13u w=0.28u m=1
M14 N_113 N_7 N_14 GND mn15  l=0.13u w=0.17u m=1
M15 N_36 N_21 N_14 GND mn15  l=0.13u w=0.2u m=1
M16 N_113 N_26 N_36 GND mn15  l=0.13u w=0.17u m=1
M17 QN N_14 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_26 N_14 GND GND mn15  l=0.13u w=0.18u m=1
M19 GND RN N_21 GND mn15  l=0.13u w=0.18u m=1
M20 N_36 SN GND GND mn15  l=0.13u w=0.19u m=1
M21 N_36 SN GND GND mn15  l=0.13u w=0.17u m=1
M22 Q N_26 GND GND mn15  l=0.13u w=0.26u m=1
M23 N_27 D VDD VDD mp15  l=0.13u w=0.37u m=1
M24 N_27 SE N_6 VDD mp15  l=0.13u w=0.37u m=1
M25 N_5 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M26 N_28 N_5 N_6 VDD mp15  l=0.13u w=0.28u m=1
M27 N_28 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M28 N_3 CKN VDD VDD mp15  l=0.13u w=0.46u m=1
M29 N_29 N_12 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 N_10 N_3 N_6 VDD mp15  l=0.13u w=0.5u m=1
M31 VDD N_3 N_7 VDD mp15  l=0.13u w=0.42u m=1
M32 N_29 N_7 N_10 VDD mp15  l=0.13u w=0.17u m=1
M33 N_12 N_10 N_11 VDD mp15  l=0.13u w=0.3u m=1
M34 N_11 N_10 N_12 VDD mp15  l=0.13u w=0.17u m=1
M35 N_14 N_3 N_30 VDD mp15  l=0.13u w=0.17u m=1
M36 N_30 N_26 N_11 VDD mp15  l=0.13u w=0.17u m=1
M37 N_12 N_7 N_14 VDD mp15  l=0.13u w=0.46u m=1
M38 N_11 N_21 VDD VDD mp15  l=0.13u w=0.315u m=1
M39 VDD N_21 N_11 VDD mp15  l=0.13u w=0.315u m=1
M40 N_21 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M41 N_14 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M42 Q N_26 VDD VDD mp15  l=0.13u w=0.4u m=1
M43 QN N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M44 N_26 N_14 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends sdbfb0
* SPICE INPUT		Tue Jul 31 20:21:38 2018	sdbfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb1
.subckt sdbfb1 VDD QN Q GND CKN RN SI SN D SE
M1 N_110 D GND GND mn15  l=0.13u w=0.28u m=1
M2 N_110 N_5 N_6 GND mn15  l=0.13u w=0.28u m=1
M3 N_111 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_5 GND mn15  l=0.13u w=0.18u m=1
M5 N_111 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CKN N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_112 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M8 GND N_2 N_7 GND mn15  l=0.13u w=0.2u m=1
M9 N_112 N_2 N_10 GND mn15  l=0.13u w=0.17u m=1
M10 N_10 N_7 N_6 GND mn15  l=0.13u w=0.3u m=1
M11 N_113 N_18 N_39 GND mn15  l=0.13u w=0.17u m=1
M12 N_12 N_10 N_39 GND mn15  l=0.13u w=0.165u m=1
M13 N_39 N_10 N_12 GND mn15  l=0.13u w=0.165u m=1
M14 N_14 N_2 N_12 GND mn15  l=0.13u w=0.4u m=1
M15 N_113 N_7 N_14 GND mn15  l=0.13u w=0.17u m=1
M16 N_14 N_24 N_39 GND mn15  l=0.13u w=0.27u m=1
M17 QN N_14 GND GND mn15  l=0.13u w=0.46u m=1
M18 N_18 N_14 GND GND mn15  l=0.13u w=0.27u m=1
M19 GND RN N_24 GND mn15  l=0.13u w=0.17u m=1
M20 N_39 SN GND GND mn15  l=0.13u w=0.27u m=1
M21 N_39 SN GND GND mn15  l=0.13u w=0.19u m=1
M22 Q N_18 GND GND mn15  l=0.13u w=0.46u m=1
M23 N_27 D VDD VDD mp15  l=0.13u w=0.42u m=1
M24 N_27 SE N_6 VDD mp15  l=0.13u w=0.42u m=1
M25 N_5 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M26 N_28 N_5 N_6 VDD mp15  l=0.13u w=0.28u m=1
M27 N_28 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M28 VDD CKN N_2 VDD mp15  l=0.13u w=0.51u m=1
M29 N_29 N_12 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 VDD N_2 N_7 VDD mp15  l=0.13u w=0.51u m=1
M31 N_10 N_2 N_6 VDD mp15  l=0.13u w=0.48u m=1
M32 N_29 N_7 N_10 VDD mp15  l=0.13u w=0.17u m=1
M33 N_12 N_10 N_11 VDD mp15  l=0.13u w=0.315u m=1
M34 N_11 N_10 N_12 VDD mp15  l=0.13u w=0.315u m=1
M35 N_14 N_2 N_30 VDD mp15  l=0.13u w=0.17u m=1
M36 N_30 N_18 N_11 VDD mp15  l=0.13u w=0.17u m=1
M37 N_12 N_7 N_14 VDD mp15  l=0.13u w=0.565u m=1
M38 QN N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 N_18 N_14 VDD VDD mp15  l=0.13u w=0.39u m=1
M40 N_11 N_24 VDD VDD mp15  l=0.13u w=0.35u m=1
M41 VDD N_24 N_11 VDD mp15  l=0.13u w=0.35u m=1
M42 N_24 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M43 N_14 SN VDD VDD mp15  l=0.13u w=0.35u m=1
M44 Q N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends sdbfb1
* SPICE INPUT		Tue Jul 31 20:21:51 2018	sdbfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbfb2
.subckt sdbfb2 Q VDD QN SE SI SN RN CKN GND D
M1 GND N_9 QN GND mn15  l=0.13u w=0.46u m=1
M2 QN N_9 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND N_9 N_5 GND mn15  l=0.13u w=0.36u m=1
M4 GND N_5 Q GND mn15  l=0.13u w=0.46u m=1
M5 GND N_5 Q GND mn15  l=0.13u w=0.43u m=1
M6 GND SN N_46 GND mn15  l=0.13u w=0.28u m=1
M7 N_46 SN GND GND mn15  l=0.13u w=0.32u m=1
M8 N_46 SN GND GND mn15  l=0.13u w=0.32u m=1
M9 N_10 RN GND GND mn15  l=0.13u w=0.27u m=1
M10 N_27 CKN GND GND mn15  l=0.13u w=0.27u m=1
M11 N_128 SE N_24 GND mn15  l=0.13u w=0.27u m=1
M12 GND SE N_29 GND mn15  l=0.13u w=0.24u m=1
M13 N_127 N_29 N_24 GND mn15  l=0.13u w=0.36u m=1
M14 N_128 SI GND GND mn15  l=0.13u w=0.27u m=1
M15 N_127 D GND GND mn15  l=0.13u w=0.36u m=1
M16 N_129 N_5 N_46 GND mn15  l=0.13u w=0.17u m=1
M17 N_9 N_10 N_46 GND mn15  l=0.13u w=0.36u m=1
M18 N_129 N_22 N_9 GND mn15  l=0.13u w=0.17u m=1
M19 N_9 N_27 N_13 GND mn15  l=0.13u w=0.46u m=1
M20 N_13 N_25 N_46 GND mn15  l=0.13u w=0.22u m=1
M21 N_46 N_25 N_13 GND mn15  l=0.13u w=0.22u m=1
M22 N_13 N_25 N_46 GND mn15  l=0.13u w=0.22u m=1
M23 N_25 N_22 N_24 GND mn15  l=0.13u w=0.35u m=1
M24 GND N_27 N_22 GND mn15  l=0.13u w=0.22u m=1
M25 N_130 N_27 N_25 GND mn15  l=0.13u w=0.17u m=1
M26 N_130 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M27 QN N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 QN N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 N_5 N_9 VDD VDD mp15  l=0.13u w=0.52u m=1
M30 VDD N_5 Q VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_5 Q VDD mp15  l=0.13u w=0.69u m=1
M32 N_9 SN VDD VDD mp15  l=0.13u w=0.55u m=1
M33 N_10 RN VDD VDD mp15  l=0.13u w=0.4u m=1
M34 N_14 N_5 N_31 VDD mp15  l=0.13u w=0.17u m=1
M35 N_14 N_10 VDD VDD mp15  l=0.13u w=0.45u m=1
M36 N_14 N_10 VDD VDD mp15  l=0.13u w=0.45u m=1
M37 VDD N_10 N_14 VDD mp15  l=0.13u w=0.44u m=1
M38 N_31 N_27 N_9 VDD mp15  l=0.13u w=0.17u m=1
M39 N_13 N_22 N_9 VDD mp15  l=0.13u w=0.7u m=1
M40 N_13 N_25 N_14 VDD mp15  l=0.13u w=0.315u m=1
M41 N_14 N_25 N_13 VDD mp15  l=0.13u w=0.315u m=1
M42 N_13 N_25 N_14 VDD mp15  l=0.13u w=0.315u m=1
M43 N_13 N_25 N_14 VDD mp15  l=0.13u w=0.315u m=1
M44 N_32 N_22 N_25 VDD mp15  l=0.13u w=0.17u m=1
M45 VDD N_27 N_22 VDD mp15  l=0.13u w=0.55u m=1
M46 N_25 N_27 N_24 VDD mp15  l=0.13u w=0.52u m=1
M47 N_32 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M48 N_27 CKN VDD VDD mp15  l=0.13u w=0.69u m=1
M49 N_24 SE N_33 VDD mp15  l=0.13u w=0.51u m=1
M50 N_29 SE VDD VDD mp15  l=0.13u w=0.37u m=1
M51 N_34 N_29 N_24 VDD mp15  l=0.13u w=0.4u m=1
M52 N_34 SI VDD VDD mp15  l=0.13u w=0.4u m=1
M53 N_33 D VDD VDD mp15  l=0.13u w=0.51u m=1
.ends sdbfb2
* SPICE INPUT		Tue Jul 31 20:22:05 2018	sdbrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb0
.subckt sdbrb0 VDD Q QN SN RN GND CK SI D SE
M1 N_106 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_106 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 N_107 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_5 GND mn15  l=0.13u w=0.18u m=1
M5 N_107 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_3 GND mn15  l=0.13u w=0.18u m=1
M7 N_10 N_3 N_6 GND mn15  l=0.13u w=0.18u m=1
M8 N_108 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_108 N_7 N_10 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_3 N_7 GND mn15  l=0.13u w=0.17u m=1
M11 QN N_14 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_24 N_14 GND GND mn15  l=0.13u w=0.18u m=1
M13 N_34 N_10 N_12 GND mn15  l=0.13u w=0.14u m=1
M14 N_12 N_10 N_34 GND mn15  l=0.13u w=0.14u m=1
M15 N_14 N_7 N_12 GND mn15  l=0.13u w=0.28u m=1
M16 N_109 N_3 N_14 GND mn15  l=0.13u w=0.17u m=1
M17 N_34 N_19 N_14 GND mn15  l=0.13u w=0.2u m=1
M18 N_109 N_24 N_34 GND mn15  l=0.13u w=0.17u m=1
M19 N_19 RN GND GND mn15  l=0.13u w=0.18u m=1
M20 GND SN N_34 GND mn15  l=0.13u w=0.28u m=1
M21 Q N_24 GND GND mn15  l=0.13u w=0.26u m=1
M22 N_25 D VDD VDD mp15  l=0.13u w=0.28u m=1
M23 N_26 N_5 N_6 VDD mp15  l=0.13u w=0.28u m=1
M24 N_25 SE N_6 VDD mp15  l=0.13u w=0.28u m=1
M25 N_5 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M26 N_26 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M27 N_3 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M28 N_27 N_12 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_10 N_7 N_6 VDD mp15  l=0.13u w=0.28u m=1
M30 VDD N_3 N_7 VDD mp15  l=0.13u w=0.42u m=1
M31 N_27 N_3 N_10 VDD mp15  l=0.13u w=0.17u m=1
M32 N_11 N_10 N_12 VDD mp15  l=0.13u w=0.47u m=1
M33 N_14 N_7 N_28 VDD mp15  l=0.13u w=0.17u m=1
M34 N_28 N_24 N_11 VDD mp15  l=0.13u w=0.17u m=1
M35 N_14 N_3 N_12 VDD mp15  l=0.13u w=0.46u m=1
M36 VDD N_19 N_11 VDD mp15  l=0.13u w=0.47u m=1
M37 N_19 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M38 N_14 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M39 Q N_24 VDD VDD mp15  l=0.13u w=0.4u m=1
M40 QN N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M41 N_24 N_14 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends sdbrb0
* SPICE INPUT		Tue Jul 31 20:22:18 2018	sdbrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb1
.subckt sdbrb1 GND Q QN VDD SN RN CK SI D SE
M1 N_25 D GND GND mn15  l=0.13u w=0.28u m=1
M2 N_25 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M3 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M4 N_26 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M5 N_26 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_6 N_2 N_9 GND mn15  l=0.13u w=0.31u m=1
M8 N_27 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_27 N_7 N_9 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_2 N_7 GND mn15  l=0.13u w=0.17u m=1
M11 N_13 N_9 N_11 GND mn15  l=0.13u w=0.18u m=1
M12 N_11 N_9 N_13 GND mn15  l=0.13u w=0.18u m=1
M13 N_12 N_7 N_13 GND mn15  l=0.13u w=0.4u m=1
M14 N_28 N_2 N_12 GND mn15  l=0.13u w=0.17u m=1
M15 N_12 N_19 N_11 GND mn15  l=0.13u w=0.28u m=1
M16 N_28 N_24 N_11 GND mn15  l=0.13u w=0.17u m=1
M17 GND RN N_19 GND mn15  l=0.13u w=0.18u m=1
M18 N_11 SN GND GND mn15  l=0.13u w=0.27u m=1
M19 N_11 SN GND GND mn15  l=0.13u w=0.19u m=1
M20 Q N_24 GND GND mn15  l=0.13u w=0.46u m=1
M21 QN N_12 GND GND mn15  l=0.13u w=0.46u m=1
M22 N_24 N_12 GND GND mn15  l=0.13u w=0.28u m=1
M23 N_115 D VDD VDD mp15  l=0.13u w=0.42u m=1
M24 N_115 SE N_6 VDD mp15  l=0.13u w=0.42u m=1
M25 N_4 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M26 N_116 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M27 N_116 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M28 VDD CK N_2 VDD mp15  l=0.13u w=0.51u m=1
M29 N_117 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 N_6 N_7 N_9 VDD mp15  l=0.13u w=0.48u m=1
M31 VDD N_2 N_7 VDD mp15  l=0.13u w=0.42u m=1
M32 N_117 N_2 N_9 VDD mp15  l=0.13u w=0.17u m=1
M33 N_13 N_9 N_37 VDD mp15  l=0.13u w=0.32u m=1
M34 N_13 N_9 N_37 VDD mp15  l=0.13u w=0.31u m=1
M35 N_12 N_7 N_118 VDD mp15  l=0.13u w=0.17u m=1
M36 N_118 N_24 N_37 VDD mp15  l=0.13u w=0.17u m=1
M37 N_13 N_2 N_12 VDD mp15  l=0.13u w=0.55u m=1
M38 N_37 N_19 VDD VDD mp15  l=0.13u w=0.35u m=1
M39 VDD N_19 N_37 VDD mp15  l=0.13u w=0.35u m=1
M40 N_19 RN VDD VDD mp15  l=0.13u w=0.28u m=1
M41 N_12 SN VDD VDD mp15  l=0.13u w=0.37u m=1
M42 Q N_24 VDD VDD mp15  l=0.13u w=0.69u m=1
M43 QN N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M44 N_24 N_12 VDD VDD mp15  l=0.13u w=0.41u m=1
.ends sdbrb1
* SPICE INPUT		Tue Jul 31 20:22:32 2018	sdbrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrb2
.subckt sdbrb2 VDD QN Q SE SN RN CK SI D GND
M1 GND SE N_3 GND mn15  l=0.13u w=0.24u m=1
M2 N_56 SE N_6 GND mn15  l=0.13u w=0.28u m=1
M3 N_5 CK GND GND mn15  l=0.13u w=0.28u m=1
M4 N_55 D GND GND mn15  l=0.13u w=0.21u m=1
M5 N_54 D GND GND mn15  l=0.13u w=0.21u m=1
M6 N_54 N_3 N_6 GND mn15  l=0.13u w=0.21u m=1
M7 N_6 N_3 N_55 GND mn15  l=0.13u w=0.21u m=1
M8 N_56 SI GND GND mn15  l=0.13u w=0.28u m=1
M9 N_6 N_5 N_11 GND mn15  l=0.13u w=0.37u m=1
M10 N_57 N_26 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_57 N_9 N_11 GND mn15  l=0.13u w=0.17u m=1
M12 GND N_5 N_9 GND mn15  l=0.13u w=0.17u m=1
M13 N_26 N_11 N_53 GND mn15  l=0.13u w=0.32u m=1
M14 N_26 N_11 N_53 GND mn15  l=0.13u w=0.32u m=1
M15 N_15 N_9 N_26 GND mn15  l=0.13u w=0.54u m=1
M16 N_58 N_5 N_15 GND mn15  l=0.13u w=0.17u m=1
M17 N_53 N_19 N_15 GND mn15  l=0.13u w=0.18u m=1
M18 N_15 N_19 N_53 GND mn15  l=0.13u w=0.19u m=1
M19 N_53 N_23 N_58 GND mn15  l=0.13u w=0.17u m=1
M20 N_19 RN GND GND mn15  l=0.13u w=0.28u m=1
M21 GND SN N_53 GND mn15  l=0.13u w=0.205u m=1
M22 N_53 SN GND GND mn15  l=0.13u w=0.33u m=1
M23 N_53 SN GND GND mn15  l=0.13u w=0.33u m=1
M24 GND N_15 N_23 GND mn15  l=0.13u w=0.37u m=1
M25 GND N_23 Q GND mn15  l=0.13u w=0.455u m=1
M26 Q N_23 GND GND mn15  l=0.13u w=0.455u m=1
M27 GND N_15 QN GND mn15  l=0.13u w=0.46u m=1
M28 GND N_15 QN GND mn15  l=0.13u w=0.46u m=1
M29 N_3 SE VDD VDD mp15  l=0.13u w=0.37u m=1
M30 N_35 N_3 N_6 VDD mp15  l=0.13u w=0.42u m=1
M31 N_34 SE N_6 VDD mp15  l=0.13u w=0.31u m=1
M32 N_33 SE N_6 VDD mp15  l=0.13u w=0.31u m=1
M33 N_5 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M34 N_34 D VDD VDD mp15  l=0.13u w=0.31u m=1
M35 N_33 D VDD VDD mp15  l=0.13u w=0.31u m=1
M36 N_35 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M37 N_36 N_26 VDD VDD mp15  l=0.13u w=0.17u m=1
M38 N_6 N_9 N_11 VDD mp15  l=0.13u w=0.55u m=1
M39 VDD N_5 N_9 VDD mp15  l=0.13u w=0.42u m=1
M40 N_36 N_5 N_11 VDD mp15  l=0.13u w=0.17u m=1
M41 N_37 N_9 N_15 VDD mp15  l=0.13u w=0.17u m=1
M42 N_14 N_19 VDD VDD mp15  l=0.13u w=0.59u m=1
M43 N_14 N_19 VDD VDD mp15  l=0.13u w=0.59u m=1
M44 N_14 N_23 N_37 VDD mp15  l=0.13u w=0.17u m=1
M45 N_19 RN VDD VDD mp15  l=0.13u w=0.42u m=1
M46 N_15 SN VDD VDD mp15  l=0.13u w=0.55u m=1
M47 N_23 N_15 VDD VDD mp15  l=0.13u w=0.55u m=1
M48 Q N_23 VDD VDD mp15  l=0.13u w=0.69u m=1
M49 Q N_23 VDD VDD mp15  l=0.13u w=0.69u m=1
M50 VDD N_15 QN VDD mp15  l=0.13u w=0.69u m=1
M51 VDD N_15 QN VDD mp15  l=0.13u w=0.69u m=1
M52 N_26 N_11 N_14 VDD mp15  l=0.13u w=0.28u m=1
M53 N_14 N_11 N_26 VDD mp15  l=0.13u w=0.28u m=1
M54 N_26 N_11 N_14 VDD mp15  l=0.13u w=0.28u m=1
M55 N_14 N_11 N_26 VDD mp15  l=0.13u w=0.28u m=1
M56 N_15 N_5 N_26 VDD mp15  l=0.13u w=0.5u m=1
M57 N_26 N_5 N_15 VDD mp15  l=0.13u w=0.5u m=1
.ends sdbrb2
* SPICE INPUT		Tue Jul 31 20:22:46 2018	sdbrbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrbm
.subckt sdbrbm VDD Q QN GND SN RN CK SI D SE
M1 N_111 D GND GND mn15  l=0.13u w=0.24u m=1
M2 N_111 N_5 N_6 GND mn15  l=0.13u w=0.24u m=1
M3 N_112 SE N_6 GND mn15  l=0.13u w=0.24u m=1
M4 GND SE N_5 GND mn15  l=0.13u w=0.18u m=1
M5 N_112 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND CK N_3 GND mn15  l=0.13u w=0.2u m=1
M7 N_6 N_3 N_9 GND mn15  l=0.13u w=0.28u m=1
M8 N_113 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_113 N_7 N_9 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_3 N_7 GND mn15  l=0.13u w=0.17u m=1
M11 N_37 N_9 N_12 GND mn15  l=0.13u w=0.18u m=1
M12 N_12 N_9 N_37 GND mn15  l=0.13u w=0.18u m=1
M13 N_14 N_7 N_12 GND mn15  l=0.13u w=0.37u m=1
M14 N_114 N_3 N_14 GND mn15  l=0.13u w=0.17u m=1
M15 N_37 N_21 N_14 GND mn15  l=0.13u w=0.22u m=1
M16 N_114 N_26 N_37 GND mn15  l=0.13u w=0.17u m=1
M17 GND RN N_21 GND mn15  l=0.13u w=0.17u m=1
M18 N_37 SN GND GND mn15  l=0.13u w=0.21u m=1
M19 N_37 SN GND GND mn15  l=0.13u w=0.21u m=1
M20 Q N_26 GND GND mn15  l=0.13u w=0.36u m=1
M21 QN N_14 GND GND mn15  l=0.13u w=0.36u m=1
M22 N_26 N_14 GND GND mn15  l=0.13u w=0.22u m=1
M23 N_27 D VDD VDD mp15  l=0.13u w=0.37u m=1
M24 N_28 N_5 N_6 VDD mp15  l=0.13u w=0.37u m=1
M25 N_5 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M26 N_27 SE N_6 VDD mp15  l=0.13u w=0.37u m=1
M27 N_28 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M28 N_3 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M29 N_29 N_12 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 N_6 N_7 N_9 VDD mp15  l=0.13u w=0.42u m=1
M31 VDD N_3 N_7 VDD mp15  l=0.13u w=0.42u m=1
M32 N_29 N_3 N_9 VDD mp15  l=0.13u w=0.17u m=1
M33 N_12 N_9 N_11 VDD mp15  l=0.13u w=0.28u m=1
M34 N_11 N_9 N_12 VDD mp15  l=0.13u w=0.28u m=1
M35 N_14 N_7 N_30 VDD mp15  l=0.13u w=0.17u m=1
M36 N_30 N_26 N_11 VDD mp15  l=0.13u w=0.17u m=1
M37 N_12 N_3 N_14 VDD mp15  l=0.13u w=0.55u m=1
M38 VDD N_21 N_11 VDD mp15  l=0.13u w=0.28u m=1
M39 VDD N_21 N_11 VDD mp15  l=0.13u w=0.28u m=1
M40 N_21 RN VDD VDD mp15  l=0.13u w=0.24u m=1
M41 N_14 SN VDD VDD mp15  l=0.13u w=0.31u m=1
M42 Q N_26 VDD VDD mp15  l=0.13u w=0.55u m=1
M43 QN N_14 VDD VDD mp15  l=0.13u w=0.55u m=1
M44 N_26 N_14 VDD VDD mp15  l=0.13u w=0.31u m=1
.ends sdbrbm
* SPICE INPUT		Tue Jul 31 20:22:59 2018	sdbrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq0
.subckt sdbrq0 GND Q SE D SI CK SN RN VDD
M1 N_23 SI GND GND mn15  l=0.13u w=0.18u m=1
M2 N_22 N_4 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 N_22 D GND GND mn15  l=0.13u w=0.18u m=1
M4 N_23 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M5 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.18u m=1
M7 N_24 N_7 N_10 GND mn15  l=0.13u w=0.17u m=1
M8 N_10 N_2 N_6 GND mn15  l=0.13u w=0.18u m=1
M9 N_24 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M10 GND N_2 N_7 GND mn15  l=0.13u w=0.17u m=1
M11 N_25 N_21 N_11 GND mn15  l=0.13u w=0.17u m=1
M12 N_14 N_7 N_13 GND mn15  l=0.13u w=0.28u m=1
M13 N_13 N_2 N_25 GND mn15  l=0.13u w=0.17u m=1
M14 N_14 N_10 N_11 GND mn15  l=0.13u w=0.28u m=1
M15 GND RN N_15 GND mn15  l=0.13u w=0.18u m=1
M16 N_11 SN GND GND mn15  l=0.13u w=0.28u m=1
M17 N_11 N_15 N_13 GND mn15  l=0.13u w=0.2u m=1
M18 Q N_21 GND GND mn15  l=0.13u w=0.26u m=1
M19 N_21 N_13 GND GND mn15  l=0.13u w=0.18u m=1
M20 Q N_21 VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_21 N_13 VDD VDD mp15  l=0.13u w=0.26u m=1
M22 N_44 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M23 N_44 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M24 N_43 D VDD VDD mp15  l=0.13u w=0.28u m=1
M25 N_6 SE N_43 VDD mp15  l=0.13u w=0.28u m=1
M26 N_4 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M27 N_2 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M28 VDD RN N_15 VDD mp15  l=0.13u w=0.26u m=1
M29 N_13 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M30 N_10 N_7 N_6 VDD mp15  l=0.13u w=0.28u m=1
M31 N_45 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_7 N_2 VDD VDD mp15  l=0.13u w=0.42u m=1
M33 N_45 N_2 N_10 VDD mp15  l=0.13u w=0.17u m=1
M34 N_46 N_21 N_37 VDD mp15  l=0.13u w=0.17u m=1
M35 N_46 N_7 N_13 VDD mp15  l=0.13u w=0.17u m=1
M36 N_13 N_2 N_14 VDD mp15  l=0.13u w=0.44u m=1
M37 N_37 N_15 VDD VDD mp15  l=0.13u w=0.47u m=1
M38 N_14 N_10 N_37 VDD mp15  l=0.13u w=0.26u m=1
M39 N_14 N_10 N_37 VDD mp15  l=0.13u w=0.19u m=1
.ends sdbrq0
* SPICE INPUT		Tue Jul 31 20:23:12 2018	sdbrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq1
.subckt sdbrq1 GND Q SI SE SN RN VDD D CK
M1 GND N_18 N_2 GND mn15  l=0.13u w=0.17u m=1
M2 N_23 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M3 N_23 N_2 N_5 GND mn15  l=0.13u w=0.17u m=1
M4 N_5 N_18 N_4 GND mn15  l=0.13u w=0.31u m=1
M5 GND RN N_6 GND mn15  l=0.13u w=0.18u m=1
M6 N_8 SN GND GND mn15  l=0.13u w=0.46u m=1
M7 Q N_11 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_11 N_12 GND GND mn15  l=0.13u w=0.28u m=1
M9 N_24 N_11 N_8 GND mn15  l=0.13u w=0.17u m=1
M10 N_24 N_18 N_12 GND mn15  l=0.13u w=0.17u m=1
M11 N_12 N_2 N_14 GND mn15  l=0.13u w=0.4u m=1
M12 N_8 N_5 N_14 GND mn15  l=0.13u w=0.185u m=1
M13 N_14 N_5 N_8 GND mn15  l=0.13u w=0.185u m=1
M14 N_8 N_6 N_12 GND mn15  l=0.13u w=0.28u m=1
M15 GND CK N_18 GND mn15  l=0.13u w=0.2u m=1
M16 N_26 SE N_4 GND mn15  l=0.13u w=0.18u m=1
M17 GND SE N_20 GND mn15  l=0.13u w=0.18u m=1
M18 N_25 N_20 N_4 GND mn15  l=0.13u w=0.28u m=1
M19 N_25 D GND GND mn15  l=0.13u w=0.28u m=1
M20 N_26 SI GND GND mn15  l=0.13u w=0.18u m=1
M21 N_18 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M22 N_103 SE N_4 VDD mp15  l=0.13u w=0.42u m=1
M23 N_20 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M24 N_103 D VDD VDD mp15  l=0.13u w=0.42u m=1
M25 N_104 N_20 N_4 VDD mp15  l=0.13u w=0.28u m=1
M26 N_104 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M27 N_2 N_18 VDD VDD mp15  l=0.13u w=0.42u m=1
M28 N_105 N_18 N_5 VDD mp15  l=0.13u w=0.17u m=1
M29 N_105 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 N_4 N_2 N_5 VDD mp15  l=0.13u w=0.48u m=1
M31 N_14 N_18 N_12 VDD mp15  l=0.13u w=0.55u m=1
M32 N_12 N_2 N_106 VDD mp15  l=0.13u w=0.17u m=1
M33 N_14 N_5 N_36 VDD mp15  l=0.13u w=0.315u m=1
M34 N_36 N_5 N_14 VDD mp15  l=0.13u w=0.315u m=1
M35 N_106 N_11 N_36 VDD mp15  l=0.13u w=0.17u m=1
M36 N_36 N_6 VDD VDD mp15  l=0.13u w=0.35u m=1
M37 VDD N_6 N_36 VDD mp15  l=0.13u w=0.35u m=1
M38 VDD RN N_6 VDD mp15  l=0.13u w=0.28u m=1
M39 N_12 SN VDD VDD mp15  l=0.13u w=0.37u m=1
M40 Q N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 N_11 N_12 VDD VDD mp15  l=0.13u w=0.41u m=1
.ends sdbrq1
* SPICE INPUT		Tue Jul 31 20:23:25 2018	sdbrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdbrq2
.subckt sdbrq2 GND Q SE D SI CK SN RN VDD
M1 GND SE N_2 GND mn15  l=0.13u w=0.24u m=1
M2 N_29 SI GND GND mn15  l=0.13u w=0.28u m=1
M3 N_29 SE N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_27 N_2 N_6 GND mn15  l=0.13u w=0.21u m=1
M5 N_5 CK GND GND mn15  l=0.13u w=0.28u m=1
M6 N_28 D GND GND mn15  l=0.13u w=0.21u m=1
M7 N_27 D GND GND mn15  l=0.13u w=0.21u m=1
M8 N_6 N_2 N_28 GND mn15  l=0.13u w=0.21u m=1
M9 GND N_5 N_9 GND mn15  l=0.13u w=0.17u m=1
M10 N_30 N_9 N_11 GND mn15  l=0.13u w=0.17u m=1
M11 N_30 N_24 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_6 N_5 N_11 GND mn15  l=0.13u w=0.37u m=1
M13 GND RN N_13 GND mn15  l=0.13u w=0.28u m=1
M14 N_16 SN GND GND mn15  l=0.13u w=0.435u m=1
M15 N_16 SN GND GND mn15  l=0.13u w=0.435u m=1
M16 GND N_21 N_19 GND mn15  l=0.13u w=0.37u m=1
M17 GND N_19 Q GND mn15  l=0.13u w=0.46u m=1
M18 GND N_19 Q GND mn15  l=0.13u w=0.46u m=1
M19 N_16 N_13 N_21 GND mn15  l=0.13u w=0.37u m=1
M20 N_31 N_5 N_21 GND mn15  l=0.13u w=0.17u m=1
M21 N_21 N_9 N_24 GND mn15  l=0.13u w=0.54u m=1
M22 N_24 N_11 N_16 GND mn15  l=0.13u w=0.325u m=1
M23 N_24 N_11 N_16 GND mn15  l=0.13u w=0.325u m=1
M24 N_31 N_19 N_16 GND mn15  l=0.13u w=0.17u m=1
M25 N_2 SE VDD VDD mp15  l=0.13u w=0.37u m=1
M26 N_133 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M27 N_132 SE N_6 VDD mp15  l=0.13u w=0.31u m=1
M28 N_131 SE N_6 VDD mp15  l=0.13u w=0.31u m=1
M29 N_133 N_2 N_6 VDD mp15  l=0.13u w=0.42u m=1
M30 VDD CK N_5 VDD mp15  l=0.13u w=0.69u m=1
M31 N_132 D VDD VDD mp15  l=0.13u w=0.31u m=1
M32 N_131 D VDD VDD mp15  l=0.13u w=0.31u m=1
M33 N_21 N_5 N_24 VDD mp15  l=0.13u w=0.5u m=1
M34 N_24 N_5 N_21 VDD mp15  l=0.13u w=0.5u m=1
M35 N_24 N_11 N_45 VDD mp15  l=0.13u w=0.28u m=1
M36 N_24 N_11 N_45 VDD mp15  l=0.13u w=0.28u m=1
M37 N_24 N_11 N_45 VDD mp15  l=0.13u w=0.28u m=1
M38 N_24 N_11 N_45 VDD mp15  l=0.13u w=0.28u m=1
M39 N_45 N_13 VDD VDD mp15  l=0.13u w=0.58u m=1
M40 N_45 N_13 VDD VDD mp15  l=0.13u w=0.58u m=1
M41 N_134 N_9 N_21 VDD mp15  l=0.13u w=0.17u m=1
M42 N_45 N_19 N_134 VDD mp15  l=0.13u w=0.17u m=1
M43 N_13 RN VDD VDD mp15  l=0.13u w=0.42u m=1
M44 N_21 SN VDD VDD mp15  l=0.13u w=0.53u m=1
M45 N_19 N_21 VDD VDD mp15  l=0.13u w=0.55u m=1
M46 VDD N_19 Q VDD mp15  l=0.13u w=0.69u m=1
M47 VDD N_19 Q VDD mp15  l=0.13u w=0.69u m=1
M48 N_9 N_5 VDD VDD mp15  l=0.13u w=0.42u m=1
M49 N_135 N_5 N_11 VDD mp15  l=0.13u w=0.17u m=1
M50 N_6 N_9 N_11 VDD mp15  l=0.13u w=0.55u m=1
M51 N_135 N_24 VDD VDD mp15  l=0.13u w=0.17u m=1
.ends sdbrq2
* SPICE INPUT		Tue Jul 31 20:23:39 2018	sdcfb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb0
.subckt sdcfb0 VDD QN Q D SI CKN RN SE GND
M1 QN N_16 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 N_16 GND GND mn15  l=0.13u w=0.18u m=1
M3 N_7 RN GND GND mn15  l=0.13u w=0.17u m=1
M4 Q N_4 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_37 D GND GND mn15  l=0.13u w=0.26u m=1
M6 N_37 N_11 N_12 GND mn15  l=0.13u w=0.26u m=1
M7 N_38 SE N_12 GND mn15  l=0.13u w=0.18u m=1
M8 GND SE N_11 GND mn15  l=0.13u w=0.18u m=1
M9 GND CKN N_9 GND mn15  l=0.13u w=0.18u m=1
M10 N_38 SI GND GND mn15  l=0.13u w=0.18u m=1
M11 N_39 N_18 N_16 GND mn15  l=0.13u w=0.16u m=1
M12 N_16 N_9 N_15 GND mn15  l=0.13u w=0.23u m=1
M13 GND N_7 N_16 GND mn15  l=0.13u w=0.17u m=1
M14 GND N_4 N_39 GND mn15  l=0.13u w=0.16u m=1
M15 N_19 N_18 N_12 GND mn15  l=0.13u w=0.18u m=1
M16 GND N_9 N_18 GND mn15  l=0.13u w=0.17u m=1
M17 N_40 N_9 N_19 GND mn15  l=0.13u w=0.17u m=1
M18 N_40 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M19 N_15 N_19 GND GND mn15  l=0.13u w=0.23u m=1
M20 QN N_16 VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_4 N_16 VDD VDD mp15  l=0.13u w=0.26u m=1
M22 N_7 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M23 Q N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M24 N_23 D VDD VDD mp15  l=0.13u w=0.37u m=1
M25 N_24 N_11 N_12 VDD mp15  l=0.13u w=0.28u m=1
M26 N_23 SE N_12 VDD mp15  l=0.13u w=0.37u m=1
M27 N_11 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M28 N_9 CKN VDD VDD mp15  l=0.13u w=0.46u m=1
M29 N_24 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M30 N_16 N_18 N_15 VDD mp15  l=0.13u w=0.44u m=1
M31 N_15 N_19 N_13 VDD mp15  l=0.13u w=0.39u m=1
M32 N_16 N_9 N_25 VDD mp15  l=0.13u w=0.17u m=1
M33 N_25 N_4 N_13 VDD mp15  l=0.13u w=0.17u m=1
M34 N_26 N_18 N_19 VDD mp15  l=0.13u w=0.17u m=1
M35 N_18 N_9 VDD VDD mp15  l=0.13u w=0.42u m=1
M36 N_12 N_9 N_19 VDD mp15  l=0.13u w=0.5u m=1
M37 N_26 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M38 N_13 N_7 VDD VDD mp15  l=0.13u w=0.59u m=1
.ends sdcfb0
* SPICE INPUT		Tue Jul 31 20:23:51 2018	sdcfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb1
.subckt sdcfb1 VDD QN Q RN GND CKN SI D SE
M1 QN N_9 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_17 N_9 GND GND mn15  l=0.13u w=0.27u m=1
M3 N_37 D GND GND mn15  l=0.13u w=0.28u m=1
M4 N_37 N_5 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_38 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M6 GND SE N_5 GND mn15  l=0.13u w=0.18u m=1
M7 N_38 SI GND GND mn15  l=0.13u w=0.18u m=1
M8 GND CKN N_3 GND mn15  l=0.13u w=0.2u m=1
M9 GND N_17 Q GND mn15  l=0.13u w=0.45u m=1
M10 N_22 RN GND GND mn15  l=0.13u w=0.17u m=1
M11 GND N_3 N_12 GND mn15  l=0.13u w=0.2u m=1
M12 N_39 N_3 N_13 GND mn15  l=0.13u w=0.17u m=1
M13 N_39 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M14 N_13 N_12 N_6 GND mn15  l=0.13u w=0.28u m=1
M15 N_10 N_13 GND GND mn15  l=0.13u w=0.33u m=1
M16 GND N_22 N_9 GND mn15  l=0.13u w=0.28u m=1
M17 GND N_17 N_40 GND mn15  l=0.13u w=0.17u m=1
M18 N_10 N_3 N_9 GND mn15  l=0.13u w=0.41u m=1
M19 N_40 N_12 N_9 GND mn15  l=0.13u w=0.17u m=1
M20 N_23 D VDD VDD mp15  l=0.13u w=0.42u m=1
M21 N_24 N_5 N_6 VDD mp15  l=0.13u w=0.28u m=1
M22 N_23 SE N_6 VDD mp15  l=0.13u w=0.42u m=1
M23 N_5 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M24 N_24 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M25 N_3 CKN VDD VDD mp15  l=0.13u w=0.51u m=1
M26 N_25 N_17 N_7 VDD mp15  l=0.13u w=0.17u m=1
M27 N_25 N_3 N_9 VDD mp15  l=0.13u w=0.17u m=1
M28 N_10 N_12 N_9 VDD mp15  l=0.13u w=0.65u m=1
M29 N_10 N_13 N_7 VDD mp15  l=0.13u w=0.65u m=1
M30 N_12 N_3 VDD VDD mp15  l=0.13u w=0.51u m=1
M31 N_6 N_3 N_13 VDD mp15  l=0.13u w=0.42u m=1
M32 N_26 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M33 N_26 N_12 N_13 VDD mp15  l=0.13u w=0.17u m=1
M34 QN N_9 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 N_17 N_9 VDD VDD mp15  l=0.13u w=0.39u m=1
M36 N_7 N_22 VDD VDD mp15  l=0.13u w=0.69u m=1
M37 Q N_17 VDD VDD mp15  l=0.13u w=0.67u m=1
M38 N_22 RN VDD VDD mp15  l=0.13u w=0.28u m=1
.ends sdcfb1
* SPICE INPUT		Tue Jul 31 20:24:05 2018	sdcfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcfb2
.subckt sdcfb2 GND Q QN D VDD SE SI RN CKN
M1 N_27 D GND GND mn15  l=0.13u w=0.37u m=1
M2 N_27 N_4 N_6 GND mn15  l=0.13u w=0.37u m=1
M3 N_28 SE N_6 GND mn15  l=0.13u w=0.28u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.24u m=1
M5 N_28 SI GND GND mn15  l=0.13u w=0.28u m=1
M6 GND CKN N_2 GND mn15  l=0.13u w=0.27u m=1
M7 N_10 N_7 N_6 GND mn15  l=0.13u w=0.36u m=1
M8 N_29 N_11 GND GND mn15  l=0.13u w=0.17u m=1
M9 GND N_2 N_7 GND mn15  l=0.13u w=0.22u m=1
M10 N_29 N_2 N_10 GND mn15  l=0.13u w=0.17u m=1
M11 GND N_10 N_11 GND mn15  l=0.13u w=0.325u m=1
M12 N_11 N_10 GND GND mn15  l=0.13u w=0.325u m=1
M13 N_14 N_2 N_11 GND mn15  l=0.13u w=0.46u m=1
M14 GND N_21 N_14 GND mn15  l=0.13u w=0.37u m=1
M15 N_30 N_7 N_14 GND mn15  l=0.13u w=0.17u m=1
M16 GND N_25 N_30 GND mn15  l=0.13u w=0.17u m=1
M17 GND RN N_21 GND mn15  l=0.13u w=0.14u m=1
M18 N_21 RN GND GND mn15  l=0.13u w=0.14u m=1
M19 Q N_25 GND GND mn15  l=0.13u w=0.44u m=1
M20 GND N_25 Q GND mn15  l=0.13u w=0.44u m=1
M21 GND N_14 QN GND mn15  l=0.13u w=0.46u m=1
M22 GND N_14 QN GND mn15  l=0.13u w=0.46u m=1
M23 GND N_14 N_25 GND mn15  l=0.13u w=0.37u m=1
M24 N_46 D VDD VDD mp15  l=0.13u w=0.53u m=1
M25 N_6 N_4 N_42 VDD mp15  l=0.13u w=0.42u m=1
M26 N_46 SE N_6 VDD mp15  l=0.13u w=0.53u m=1
M27 N_4 SE VDD VDD mp15  l=0.13u w=0.37u m=1
M28 N_42 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M29 N_2 CKN VDD VDD mp15  l=0.13u w=0.67u m=1
M30 N_47 N_7 N_10 VDD mp15  l=0.13u w=0.17u m=1
M31 N_47 N_11 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_7 N_2 VDD VDD mp15  l=0.13u w=0.55u m=1
M33 N_6 N_2 N_10 VDD mp15  l=0.13u w=0.54u m=1
M34 N_11 N_10 N_40 VDD mp15  l=0.13u w=0.69u m=1
M35 N_40 N_10 N_11 VDD mp15  l=0.13u w=0.275u m=1
M36 N_11 N_10 N_40 VDD mp15  l=0.13u w=0.275u m=1
M37 N_48 N_2 N_14 VDD mp15  l=0.13u w=0.17u m=1
M38 N_11 N_7 N_14 VDD mp15  l=0.13u w=0.69u m=1
M39 N_48 N_25 N_40 VDD mp15  l=0.13u w=0.17u m=1
M40 N_40 N_21 VDD VDD mp15  l=0.13u w=0.625u m=1
M41 VDD N_21 N_40 VDD mp15  l=0.13u w=0.625u m=1
M42 VDD RN N_21 VDD mp15  l=0.13u w=0.42u m=1
M43 Q N_25 VDD VDD mp15  l=0.13u w=0.68u m=1
M44 VDD N_25 Q VDD mp15  l=0.13u w=0.68u m=1
M45 VDD N_14 QN VDD mp15  l=0.13u w=0.69u m=1
M46 VDD N_14 QN VDD mp15  l=0.13u w=0.69u m=1
M47 N_25 N_14 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends sdcfb2
* SPICE INPUT		Tue Jul 31 20:24:18 2018	sdcrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb0
.subckt sdcrb0 GND Q QN VDD SE CK RN SI D
M1 N_22 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_22 N_4 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 N_23 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M5 N_23 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.18u m=1
M7 N_24 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_24 N_7 N_10 GND mn15  l=0.13u w=0.17u m=1
M9 N_10 N_2 N_6 GND mn15  l=0.13u w=0.18u m=1
M10 GND N_2 N_7 GND mn15  l=0.13u w=0.17u m=1
M11 N_14 N_10 GND GND mn15  l=0.13u w=0.24u m=1
M12 N_11 N_7 N_14 GND mn15  l=0.13u w=0.22u m=1
M13 N_25 N_2 N_11 GND mn15  l=0.13u w=0.17u m=1
M14 GND N_18 N_11 GND mn15  l=0.13u w=0.18u m=1
M15 N_25 N_21 GND GND mn15  l=0.13u w=0.17u m=1
M16 N_18 RN GND GND mn15  l=0.13u w=0.18u m=1
M17 Q N_21 GND GND mn15  l=0.13u w=0.26u m=1
M18 QN N_11 GND GND mn15  l=0.13u w=0.26u m=1
M19 N_21 N_11 GND GND mn15  l=0.13u w=0.18u m=1
M20 N_104 D VDD VDD mp15  l=0.13u w=0.28u m=1
M21 N_6 SE N_104 VDD mp15  l=0.13u w=0.28u m=1
M22 N_4 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M23 N_105 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M24 N_105 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M25 N_2 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M26 N_106 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_10 N_7 N_6 VDD mp15  l=0.13u w=0.5u m=1
M28 VDD N_2 N_7 VDD mp15  l=0.13u w=0.42u m=1
M29 N_106 N_2 N_10 VDD mp15  l=0.13u w=0.17u m=1
M30 N_14 N_10 N_34 VDD mp15  l=0.13u w=0.19u m=1
M31 N_14 N_10 N_34 VDD mp15  l=0.13u w=0.26u m=1
M32 N_11 N_7 N_107 VDD mp15  l=0.13u w=0.17u m=1
M33 N_107 N_21 N_34 VDD mp15  l=0.13u w=0.17u m=1
M34 N_11 N_2 N_14 VDD mp15  l=0.13u w=0.42u m=1
M35 N_34 N_18 VDD VDD mp15  l=0.13u w=0.305u m=1
M36 VDD N_18 N_34 VDD mp15  l=0.13u w=0.305u m=1
M37 N_18 RN VDD VDD mp15  l=0.13u w=0.26u m=1
M38 Q N_21 VDD VDD mp15  l=0.13u w=0.4u m=1
M39 QN N_11 VDD VDD mp15  l=0.13u w=0.4u m=1
M40 N_21 N_11 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends sdcrb0
* SPICE INPUT		Tue Jul 31 20:24:31 2018	sdcrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb1
.subckt sdcrb1 GND QN Q RN CK SI D SE VDD
M1 N_23 D GND GND mn15  l=0.13u w=0.24u m=1
M2 N_23 N_4 N_6 GND mn15  l=0.13u w=0.24u m=1
M3 N_24 SE N_6 GND mn15  l=0.13u w=0.24u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.17u m=1
M5 N_24 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_25 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_25 N_7 N_10 GND mn15  l=0.13u w=0.17u m=1
M9 N_10 N_2 N_6 GND mn15  l=0.13u w=0.24u m=1
M10 GND N_2 N_7 GND mn15  l=0.13u w=0.17u m=1
M11 N_13 N_10 GND GND mn15  l=0.13u w=0.14u m=1
M12 GND N_10 N_13 GND mn15  l=0.13u w=0.14u m=1
M13 N_12 N_7 N_13 GND mn15  l=0.13u w=0.28u m=1
M14 N_26 N_2 N_12 GND mn15  l=0.13u w=0.17u m=1
M15 N_12 N_22 GND GND mn15  l=0.13u w=0.28u m=1
M16 N_26 N_19 GND GND mn15  l=0.13u w=0.17u m=1
M17 QN N_12 GND GND mn15  l=0.13u w=0.46u m=1
M18 N_19 N_12 GND GND mn15  l=0.13u w=0.28u m=1
M19 N_22 RN GND GND mn15  l=0.13u w=0.19u m=1
M20 Q N_19 GND GND mn15  l=0.13u w=0.43u m=1
M21 N_105 D VDD VDD mp15  l=0.13u w=0.37u m=1
M22 N_6 SE N_105 VDD mp15  l=0.13u w=0.37u m=1
M23 VDD SE N_4 VDD mp15  l=0.13u w=0.24u m=1
M24 N_106 N_4 N_6 VDD mp15  l=0.13u w=0.37u m=1
M25 N_106 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M26 N_2 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M27 N_107 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 N_6 N_7 N_10 VDD mp15  l=0.13u w=0.37u m=1
M29 N_7 N_2 VDD VDD mp15  l=0.13u w=0.42u m=1
M30 N_107 N_2 N_10 VDD mp15  l=0.13u w=0.17u m=1
M31 N_13 N_10 N_33 VDD mp15  l=0.13u w=0.35u m=1
M32 N_33 N_10 N_13 VDD mp15  l=0.13u w=0.35u m=1
M33 N_12 N_7 N_108 VDD mp15  l=0.13u w=0.17u m=1
M34 N_108 N_19 N_33 VDD mp15  l=0.13u w=0.17u m=1
M35 N_12 N_2 N_13 VDD mp15  l=0.13u w=0.42u m=1
M36 N_19 N_12 VDD VDD mp15  l=0.13u w=0.41u m=1
M37 QN N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M38 N_33 N_22 VDD VDD mp15  l=0.13u w=0.35u m=1
M39 N_33 N_22 VDD VDD mp15  l=0.13u w=0.35u m=1
M40 N_22 RN VDD VDD mp15  l=0.13u w=0.29u m=1
M41 Q N_19 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends sdcrb1
* SPICE INPUT		Tue Jul 31 20:24:44 2018	sdcrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrb2
.subckt sdcrb2 GND QN Q SE RN CK SI VDD D
M1 N_20 D GND GND mn15  l=0.13u w=0.24u m=1
M2 N_20 N_4 N_6 GND mn15  l=0.13u w=0.24u m=1
M3 N_21 SE N_6 GND mn15  l=0.13u w=0.24u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.17u m=1
M5 N_21 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.23u m=1
M7 N_23 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_24 N_8 N_10 GND mn15  l=0.13u w=0.17u m=1
M9 N_24 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M10 N_13 N_8 N_12 GND mn15  l=0.13u w=0.37u m=1
M11 N_25 N_10 N_12 GND mn15  l=0.13u w=0.39u m=1
M12 GND N_2 N_8 GND mn15  l=0.13u w=0.18u m=1
M13 N_26 N_2 N_13 GND mn15  l=0.13u w=0.17u m=1
M14 N_23 N_2 N_10 GND mn15  l=0.13u w=0.28u m=1
M15 N_26 N_16 N_22 GND mn15  l=0.13u w=0.17u m=1
M16 N_25 RN GND GND mn15  l=0.13u w=0.39u m=1
M17 N_22 RN GND GND mn15  l=0.13u w=0.17u m=1
M18 GND N_13 Q GND mn15  l=0.13u w=0.46u m=1
M19 Q N_13 GND GND mn15  l=0.13u w=0.46u m=1
M20 GND N_13 N_16 GND mn15  l=0.13u w=0.37u m=1
M21 GND N_16 QN GND mn15  l=0.13u w=0.46u m=1
M22 GND N_16 QN GND mn15  l=0.13u w=0.46u m=1
M23 N_45 D VDD VDD mp15  l=0.13u w=0.37u m=1
M24 N_46 N_4 N_6 VDD mp15  l=0.13u w=0.37u m=1
M25 N_6 SE N_45 VDD mp15  l=0.13u w=0.37u m=1
M26 VDD SE N_4 VDD mp15  l=0.13u w=0.24u m=1
M27 N_46 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M28 N_2 CK VDD VDD mp15  l=0.13u w=0.57u m=1
M29 N_47 N_6 VDD VDD mp15  l=0.13u w=0.39u m=1
M30 N_47 N_8 N_10 VDD mp15  l=0.13u w=0.39u m=1
M31 N_48 N_12 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_8 N_2 VDD VDD mp15  l=0.13u w=0.46u m=1
M33 N_48 N_2 N_10 VDD mp15  l=0.13u w=0.17u m=1
M34 N_12 RN VDD VDD mp15  l=0.13u w=0.23u m=1
M35 N_12 RN VDD VDD mp15  l=0.13u w=0.23u m=1
M36 N_12 N_10 VDD VDD mp15  l=0.13u w=0.23u m=1
M37 VDD N_10 N_12 VDD mp15  l=0.13u w=0.23u m=1
M38 N_13 N_2 N_12 VDD mp15  l=0.13u w=0.55u m=1
M39 N_49 N_8 N_13 VDD mp15  l=0.13u w=0.28u m=1
M40 N_49 N_16 VDD VDD mp15  l=0.13u w=0.28u m=1
M41 N_13 RN VDD VDD mp15  l=0.13u w=0.56u m=1
M42 Q N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M43 Q N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M44 N_16 N_13 VDD VDD mp15  l=0.13u w=0.55u m=1
M45 VDD N_16 QN VDD mp15  l=0.13u w=0.69u m=1
M46 VDD N_16 QN VDD mp15  l=0.13u w=0.69u m=1
.ends sdcrb2
* SPICE INPUT		Tue Jul 31 20:24:57 2018	sdcrbm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrbm
.subckt sdcrbm GND Q QN RN VDD CK SI D SE
M1 N_23 D GND GND mn15  l=0.13u w=0.24u m=1
M2 N_23 N_4 N_6 GND mn15  l=0.13u w=0.24u m=1
M3 N_24 SE N_6 GND mn15  l=0.13u w=0.24u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M5 N_24 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_25 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_25 N_7 N_10 GND mn15  l=0.13u w=0.17u m=1
M9 N_10 N_2 N_6 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_2 N_7 GND mn15  l=0.13u w=0.17u m=1
M11 N_13 N_10 GND GND mn15  l=0.13u w=0.14u m=1
M12 GND N_10 N_13 GND mn15  l=0.13u w=0.14u m=1
M13 N_11 N_7 N_13 GND mn15  l=0.13u w=0.28u m=1
M14 N_26 N_2 N_11 GND mn15  l=0.13u w=0.17u m=1
M15 GND N_19 N_11 GND mn15  l=0.13u w=0.22u m=1
M16 N_26 N_22 GND GND mn15  l=0.13u w=0.17u m=1
M17 N_19 RN GND GND mn15  l=0.13u w=0.17u m=1
M18 Q N_22 GND GND mn15  l=0.13u w=0.36u m=1
M19 QN N_11 GND GND mn15  l=0.13u w=0.36u m=1
M20 N_22 N_11 GND GND mn15  l=0.13u w=0.22u m=1
M21 N_43 D VDD VDD mp15  l=0.13u w=0.37u m=1
M22 N_6 SE N_43 VDD mp15  l=0.13u w=0.37u m=1
M23 N_4 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M24 N_44 N_4 N_6 VDD mp15  l=0.13u w=0.37u m=1
M25 N_44 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M26 N_2 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M27 N_45 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 N_6 N_7 N_10 VDD mp15  l=0.13u w=0.5u m=1
M29 VDD N_2 N_7 VDD mp15  l=0.13u w=0.42u m=1
M30 N_45 N_2 N_10 VDD mp15  l=0.13u w=0.17u m=1
M31 N_13 N_10 N_34 VDD mp15  l=0.13u w=0.29u m=1
M32 N_34 N_10 N_13 VDD mp15  l=0.13u w=0.29u m=1
M33 N_11 N_7 N_46 VDD mp15  l=0.13u w=0.17u m=1
M34 N_46 N_22 N_34 VDD mp15  l=0.13u w=0.17u m=1
M35 N_11 N_2 N_13 VDD mp15  l=0.13u w=0.42u m=1
M36 N_22 N_11 VDD VDD mp15  l=0.13u w=0.31u m=1
M37 QN N_11 VDD VDD mp15  l=0.13u w=0.55u m=1
M38 N_34 N_19 VDD VDD mp15  l=0.13u w=0.28u m=1
M39 N_34 N_19 VDD VDD mp15  l=0.13u w=0.28u m=1
M40 N_19 RN VDD VDD mp15  l=0.13u w=0.24u m=1
M41 Q N_22 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends sdcrbm
* SPICE INPUT		Tue Jul 31 20:25:09 2018	sdcrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq0
.subckt sdcrq0 GND Q SE D SI CK RN VDD
M1 N_19 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_19 N_4 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 N_20 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M5 N_20 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.18u m=1
M7 N_22 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_21 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_10 N_8 N_21 GND mn15  l=0.13u w=0.17u m=1
M10 N_22 N_2 N_10 GND mn15  l=0.13u w=0.28u m=1
M11 GND N_2 N_8 GND mn15  l=0.13u w=0.17u m=1
M12 N_11 N_10 N_13 GND mn15  l=0.13u w=0.3u m=1
M13 N_15 N_8 N_13 GND mn15  l=0.13u w=0.29u m=1
M14 N_23 N_2 N_15 GND mn15  l=0.13u w=0.17u m=1
M15 N_23 N_18 N_11 GND mn15  l=0.13u w=0.17u m=1
M16 GND RN N_11 GND mn15  l=0.13u w=0.46u m=1
M17 Q N_15 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_18 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M19 N_41 D VDD VDD mp15  l=0.13u w=0.28u m=1
M20 N_6 SE N_41 VDD mp15  l=0.13u w=0.28u m=1
M21 N_4 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M22 N_42 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M23 N_42 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M24 N_2 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M25 N_44 N_6 VDD VDD mp15  l=0.13u w=0.39u m=1
M26 N_44 N_8 N_10 VDD mp15  l=0.13u w=0.39u m=1
M27 N_43 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 VDD N_2 N_8 VDD mp15  l=0.13u w=0.42u m=1
M29 N_10 N_2 N_43 VDD mp15  l=0.13u w=0.17u m=1
M30 Q N_15 VDD VDD mp15  l=0.13u w=0.4u m=1
M31 N_18 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_13 N_10 VDD VDD mp15  l=0.13u w=0.19u m=1
M33 VDD N_10 N_13 VDD mp15  l=0.13u w=0.18u m=1
M34 N_15 N_2 N_13 VDD mp15  l=0.13u w=0.35u m=1
M35 N_45 N_8 N_15 VDD mp15  l=0.13u w=0.17u m=1
M36 N_45 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M37 VDD RN N_15 VDD mp15  l=0.13u w=0.21u m=1
.ends sdcrq0
* SPICE INPUT		Tue Jul 31 20:25:22 2018	sdcrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq1
.subckt sdcrq1 GND Q SE D SI CK RN VDD
M1 N_19 D GND GND mn15  l=0.13u w=0.28u m=1
M2 N_19 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M3 N_20 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M5 N_20 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_22 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_21 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_10 N_8 N_21 GND mn15  l=0.13u w=0.17u m=1
M10 N_22 N_2 N_10 GND mn15  l=0.13u w=0.28u m=1
M11 GND N_2 N_8 GND mn15  l=0.13u w=0.2u m=1
M12 N_11 N_10 N_13 GND mn15  l=0.13u w=0.37u m=1
M13 N_15 N_8 N_13 GND mn15  l=0.13u w=0.34u m=1
M14 N_23 N_2 N_15 GND mn15  l=0.13u w=0.17u m=1
M15 N_23 N_18 N_11 GND mn15  l=0.13u w=0.17u m=1
M16 GND RN N_11 GND mn15  l=0.13u w=0.46u m=1
M17 Q N_15 GND GND mn15  l=0.13u w=0.46u m=1
M18 N_18 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M19 N_41 D VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_41 SE N_6 VDD mp15  l=0.13u w=0.42u m=1
M21 N_4 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M22 N_42 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M23 N_42 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M24 VDD CK N_2 VDD mp15  l=0.13u w=0.51u m=1
M25 N_44 N_6 VDD VDD mp15  l=0.13u w=0.42u m=1
M26 N_44 N_8 N_10 VDD mp15  l=0.13u w=0.42u m=1
M27 N_43 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M28 VDD N_2 N_8 VDD mp15  l=0.13u w=0.51u m=1
M29 N_10 N_2 N_43 VDD mp15  l=0.13u w=0.17u m=1
M30 Q N_15 VDD VDD mp15  l=0.13u w=0.69u m=1
M31 N_18 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M32 N_13 N_10 VDD VDD mp15  l=0.13u w=0.19u m=1
M33 VDD N_10 N_13 VDD mp15  l=0.13u w=0.2u m=1
M34 N_15 N_2 N_13 VDD mp15  l=0.13u w=0.52u m=1
M35 N_45 N_8 N_15 VDD mp15  l=0.13u w=0.17u m=1
M36 N_45 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M37 VDD RN N_15 VDD mp15  l=0.13u w=0.39u m=1
.ends sdcrq1
* SPICE INPUT		Tue Jul 31 20:25:35 2018	sdcrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrq2
.subckt sdcrq2 GND Q SE D SI CK RN VDD
M1 N_20 D GND GND mn15  l=0.13u w=0.28u m=1
M2 N_6 N_4 N_20 GND mn15  l=0.13u w=0.28u m=1
M3 N_21 SE N_6 GND mn15  l=0.13u w=0.28u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M5 N_21 SI GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 CK GND GND mn15  l=0.13u w=0.28u m=1
M7 N_23 N_6 GND GND mn15  l=0.13u w=0.3u m=1
M8 N_22 N_13 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_10 N_8 N_22 GND mn15  l=0.13u w=0.17u m=1
M10 N_23 N_3 N_10 GND mn15  l=0.13u w=0.3u m=1
M11 GND N_3 N_8 GND mn15  l=0.13u w=0.2u m=1
M12 N_11 N_10 N_13 GND mn15  l=0.13u w=0.42u m=1
M13 N_15 N_8 N_13 GND mn15  l=0.13u w=0.37u m=1
M14 N_24 N_3 N_15 GND mn15  l=0.13u w=0.17u m=1
M15 N_24 N_18 N_11 GND mn15  l=0.13u w=0.17u m=1
M16 GND RN N_11 GND mn15  l=0.13u w=0.46u m=1
M17 GND N_15 Q GND mn15  l=0.13u w=0.46u m=1
M18 GND N_15 Q GND mn15  l=0.13u w=0.46u m=1
M19 GND N_15 N_18 GND mn15  l=0.13u w=0.17u m=1
M20 N_42 D VDD VDD mp15  l=0.13u w=0.42u m=1
M21 N_42 SE N_6 VDD mp15  l=0.13u w=0.42u m=1
M22 N_4 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M23 N_43 N_4 N_6 VDD mp15  l=0.13u w=0.42u m=1
M24 N_43 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M25 N_3 CK VDD VDD mp15  l=0.13u w=0.7u m=1
M26 N_44 N_6 VDD VDD mp15  l=0.13u w=0.46u m=1
M27 N_44 N_8 N_10 VDD mp15  l=0.13u w=0.46u m=1
M28 N_45 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_13 N_10 VDD VDD mp15  l=0.13u w=0.18u m=1
M30 VDD N_10 N_13 VDD mp15  l=0.13u w=0.18u m=1
M31 N_13 N_10 VDD VDD mp15  l=0.13u w=0.18u m=1
M32 N_15 N_3 N_13 VDD mp15  l=0.13u w=0.55u m=1
M33 VDD N_3 N_8 VDD mp15  l=0.13u w=0.51u m=1
M34 N_45 N_3 N_10 VDD mp15  l=0.13u w=0.17u m=1
M35 N_46 N_8 N_15 VDD mp15  l=0.13u w=0.17u m=1
M36 N_46 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M37 N_15 RN VDD VDD mp15  l=0.13u w=0.47u m=1
M38 VDD N_15 Q VDD mp15  l=0.13u w=0.69u m=1
M39 VDD N_15 Q VDD mp15  l=0.13u w=0.69u m=1
M40 VDD N_15 N_18 VDD mp15  l=0.13u w=0.17u m=1
.ends sdcrq2
* SPICE INPUT		Tue Jul 31 20:25:48 2018	sdcrqm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdcrqm
.subckt sdcrqm GND Q SI D SE CK RN VDD
M1 N_19 D GND GND mn15  l=0.13u w=0.24u m=1
M2 N_19 N_4 N_6 GND mn15  l=0.13u w=0.24u m=1
M3 N_20 SE N_6 GND mn15  l=0.13u w=0.24u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M5 N_20 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_21 N_2 N_11 GND mn15  l=0.13u w=0.17u m=1
M8 N_7 N_18 N_9 GND mn15  l=0.13u w=0.35u m=1
M9 N_11 N_16 N_9 GND mn15  l=0.13u w=0.27u m=1
M10 N_21 N_14 N_7 GND mn15  l=0.13u w=0.17u m=1
M11 GND RN N_7 GND mn15  l=0.13u w=0.42u m=1
M12 Q N_11 GND GND mn15  l=0.13u w=0.32u m=1
M13 N_14 N_11 GND GND mn15  l=0.13u w=0.17u m=1
M14 N_23 N_2 N_18 GND mn15  l=0.13u w=0.28u m=1
M15 GND N_2 N_16 GND mn15  l=0.13u w=0.17u m=1
M16 N_22 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M17 N_18 N_16 N_22 GND mn15  l=0.13u w=0.17u m=1
M18 N_23 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M19 N_41 D VDD VDD mp15  l=0.13u w=0.37u m=1
M20 N_6 SE N_41 VDD mp15  l=0.13u w=0.37u m=1
M21 N_4 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M22 N_42 N_4 N_6 VDD mp15  l=0.13u w=0.37u m=1
M23 N_42 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M24 N_2 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M25 N_11 N_2 N_9 VDD mp15  l=0.13u w=0.4u m=1
M26 N_9 N_18 VDD VDD mp15  l=0.13u w=0.21u m=1
M27 VDD N_18 N_9 VDD mp15  l=0.13u w=0.21u m=1
M28 N_43 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_43 N_16 N_11 VDD mp15  l=0.13u w=0.17u m=1
M30 VDD RN N_11 VDD mp15  l=0.13u w=0.31u m=1
M31 Q N_11 VDD VDD mp15  l=0.13u w=0.48u m=1
M32 N_14 N_11 VDD VDD mp15  l=0.13u w=0.17u m=1
M33 N_45 N_16 N_18 VDD mp15  l=0.13u w=0.42u m=1
M34 VDD N_2 N_16 VDD mp15  l=0.13u w=0.42u m=1
M35 N_18 N_2 N_44 VDD mp15  l=0.13u w=0.17u m=1
M36 N_44 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M37 N_45 N_6 VDD VDD mp15  l=0.13u w=0.42u m=1
.ends sdcrqm
* SPICE INPUT		Tue Jul 31 20:26:01 2018	sdmnrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdmnrq0
.subckt sdmnrq0 VDD Q GND CK SI SE D0 D1 S0
M1 N_43 D1 GND GND mn15  l=0.13u w=0.18u m=1
M2 GND S0 N_5 GND mn15  l=0.13u w=0.18u m=1
M3 N_43 S0 N_6 GND mn15  l=0.13u w=0.18u m=1
M4 N_44 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M5 N_44 D0 GND GND mn15  l=0.13u w=0.18u m=1
M6 GND SE N_3 GND mn15  l=0.13u w=0.18u m=1
M7 N_6 N_3 N_9 GND mn15  l=0.13u w=0.28u m=1
M8 N_45 SE N_9 GND mn15  l=0.13u w=0.24u m=1
M9 GND SI N_45 GND mn15  l=0.13u w=0.24u m=1
M10 N_46 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M11 N_47 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_14 N_12 GND GND mn15  l=0.13u w=0.14u m=1
M13 N_14 N_12 GND GND mn15  l=0.13u w=0.14u m=1
M14 N_47 N_8 N_12 GND mn15  l=0.13u w=0.17u m=1
M15 N_12 N_20 N_46 GND mn15  l=0.13u w=0.28u m=1
M16 GND N_20 N_8 GND mn15  l=0.13u w=0.17u m=1
M17 N_14 N_8 N_16 GND mn15  l=0.13u w=0.28u m=1
M18 N_48 N_20 N_16 GND mn15  l=0.13u w=0.17u m=1
M19 N_48 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M20 GND N_16 N_15 GND mn15  l=0.13u w=0.18u m=1
M21 Q N_16 GND GND mn15  l=0.13u w=0.26u m=1
M22 GND CK N_20 GND mn15  l=0.13u w=0.17u m=1
M23 N_22 D1 VDD VDD mp15  l=0.13u w=0.28u m=1
M24 N_6 N_5 N_22 VDD mp15  l=0.13u w=0.28u m=1
M25 N_23 S0 N_6 VDD mp15  l=0.13u w=0.28u m=1
M26 N_5 S0 VDD VDD mp15  l=0.13u w=0.26u m=1
M27 N_23 D0 VDD VDD mp15  l=0.13u w=0.28u m=1
M28 N_3 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M29 N_24 N_3 N_9 VDD mp15  l=0.13u w=0.37u m=1
M30 N_6 SE N_9 VDD mp15  l=0.13u w=0.42u m=1
M31 VDD SI N_24 VDD mp15  l=0.13u w=0.37u m=1
M32 N_25 N_9 VDD VDD mp15  l=0.13u w=0.42u m=1
M33 N_25 N_8 N_12 VDD mp15  l=0.13u w=0.42u m=1
M34 VDD N_14 N_26 VDD mp15  l=0.13u w=0.17u m=1
M35 N_14 N_12 VDD VDD mp15  l=0.13u w=0.21u m=1
M36 N_14 N_12 VDD VDD mp15  l=0.13u w=0.21u m=1
M37 N_8 N_20 VDD VDD mp15  l=0.13u w=0.42u m=1
M38 N_26 N_20 N_12 VDD mp15  l=0.13u w=0.17u m=1
M39 N_27 N_8 N_16 VDD mp15  l=0.13u w=0.17u m=1
M40 N_27 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M41 N_14 N_20 N_16 VDD mp15  l=0.13u w=0.42u m=1
M42 VDD N_16 N_15 VDD mp15  l=0.13u w=0.26u m=1
M43 Q N_16 VDD VDD mp15  l=0.13u w=0.4u m=1
M44 N_20 CK VDD VDD mp15  l=0.13u w=0.42u m=1
.ends sdmnrq0
* SPICE INPUT		Tue Jul 31 20:26:14 2018	sdmnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdmnrq1
.subckt sdmnrq1 VDD Q GND CK SI SE D0 D1 S0
M1 N_43 D1 GND GND mn15  l=0.13u w=0.27u m=1
M2 N_43 S0 N_6 GND mn15  l=0.13u w=0.27u m=1
M3 GND S0 N_4 GND mn15  l=0.13u w=0.16u m=1
M4 N_44 N_4 N_6 GND mn15  l=0.13u w=0.27u m=1
M5 N_44 D0 GND GND mn15  l=0.13u w=0.27u m=1
M6 GND SE N_3 GND mn15  l=0.13u w=0.17u m=1
M7 N_6 N_3 N_9 GND mn15  l=0.13u w=0.27u m=1
M8 N_45 SE N_9 GND mn15  l=0.13u w=0.23u m=1
M9 GND SI N_45 GND mn15  l=0.13u w=0.23u m=1
M10 N_46 N_9 GND GND mn15  l=0.13u w=0.27u m=1
M11 N_47 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_14 N_12 GND GND mn15  l=0.13u w=0.18u m=1
M13 N_14 N_12 GND GND mn15  l=0.13u w=0.18u m=1
M14 N_47 N_8 N_12 GND mn15  l=0.13u w=0.17u m=1
M15 N_12 N_20 N_46 GND mn15  l=0.13u w=0.27u m=1
M16 GND N_20 N_8 GND mn15  l=0.13u w=0.19u m=1
M17 N_14 N_8 N_16 GND mn15  l=0.13u w=0.36u m=1
M18 N_48 N_20 N_16 GND mn15  l=0.13u w=0.17u m=1
M19 N_48 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M20 N_15 N_16 GND GND mn15  l=0.13u w=0.27u m=1
M21 Q N_16 GND GND mn15  l=0.13u w=0.46u m=1
M22 GND CK N_20 GND mn15  l=0.13u w=0.19u m=1
M23 N_22 D1 VDD VDD mp15  l=0.13u w=0.4u m=1
M24 N_22 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M25 N_23 S0 N_6 VDD mp15  l=0.13u w=0.39u m=1
M26 VDD S0 N_4 VDD mp15  l=0.13u w=0.22u m=1
M27 N_23 D0 VDD VDD mp15  l=0.13u w=0.39u m=1
M28 N_3 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M29 N_24 N_3 N_9 VDD mp15  l=0.13u w=0.35u m=1
M30 N_6 SE N_9 VDD mp15  l=0.13u w=0.4u m=1
M31 VDD SI N_24 VDD mp15  l=0.13u w=0.35u m=1
M32 N_25 N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M33 N_25 N_8 N_12 VDD mp15  l=0.13u w=0.4u m=1
M34 VDD N_14 N_26 VDD mp15  l=0.13u w=0.17u m=1
M35 N_14 N_12 VDD VDD mp15  l=0.13u w=0.26u m=1
M36 N_14 N_12 VDD VDD mp15  l=0.13u w=0.26u m=1
M37 N_8 N_20 VDD VDD mp15  l=0.13u w=0.49u m=1
M38 N_26 N_20 N_12 VDD mp15  l=0.13u w=0.17u m=1
M39 N_27 N_8 N_16 VDD mp15  l=0.13u w=0.17u m=1
M40 N_27 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M41 N_14 N_20 N_16 VDD mp15  l=0.13u w=0.52u m=1
M42 VDD N_16 N_15 VDD mp15  l=0.13u w=0.33u m=1
M43 Q N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M44 N_20 CK VDD VDD mp15  l=0.13u w=0.49u m=1
.ends sdmnrq1
* SPICE INPUT		Tue Jul 31 20:26:26 2018	sdmnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdmnrq2
.subckt sdmnrq2 GND Q VDD CK SI SE D1 S0 D0
M1 GND S0 N_3 GND mn15  l=0.13u w=0.23u m=1
M2 N_23 D0 GND GND mn15  l=0.13u w=0.27u m=1
M3 N_5 N_3 N_23 GND mn15  l=0.13u w=0.27u m=1
M4 N_5 S0 N_22 GND mn15  l=0.13u w=0.27u m=1
M5 N_22 D1 GND GND mn15  l=0.13u w=0.27u m=1
M6 N_5 N_6 N_8 GND mn15  l=0.13u w=0.41u m=1
M7 N_24 SE N_8 GND mn15  l=0.13u w=0.27u m=1
M8 GND SE N_6 GND mn15  l=0.13u w=0.23u m=1
M9 N_24 SI GND GND mn15  l=0.13u w=0.27u m=1
M10 N_12 CK GND GND mn15  l=0.13u w=0.27u m=1
M11 N_25 N_8 GND GND mn15  l=0.13u w=0.41u m=1
M12 N_25 N_12 N_13 GND mn15  l=0.13u w=0.41u m=1
M13 N_26 N_10 N_13 GND mn15  l=0.13u w=0.17u m=1
M14 GND N_15 N_26 GND mn15  l=0.13u w=0.17u m=1
M15 N_15 N_13 GND GND mn15  l=0.13u w=0.41u m=1
M16 N_16 N_10 N_15 GND mn15  l=0.13u w=0.41u m=1
M17 N_27 N_20 GND GND mn15  l=0.13u w=0.17u m=1
M18 N_27 N_12 N_16 GND mn15  l=0.13u w=0.17u m=1
M19 GND N_12 N_10 GND mn15  l=0.13u w=0.22u m=1
M20 GND N_16 Q GND mn15  l=0.13u w=0.46u m=1
M21 GND N_16 Q GND mn15  l=0.13u w=0.46u m=1
M22 GND N_16 N_20 GND mn15  l=0.13u w=0.37u m=1
M23 VDD S0 N_3 VDD mp15  l=0.13u w=0.35u m=1
M24 N_48 D0 VDD VDD mp15  l=0.13u w=0.4u m=1
M25 N_5 S0 N_48 VDD mp15  l=0.13u w=0.4u m=1
M26 N_5 N_3 N_47 VDD mp15  l=0.13u w=0.4u m=1
M27 N_47 D1 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_5 SE N_8 VDD mp15  l=0.13u w=0.63u m=1
M29 N_49 N_6 N_8 VDD mp15  l=0.13u w=0.4u m=1
M30 N_6 SE VDD VDD mp15  l=0.13u w=0.35u m=1
M31 N_49 SI VDD VDD mp15  l=0.13u w=0.4u m=1
M32 N_12 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M33 N_50 N_8 VDD VDD mp15  l=0.13u w=0.62u m=1
M34 N_51 N_12 N_13 VDD mp15  l=0.13u w=0.17u m=1
M35 N_50 N_10 N_13 VDD mp15  l=0.13u w=0.62u m=1
M36 N_51 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M37 N_15 N_13 VDD VDD mp15  l=0.13u w=0.31u m=1
M38 N_15 N_13 VDD VDD mp15  l=0.13u w=0.32u m=1
M39 N_52 N_10 N_16 VDD mp15  l=0.13u w=0.17u m=1
M40 N_52 N_20 VDD VDD mp15  l=0.13u w=0.17u m=1
M41 N_16 N_12 N_15 VDD mp15  l=0.13u w=0.63u m=1
M42 VDD N_12 N_10 VDD mp15  l=0.13u w=0.55u m=1
M43 VDD N_16 Q VDD mp15  l=0.13u w=0.69u m=1
M44 VDD N_16 Q VDD mp15  l=0.13u w=0.69u m=1
M45 N_20 N_16 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends sdmnrq2
* SPICE INPUT		Tue Jul 31 20:26:39 2018	sdnfb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb0
.subckt sdnfb0 VDD Q QN SE D SI CKN GND
M1 Q N_14 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_9 N_14 GND GND mn15  l=0.13u w=0.18u m=1
M3 QN N_9 GND GND mn15  l=0.13u w=0.26u m=1
M4 N_35 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_35 N_13 N_14 GND mn15  l=0.13u w=0.17u m=1
M6 N_14 N_3 N_34 GND mn15  l=0.13u w=0.18u m=1
M7 GND N_3 N_13 GND mn15  l=0.13u w=0.17u m=1
M8 N_34 N_15 GND GND mn15  l=0.13u w=0.18u m=1
M9 N_36 N_3 N_18 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_18 N_15 GND mn15  l=0.13u w=0.18u m=1
M11 N_36 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_18 N_13 N_6 GND mn15  l=0.13u w=0.18u m=1
M13 GND CKN N_3 GND mn15  l=0.13u w=0.17u m=1
M14 N_38 SI GND GND mn15  l=0.13u w=0.18u m=1
M15 N_38 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M16 GND SE N_5 GND mn15  l=0.13u w=0.18u m=1
M17 N_37 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M18 N_37 D GND GND mn15  l=0.13u w=0.18u m=1
M19 N_3 CKN VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_20 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M21 N_20 N_5 N_6 VDD mp15  l=0.13u w=0.28u m=1
M22 N_5 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M23 N_6 SE N_19 VDD mp15  l=0.13u w=0.28u m=1
M24 N_19 D VDD VDD mp15  l=0.13u w=0.28u m=1
M25 Q N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M26 N_9 N_14 VDD VDD mp15  l=0.13u w=0.26u m=1
M27 QN N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_22 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_13 N_3 VDD VDD mp15  l=0.13u w=0.42u m=1
M30 N_22 N_3 N_14 VDD mp15  l=0.13u w=0.17u m=1
M31 N_21 N_13 N_14 VDD mp15  l=0.13u w=0.27u m=1
M32 N_21 N_15 VDD VDD mp15  l=0.13u w=0.27u m=1
M33 N_18 N_3 N_6 VDD mp15  l=0.13u w=0.18u m=1
M34 VDD N_18 N_15 VDD mp15  l=0.13u w=0.26u m=1
M35 N_23 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M36 N_23 N_13 N_18 VDD mp15  l=0.13u w=0.17u m=1
.ends sdnfb0
* SPICE INPUT		Tue Jul 31 20:26:52 2018	sdnfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb1
.subckt sdnfb1 GND Q QN CKN SI D SE VDD
M1 Q N_18 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 N_18 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_19 D GND GND mn15  l=0.13u w=0.28u m=1
M4 N_19 N_7 N_9 GND mn15  l=0.13u w=0.28u m=1
M5 N_20 SE N_9 GND mn15  l=0.13u w=0.24u m=1
M6 GND SE N_7 GND mn15  l=0.13u w=0.18u m=1
M7 N_20 SI GND GND mn15  l=0.13u w=0.24u m=1
M8 GND CKN N_5 GND mn15  l=0.13u w=0.2u m=1
M9 N_21 N_5 N_13 GND mn15  l=0.13u w=0.17u m=1
M10 N_13 N_16 N_9 GND mn15  l=0.13u w=0.28u m=1
M11 N_21 N_11 GND GND mn15  l=0.13u w=0.17u m=1
M12 N_11 N_13 GND GND mn15  l=0.13u w=0.28u m=1
M13 GND N_5 N_16 GND mn15  l=0.13u w=0.17u m=1
M14 N_22 N_11 GND GND mn15  l=0.13u w=0.42u m=1
M15 N_22 N_5 N_18 GND mn15  l=0.13u w=0.42u m=1
M16 N_23 N_16 N_18 GND mn15  l=0.13u w=0.17u m=1
M17 QN N_4 GND GND mn15  l=0.13u w=0.46u m=1
M18 N_23 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M19 N_35 D VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_35 SE N_9 VDD mp15  l=0.13u w=0.42u m=1
M21 N_7 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M22 N_36 N_7 N_9 VDD mp15  l=0.13u w=0.37u m=1
M23 N_36 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M24 N_5 CKN VDD VDD mp15  l=0.13u w=0.51u m=1
M25 Q N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 N_4 N_18 VDD VDD mp15  l=0.13u w=0.41u m=1
M27 N_13 N_5 N_9 VDD mp15  l=0.13u w=0.39u m=1
M28 N_37 N_16 N_13 VDD mp15  l=0.13u w=0.17u m=1
M29 N_37 N_11 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 VDD N_13 N_11 VDD mp15  l=0.13u w=0.39u m=1
M31 VDD N_5 N_16 VDD mp15  l=0.13u w=0.42u m=1
M32 N_38 N_11 VDD VDD mp15  l=0.13u w=0.59u m=1
M33 N_38 N_16 N_18 VDD mp15  l=0.13u w=0.59u m=1
M34 N_39 N_5 N_18 VDD mp15  l=0.13u w=0.17u m=1
M35 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 N_39 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
.ends sdnfb1
* SPICE INPUT		Tue Jul 31 20:27:05 2018	sdnfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfb2
.subckt sdnfb2 Q GND QN VDD SE D SI CKN
M1 GND N_13 Q GND mn15  l=0.13u w=0.46u m=1
M2 GND N_13 Q GND mn15  l=0.13u w=0.46u m=1
M3 GND N_13 N_4 GND mn15  l=0.13u w=0.37u m=1
M4 N_23 N_9 N_10 GND mn15  l=0.13u w=0.37u m=1
M5 N_23 D GND GND mn15  l=0.13u w=0.37u m=1
M6 N_7 CKN GND GND mn15  l=0.13u w=0.28u m=1
M7 N_24 SE N_10 GND mn15  l=0.13u w=0.28u m=1
M8 N_9 SE GND GND mn15  l=0.13u w=0.28u m=1
M9 N_24 SI GND GND mn15  l=0.13u w=0.28u m=1
M10 GND N_4 QN GND mn15  l=0.13u w=0.46u m=1
M11 GND N_4 QN GND mn15  l=0.13u w=0.46u m=1
M12 GND N_4 N_27 GND mn15  l=0.13u w=0.17u m=1
M13 N_27 N_17 N_13 GND mn15  l=0.13u w=0.17u m=1
M14 N_26 N_7 N_13 GND mn15  l=0.13u w=0.32u m=1
M15 N_26 N_20 GND GND mn15  l=0.13u w=0.32u m=1
M16 N_25 N_20 GND GND mn15  l=0.13u w=0.32u m=1
M17 N_25 N_7 N_13 GND mn15  l=0.13u w=0.32u m=1
M18 GND N_7 N_17 GND mn15  l=0.13u w=0.23u m=1
M19 N_20 N_21 GND GND mn15  l=0.13u w=0.31u m=1
M20 N_28 N_20 GND GND mn15  l=0.13u w=0.17u m=1
M21 N_28 N_7 N_21 GND mn15  l=0.13u w=0.17u m=1
M22 N_10 N_17 N_21 GND mn15  l=0.13u w=0.37u m=1
M23 VDD N_13 Q VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_13 Q VDD mp15  l=0.13u w=0.69u m=1
M25 N_4 N_13 VDD VDD mp15  l=0.13u w=0.55u m=1
M26 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 VDD N_4 QN VDD mp15  l=0.13u w=0.69u m=1
M28 N_114 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_114 N_7 N_13 VDD mp15  l=0.13u w=0.17u m=1
M30 N_113 N_17 N_13 VDD mp15  l=0.13u w=0.49u m=1
M31 N_113 N_20 VDD VDD mp15  l=0.13u w=0.49u m=1
M32 VDD N_20 N_112 VDD mp15  l=0.13u w=0.49u m=1
M33 N_112 N_17 N_13 VDD mp15  l=0.13u w=0.49u m=1
M34 VDD N_21 N_20 VDD mp15  l=0.13u w=0.48u m=1
M35 N_115 N_20 VDD VDD mp15  l=0.13u w=0.17u m=1
M36 N_115 N_17 N_21 VDD mp15  l=0.13u w=0.17u m=1
M37 N_10 N_7 N_21 VDD mp15  l=0.13u w=0.55u m=1
M38 VDD N_7 N_17 VDD mp15  l=0.13u w=0.56u m=1
M39 N_116 D VDD VDD mp15  l=0.13u w=0.53u m=1
M40 N_7 CKN VDD VDD mp15  l=0.13u w=0.67u m=1
M41 N_9 SE VDD VDD mp15  l=0.13u w=0.39u m=1
M42 N_10 SE N_116 VDD mp15  l=0.13u w=0.53u m=1
M43 N_117 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M44 N_117 N_9 N_10 VDD mp15  l=0.13u w=0.42u m=1
.ends sdnfb2
* SPICE INPUT		Tue Jul 31 20:27:18 2018	sdnfq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfq0
.subckt sdnfq0 VDD Q GND CKN SI D SE
M1 N_33 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_33 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 N_34 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_5 GND mn15  l=0.13u w=0.18u m=1
M5 N_34 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CKN N_3 GND mn15  l=0.13u w=0.17u m=1
M7 N_35 N_3 N_10 GND mn15  l=0.13u w=0.17u m=1
M8 N_10 N_13 N_6 GND mn15  l=0.13u w=0.18u m=1
M9 N_35 N_8 GND GND mn15  l=0.13u w=0.17u m=1
M10 GND N_10 N_8 GND mn15  l=0.13u w=0.18u m=1
M11 GND N_3 N_13 GND mn15  l=0.13u w=0.17u m=1
M12 N_14 N_3 N_37 GND mn15  l=0.13u w=0.18u m=1
M13 N_14 N_13 N_36 GND mn15  l=0.13u w=0.17u m=1
M14 N_36 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M15 N_37 N_8 GND GND mn15  l=0.13u w=0.18u m=1
M16 Q N_14 GND GND mn15  l=0.13u w=0.26u m=1
M17 N_17 N_14 GND GND mn15  l=0.13u w=0.18u m=1
M18 N_18 D VDD VDD mp15  l=0.13u w=0.28u m=1
M19 N_19 N_5 N_6 VDD mp15  l=0.13u w=0.28u m=1
M20 N_6 SE N_18 VDD mp15  l=0.13u w=0.28u m=1
M21 N_5 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M22 N_19 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M23 N_3 CKN VDD VDD mp15  l=0.13u w=0.42u m=1
M24 N_10 N_3 N_6 VDD mp15  l=0.13u w=0.18u m=1
M25 N_20 N_13 N_10 VDD mp15  l=0.13u w=0.17u m=1
M26 N_20 N_8 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_8 N_10 VDD VDD mp15  l=0.13u w=0.26u m=1
M28 N_13 N_3 VDD VDD mp15  l=0.13u w=0.42u m=1
M29 N_14 N_3 N_21 VDD mp15  l=0.13u w=0.17u m=1
M30 N_21 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M31 N_22 N_8 VDD VDD mp15  l=0.13u w=0.27u m=1
M32 N_22 N_13 N_14 VDD mp15  l=0.13u w=0.27u m=1
M33 Q N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M34 N_17 N_14 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends sdnfq0
* SPICE INPUT		Tue Jul 31 20:27:32 2018	sdnfq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfq1
.subckt sdnfq1 VDD Q CKN SI GND SE D
M1 Q N_8 GND GND mn15  l=0.13u w=0.46u m=1
M2 N_4 N_8 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_34 N_11 N_12 GND mn15  l=0.13u w=0.28u m=1
M4 N_34 D GND GND mn15  l=0.13u w=0.28u m=1
M5 N_35 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND CKN N_9 GND mn15  l=0.13u w=0.2u m=1
M7 N_35 SE N_12 GND mn15  l=0.13u w=0.24u m=1
M8 GND SE N_11 GND mn15  l=0.13u w=0.18u m=1
M9 N_8 N_6 N_36 GND mn15  l=0.13u w=0.17u m=1
M10 N_36 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_37 N_9 N_8 GND mn15  l=0.13u w=0.41u m=1
M12 N_37 N_15 GND GND mn15  l=0.13u w=0.41u m=1
M13 GND N_9 N_6 GND mn15  l=0.13u w=0.17u m=1
M14 N_38 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M15 N_12 N_6 N_16 GND mn15  l=0.13u w=0.28u m=1
M16 N_15 N_16 GND GND mn15  l=0.13u w=0.28u m=1
M17 N_38 N_9 N_16 GND mn15  l=0.13u w=0.17u m=1
M18 Q N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_4 N_8 VDD VDD mp15  l=0.13u w=0.39u m=1
M20 N_18 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M21 N_8 N_9 N_18 VDD mp15  l=0.13u w=0.17u m=1
M22 N_19 N_15 VDD VDD mp15  l=0.13u w=0.57u m=1
M23 VDD N_9 N_6 VDD mp15  l=0.13u w=0.42u m=1
M24 N_19 N_6 N_8 VDD mp15  l=0.13u w=0.57u m=1
M25 N_20 D VDD VDD mp15  l=0.13u w=0.42u m=1
M26 N_21 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M27 VDD CKN N_9 VDD mp15  l=0.13u w=0.51u m=1
M28 N_20 SE N_12 VDD mp15  l=0.13u w=0.42u m=1
M29 N_11 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M30 N_21 N_11 N_12 VDD mp15  l=0.13u w=0.37u m=1
M31 N_12 N_9 N_16 VDD mp15  l=0.13u w=0.39u m=1
M32 N_22 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M33 N_22 N_6 N_16 VDD mp15  l=0.13u w=0.17u m=1
M34 N_15 N_16 VDD VDD mp15  l=0.13u w=0.39u m=1
.ends sdnfq1
* SPICE INPUT		Tue Jul 31 20:27:45 2018	sdnfq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnfq2
.subckt sdnfq2 GND Q VDD SI D CKN SE
M1 GND N_13 N_2 GND mn15  l=0.13u w=0.23u m=1
M2 N_5 N_6 GND GND mn15  l=0.13u w=0.32u m=1
M3 N_21 N_5 GND GND mn15  l=0.13u w=0.17u m=1
M4 N_21 N_13 N_6 GND mn15  l=0.13u w=0.17u m=1
M5 N_7 N_2 N_6 GND mn15  l=0.13u w=0.37u m=1
M6 GND N_18 Q GND mn15  l=0.13u w=0.46u m=1
M7 GND N_18 Q GND mn15  l=0.13u w=0.46u m=1
M8 GND N_18 N_10 GND mn15  l=0.13u w=0.37u m=1
M9 N_23 SI GND GND mn15  l=0.13u w=0.28u m=1
M10 N_13 CKN GND GND mn15  l=0.13u w=0.28u m=1
M11 N_22 D GND GND mn15  l=0.13u w=0.37u m=1
M12 N_23 SE N_7 GND mn15  l=0.13u w=0.28u m=1
M13 N_15 SE GND GND mn15  l=0.13u w=0.28u m=1
M14 N_22 N_15 N_7 GND mn15  l=0.13u w=0.37u m=1
M15 N_26 N_5 GND GND mn15  l=0.13u w=0.33u m=1
M16 N_25 N_5 GND GND mn15  l=0.13u w=0.33u m=1
M17 N_26 N_13 N_18 GND mn15  l=0.13u w=0.33u m=1
M18 N_18 N_2 N_24 GND mn15  l=0.13u w=0.17u m=1
M19 N_24 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M20 N_25 N_13 N_18 GND mn15  l=0.13u w=0.33u m=1
M21 VDD N_13 N_2 VDD mp15  l=0.13u w=0.58u m=1
M22 VDD N_18 Q VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_18 Q VDD mp15  l=0.13u w=0.69u m=1
M24 N_10 N_18 VDD VDD mp15  l=0.13u w=0.55u m=1
M25 N_47 N_5 VDD VDD mp15  l=0.13u w=0.51u m=1
M26 VDD N_5 N_46 VDD mp15  l=0.13u w=0.51u m=1
M27 N_47 N_2 N_18 VDD mp15  l=0.13u w=0.51u m=1
M28 N_18 N_13 N_45 VDD mp15  l=0.13u w=0.17u m=1
M29 N_45 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 N_46 N_2 N_18 VDD mp15  l=0.13u w=0.51u m=1
M31 N_49 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M32 N_13 CKN VDD VDD mp15  l=0.13u w=0.69u m=1
M33 N_48 D VDD VDD mp15  l=0.13u w=0.53u m=1
M34 N_15 SE VDD VDD mp15  l=0.13u w=0.39u m=1
M35 N_7 SE N_48 VDD mp15  l=0.13u w=0.53u m=1
M36 N_49 N_15 N_7 VDD mp15  l=0.13u w=0.42u m=1
M37 N_7 N_13 N_6 VDD mp15  l=0.13u w=0.55u m=1
M38 VDD N_6 N_5 VDD mp15  l=0.13u w=0.5u m=1
M39 N_50 N_5 VDD VDD mp15  l=0.13u w=0.17u m=1
M40 N_50 N_2 N_6 VDD mp15  l=0.13u w=0.17u m=1
.ends sdnfq2
* SPICE INPUT		Tue Jul 31 20:27:58 2018	sdnrb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb0
.subckt sdnrb0 GND QN Q VDD CK SI D SE
M1 N_19 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_19 N_4 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 N_20 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M5 N_20 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.17u m=1
M7 N_9 N_2 N_6 GND mn15  l=0.13u w=0.18u m=1
M8 N_21 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M9 GND N_9 N_7 GND mn15  l=0.13u w=0.18u m=1
M10 N_21 N_13 N_9 GND mn15  l=0.13u w=0.17u m=1
M11 GND N_2 N_13 GND mn15  l=0.13u w=0.17u m=1
M12 N_22 N_7 GND GND mn15  l=0.13u w=0.18u m=1
M13 N_15 N_13 N_22 GND mn15  l=0.13u w=0.18u m=1
M14 N_23 N_2 N_15 GND mn15  l=0.13u w=0.17u m=1
M15 QN N_18 GND GND mn15  l=0.13u w=0.26u m=1
M16 N_23 N_18 GND GND mn15  l=0.13u w=0.17u m=1
M17 Q N_15 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_18 N_15 GND GND mn15  l=0.13u w=0.18u m=1
M19 N_35 D VDD VDD mp15  l=0.13u w=0.28u m=1
M20 N_4 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M21 N_6 SE N_35 VDD mp15  l=0.13u w=0.28u m=1
M22 N_36 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M23 N_36 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M24 N_2 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M25 N_37 N_2 N_9 VDD mp15  l=0.13u w=0.17u m=1
M26 N_37 N_7 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 VDD N_9 N_7 VDD mp15  l=0.13u w=0.26u m=1
M28 N_9 N_13 N_6 VDD mp15  l=0.13u w=0.28u m=1
M29 VDD N_2 N_13 VDD mp15  l=0.13u w=0.42u m=1
M30 N_38 N_7 VDD VDD mp15  l=0.13u w=0.27u m=1
M31 N_39 N_13 N_15 VDD mp15  l=0.13u w=0.17u m=1
M32 N_38 N_2 N_15 VDD mp15  l=0.13u w=0.27u m=1
M33 QN N_18 VDD VDD mp15  l=0.13u w=0.4u m=1
M34 N_39 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M35 Q N_15 VDD VDD mp15  l=0.13u w=0.4u m=1
M36 N_18 N_15 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends sdnrb0
* SPICE INPUT		Tue Jul 31 20:28:11 2018	sdnrb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb1
.subckt sdnrb1 GND QN Q VDD SI CK D SE
M1 N_19 D GND GND mn15  l=0.13u w=0.28u m=1
M2 N_19 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M3 N_20 SE N_6 GND mn15  l=0.13u w=0.24u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.17u m=1
M5 N_20 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_9 N_2 N_6 GND mn15  l=0.13u w=0.24u m=1
M8 N_21 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M9 GND N_9 N_7 GND mn15  l=0.13u w=0.28u m=1
M10 N_21 N_13 N_9 GND mn15  l=0.13u w=0.17u m=1
M11 GND N_2 N_13 GND mn15  l=0.13u w=0.17u m=1
M12 N_22 N_7 GND GND mn15  l=0.13u w=0.37u m=1
M13 N_22 N_13 N_15 GND mn15  l=0.13u w=0.37u m=1
M14 N_23 N_2 N_15 GND mn15  l=0.13u w=0.17u m=1
M15 QN N_18 GND GND mn15  l=0.13u w=0.46u m=1
M16 N_23 N_18 GND GND mn15  l=0.13u w=0.17u m=1
M17 Q N_15 GND GND mn15  l=0.13u w=0.46u m=1
M18 N_18 N_15 GND GND mn15  l=0.13u w=0.28u m=1
M19 N_40 D VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_40 SE N_6 VDD mp15  l=0.13u w=0.42u m=1
M21 VDD SE N_4 VDD mp15  l=0.13u w=0.24u m=1
M22 N_41 N_4 N_6 VDD mp15  l=0.13u w=0.37u m=1
M23 N_41 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M24 N_2 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M25 N_42 N_2 N_9 VDD mp15  l=0.13u w=0.17u m=1
M26 N_42 N_7 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 VDD N_9 N_7 VDD mp15  l=0.13u w=0.39u m=1
M28 N_9 N_13 N_6 VDD mp15  l=0.13u w=0.37u m=1
M29 VDD N_2 N_13 VDD mp15  l=0.13u w=0.42u m=1
M30 N_43 N_7 VDD VDD mp15  l=0.13u w=0.55u m=1
M31 N_44 N_13 N_15 VDD mp15  l=0.13u w=0.17u m=1
M32 N_43 N_2 N_15 VDD mp15  l=0.13u w=0.55u m=1
M33 QN N_18 VDD VDD mp15  l=0.13u w=0.69u m=1
M34 N_44 N_18 VDD VDD mp15  l=0.13u w=0.17u m=1
M35 Q N_15 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 N_18 N_15 VDD VDD mp15  l=0.13u w=0.41u m=1
.ends sdnrb1
* SPICE INPUT		Tue Jul 31 20:28:23 2018	sdnrb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrb2
.subckt sdnrb2 Q GND QN SE D SI CK VDD
M1 GND N_8 Q GND mn15  l=0.13u w=0.46u m=1
M2 GND N_8 Q GND mn15  l=0.13u w=0.46u m=1
M3 GND N_8 N_4 GND mn15  l=0.13u w=0.37u m=1
M4 GND N_4 QN GND mn15  l=0.13u w=0.46u m=1
M5 GND N_4 QN GND mn15  l=0.13u w=0.46u m=1
M6 GND N_4 N_25 GND mn15  l=0.13u w=0.17u m=1
M7 N_25 N_19 N_8 GND mn15  l=0.13u w=0.17u m=1
M8 N_24 N_12 N_8 GND mn15  l=0.13u w=0.36u m=1
M9 N_24 N_17 GND GND mn15  l=0.13u w=0.36u m=1
M10 N_23 N_17 GND GND mn15  l=0.13u w=0.36u m=1
M11 N_23 N_12 N_8 GND mn15  l=0.13u w=0.36u m=1
M12 GND N_19 N_12 GND mn15  l=0.13u w=0.23u m=1
M13 N_26 N_12 N_14 GND mn15  l=0.13u w=0.17u m=1
M14 N_17 N_14 GND GND mn15  l=0.13u w=0.165u m=1
M15 N_17 N_14 GND GND mn15  l=0.13u w=0.155u m=1
M16 N_26 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M17 N_15 N_19 N_14 GND mn15  l=0.13u w=0.28u m=1
M18 N_19 CK GND GND mn15  l=0.13u w=0.28u m=1
M19 N_28 SI GND GND mn15  l=0.13u w=0.28u m=1
M20 N_28 SE N_15 GND mn15  l=0.13u w=0.28u m=1
M21 GND SE N_20 GND mn15  l=0.13u w=0.24u m=1
M22 N_15 N_20 N_27 GND mn15  l=0.13u w=0.28u m=1
M23 N_27 D GND GND mn15  l=0.13u w=0.28u m=1
M24 VDD N_8 Q VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_8 Q VDD mp15  l=0.13u w=0.69u m=1
M26 N_4 N_8 VDD VDD mp15  l=0.13u w=0.55u m=1
M27 VDD N_4 QN VDD mp15  l=0.13u w=0.69u m=1
M28 QN N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_4 N_49 VDD mp15  l=0.13u w=0.17u m=1
M30 N_47 N_19 N_8 VDD mp15  l=0.13u w=0.51u m=1
M31 N_48 N_19 N_8 VDD mp15  l=0.13u w=0.51u m=1
M32 N_49 N_12 N_8 VDD mp15  l=0.13u w=0.17u m=1
M33 N_48 N_17 VDD VDD mp15  l=0.13u w=0.51u m=1
M34 N_47 N_17 VDD VDD mp15  l=0.13u w=0.51u m=1
M35 N_12 N_19 VDD VDD mp15  l=0.13u w=0.56u m=1
M36 N_15 N_12 N_14 VDD mp15  l=0.13u w=0.42u m=1
M37 VDD N_14 N_17 VDD mp15  l=0.13u w=0.48u m=1
M38 N_50 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M39 N_50 N_19 N_14 VDD mp15  l=0.13u w=0.17u m=1
M40 N_19 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M41 N_52 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M42 N_52 N_20 N_15 VDD mp15  l=0.13u w=0.42u m=1
M43 N_15 SE N_51 VDD mp15  l=0.13u w=0.42u m=1
M44 N_20 SE VDD VDD mp15  l=0.13u w=0.37u m=1
M45 N_51 D VDD VDD mp15  l=0.13u w=0.42u m=1
.ends sdnrb2
* SPICE INPUT		Tue Jul 31 20:28:37 2018	sdnrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq0
.subckt sdnrq0 VDD Q GND SI D SE CK
M1 N_34 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_34 N_5 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 N_35 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_5 GND mn15  l=0.13u w=0.18u m=1
M5 N_35 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_3 GND mn15  l=0.13u w=0.17u m=1
M7 N_10 N_3 N_6 GND mn15  l=0.13u w=0.18u m=1
M8 N_36 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M9 GND N_10 N_7 GND mn15  l=0.13u w=0.18u m=1
M10 N_36 N_13 N_10 GND mn15  l=0.13u w=0.17u m=1
M11 Q N_14 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_17 N_14 GND GND mn15  l=0.13u w=0.18u m=1
M13 GND N_3 N_13 GND mn15  l=0.13u w=0.17u m=1
M14 N_38 N_7 GND GND mn15  l=0.13u w=0.18u m=1
M15 N_38 N_13 N_14 GND mn15  l=0.13u w=0.18u m=1
M16 N_14 N_3 N_37 GND mn15  l=0.13u w=0.17u m=1
M17 N_37 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M18 N_18 D VDD VDD mp15  l=0.13u w=0.28u m=1
M19 N_6 SE N_18 VDD mp15  l=0.13u w=0.28u m=1
M20 N_5 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M21 N_19 N_5 N_6 VDD mp15  l=0.13u w=0.28u m=1
M22 N_19 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M23 N_3 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M24 N_20 N_3 N_10 VDD mp15  l=0.13u w=0.17u m=1
M25 N_20 N_7 VDD VDD mp15  l=0.13u w=0.17u m=1
M26 VDD N_10 N_7 VDD mp15  l=0.13u w=0.26u m=1
M27 N_10 N_13 N_6 VDD mp15  l=0.13u w=0.28u m=1
M28 N_13 N_3 VDD VDD mp15  l=0.13u w=0.42u m=1
M29 N_22 N_7 VDD VDD mp15  l=0.13u w=0.27u m=1
M30 N_14 N_3 N_22 VDD mp15  l=0.13u w=0.27u m=1
M31 N_14 N_13 N_21 VDD mp15  l=0.13u w=0.17u m=1
M32 N_21 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M33 Q N_14 VDD VDD mp15  l=0.13u w=0.4u m=1
M34 N_17 N_14 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends sdnrq0
* SPICE INPUT		Tue Jul 31 20:28:50 2018	sdnrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq1
.subckt sdnrq1 GND Q SI D SE CK VDD
M1 N_5 N_6 N_18 GND mn15  l=0.13u w=0.17u m=1
M2 N_19 N_3 N_5 GND mn15  l=0.13u w=0.37u m=1
M3 GND N_6 N_3 GND mn15  l=0.13u w=0.17u m=1
M4 N_18 N_17 GND GND mn15  l=0.13u w=0.17u m=1
M5 N_19 N_11 GND GND mn15  l=0.13u w=0.37u m=1
M6 N_21 SI GND GND mn15  l=0.13u w=0.24u m=1
M7 N_21 SE N_10 GND mn15  l=0.13u w=0.24u m=1
M8 GND SE N_8 GND mn15  l=0.13u w=0.17u m=1
M9 N_20 D GND GND mn15  l=0.13u w=0.28u m=1
M10 N_20 N_8 N_10 GND mn15  l=0.13u w=0.28u m=1
M11 GND CK N_6 GND mn15  l=0.13u w=0.2u m=1
M12 N_13 N_6 N_10 GND mn15  l=0.13u w=0.24u m=1
M13 GND N_13 N_11 GND mn15  l=0.13u w=0.28u m=1
M14 N_22 N_3 N_13 GND mn15  l=0.13u w=0.17u m=1
M15 N_22 N_11 GND GND mn15  l=0.13u w=0.17u m=1
M16 Q N_5 GND GND mn15  l=0.13u w=0.46u m=1
M17 N_17 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M18 Q N_5 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_17 N_5 VDD VDD mp15  l=0.13u w=0.41u m=1
M20 N_40 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M21 N_40 N_8 N_10 VDD mp15  l=0.13u w=0.37u m=1
M22 N_10 SE N_39 VDD mp15  l=0.13u w=0.42u m=1
M23 VDD SE N_8 VDD mp15  l=0.13u w=0.24u m=1
M24 N_39 D VDD VDD mp15  l=0.13u w=0.42u m=1
M25 N_6 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M26 N_42 N_6 N_5 VDD mp15  l=0.13u w=0.55u m=1
M27 VDD N_6 N_3 VDD mp15  l=0.13u w=0.42u m=1
M28 N_41 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_42 N_11 VDD VDD mp15  l=0.13u w=0.55u m=1
M30 N_5 N_3 N_41 VDD mp15  l=0.13u w=0.17u m=1
M31 VDD N_13 N_11 VDD mp15  l=0.13u w=0.39u m=1
M32 N_43 N_6 N_13 VDD mp15  l=0.13u w=0.17u m=1
M33 N_13 N_3 N_10 VDD mp15  l=0.13u w=0.37u m=1
M34 N_43 N_11 VDD VDD mp15  l=0.13u w=0.17u m=1
.ends sdnrq1
* SPICE INPUT		Tue Jul 31 20:29:03 2018	sdnrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdnrq2
.subckt sdnrq2 GND Q CK SI D SE VDD
M1 Q N_4 GND GND mn15  l=0.13u w=0.46u m=1
M2 Q N_4 GND GND mn15  l=0.13u w=0.46u m=1
M3 N_3 N_4 GND GND mn15  l=0.13u w=0.37u m=1
M4 GND N_3 N_22 GND mn15  l=0.13u w=0.17u m=1
M5 N_22 N_16 N_4 GND mn15  l=0.13u w=0.17u m=1
M6 N_21 N_9 N_4 GND mn15  l=0.13u w=0.36u m=1
M7 N_21 N_14 GND GND mn15  l=0.13u w=0.36u m=1
M8 N_20 N_14 GND GND mn15  l=0.13u w=0.36u m=1
M9 N_20 N_9 N_4 GND mn15  l=0.13u w=0.36u m=1
M10 GND N_16 N_9 GND mn15  l=0.13u w=0.23u m=1
M11 N_23 N_9 N_12 GND mn15  l=0.13u w=0.17u m=1
M12 N_14 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M13 N_14 N_12 GND GND mn15  l=0.13u w=0.16u m=1
M14 N_23 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M15 N_12 N_16 N_11 GND mn15  l=0.13u w=0.28u m=1
M16 N_16 CK GND GND mn15  l=0.13u w=0.28u m=1
M17 N_25 SI GND GND mn15  l=0.13u w=0.28u m=1
M18 N_25 SE N_11 GND mn15  l=0.13u w=0.28u m=1
M19 GND SE N_17 GND mn15  l=0.13u w=0.24u m=1
M20 N_11 N_17 N_24 GND mn15  l=0.13u w=0.28u m=1
M21 N_24 D GND GND mn15  l=0.13u w=0.28u m=1
M22 N_9 N_16 VDD VDD mp15  l=0.13u w=0.58u m=1
M23 N_3 N_4 VDD VDD mp15  l=0.13u w=0.55u m=1
M24 Q N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 Q N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 VDD N_3 N_46 VDD mp15  l=0.13u w=0.17u m=1
M27 N_44 N_16 N_4 VDD mp15  l=0.13u w=0.51u m=1
M28 N_45 N_16 N_4 VDD mp15  l=0.13u w=0.51u m=1
M29 N_46 N_9 N_4 VDD mp15  l=0.13u w=0.17u m=1
M30 N_45 N_14 VDD VDD mp15  l=0.13u w=0.51u m=1
M31 N_44 N_14 VDD VDD mp15  l=0.13u w=0.51u m=1
M32 N_11 N_9 N_12 VDD mp15  l=0.13u w=0.42u m=1
M33 VDD N_12 N_14 VDD mp15  l=0.13u w=0.5u m=1
M34 N_47 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M35 N_47 N_16 N_12 VDD mp15  l=0.13u w=0.17u m=1
M36 N_16 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M37 N_49 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M38 N_49 N_17 N_11 VDD mp15  l=0.13u w=0.42u m=1
M39 N_17 SE VDD VDD mp15  l=0.13u w=0.37u m=1
M40 N_11 SE N_48 VDD mp15  l=0.13u w=0.42u m=1
M41 N_48 D VDD VDD mp15  l=0.13u w=0.42u m=1
.ends sdnrq2
* SPICE INPUT		Tue Jul 31 20:29:15 2018	sdpfb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb0
.subckt sdpfb0 GND QN Q VDD SN CKN SI D SE
M1 N_22 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_22 N_4 N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_23 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M5 N_23 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CKN N_2 GND mn15  l=0.13u w=0.18u m=1
M7 QN N_15 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_9 N_15 GND GND mn15  l=0.13u w=0.18u m=1
M9 N_13 N_10 N_6 GND mn15  l=0.13u w=0.18u m=1
M10 N_24 N_14 GND GND mn15  l=0.13u w=0.17u m=1
M11 GND N_2 N_10 GND mn15  l=0.13u w=0.17u m=1
M12 N_24 N_2 N_13 GND mn15  l=0.13u w=0.17u m=1
M13 N_16 N_13 N_14 GND mn15  l=0.13u w=0.29u m=1
M14 N_15 N_2 N_14 GND mn15  l=0.13u w=0.29u m=1
M15 N_25 N_10 N_15 GND mn15  l=0.13u w=0.17u m=1
M16 N_16 N_9 N_25 GND mn15  l=0.13u w=0.17u m=1
M17 N_16 SN GND GND mn15  l=0.13u w=0.31u m=1
M18 Q N_9 GND GND mn15  l=0.13u w=0.26u m=1
M19 QN N_15 VDD VDD mp15  l=0.13u w=0.4u m=1
M20 N_9 N_15 VDD VDD mp15  l=0.13u w=0.26u m=1
M21 N_41 D VDD VDD mp15  l=0.13u w=0.37u m=1
M22 N_42 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M23 N_41 SE N_6 VDD mp15  l=0.13u w=0.37u m=1
M24 N_4 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M25 N_42 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M26 VDD CKN N_2 VDD mp15  l=0.13u w=0.46u m=1
M27 N_43 N_10 N_13 VDD mp15  l=0.13u w=0.17u m=1
M28 N_43 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_6 N_2 N_13 VDD mp15  l=0.13u w=0.5u m=1
M30 VDD N_2 N_10 VDD mp15  l=0.13u w=0.42u m=1
M31 VDD N_13 N_14 VDD mp15  l=0.13u w=0.31u m=1
M32 N_15 N_2 N_44 VDD mp15  l=0.13u w=0.17u m=1
M33 N_15 N_10 N_14 VDD mp15  l=0.13u w=0.37u m=1
M34 N_44 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M35 N_15 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M36 Q N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends sdpfb0
* SPICE INPUT		Tue Jul 31 20:29:28 2018	sdpfb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb1
.subckt sdpfb1 GND Q QN VDD SN CKN SI D SE
M1 N_22 D GND GND mn15  l=0.13u w=0.27u m=1
M2 N_22 N_4 N_6 GND mn15  l=0.13u w=0.27u m=1
M3 GND SE N_4 GND mn15  l=0.13u w=0.17u m=1
M4 N_23 SE N_6 GND mn15  l=0.13u w=0.17u m=1
M5 N_23 SI GND GND mn15  l=0.13u w=0.17u m=1
M6 GND CKN N_2 GND mn15  l=0.13u w=0.19u m=1
M7 N_6 N_7 N_9 GND mn15  l=0.13u w=0.3u m=1
M8 N_24 N_11 GND GND mn15  l=0.13u w=0.16u m=1
M9 GND N_2 N_7 GND mn15  l=0.13u w=0.16u m=1
M10 N_24 N_2 N_9 GND mn15  l=0.13u w=0.16u m=1
M11 N_13 N_9 N_11 GND mn15  l=0.13u w=0.29u m=1
M12 N_12 N_2 N_11 GND mn15  l=0.13u w=0.4u m=1
M13 N_25 N_7 N_12 GND mn15  l=0.13u w=0.17u m=1
M14 N_13 N_21 N_25 GND mn15  l=0.13u w=0.17u m=1
M15 N_13 SN GND GND mn15  l=0.13u w=0.46u m=1
M16 Q N_21 GND GND mn15  l=0.13u w=0.46u m=1
M17 QN N_12 GND GND mn15  l=0.13u w=0.46u m=1
M18 N_21 N_12 GND GND mn15  l=0.13u w=0.27u m=1
M19 N_41 D VDD VDD mp15  l=0.13u w=0.4u m=1
M20 N_42 N_4 N_6 VDD mp15  l=0.13u w=0.26u m=1
M21 N_41 SE N_6 VDD mp15  l=0.13u w=0.4u m=1
M22 N_4 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M23 N_42 SI VDD VDD mp15  l=0.13u w=0.26u m=1
M24 VDD CKN N_2 VDD mp15  l=0.13u w=0.49u m=1
M25 N_43 N_7 N_9 VDD mp15  l=0.13u w=0.16u m=1
M26 N_43 N_11 VDD VDD mp15  l=0.13u w=0.16u m=1
M27 N_6 N_2 N_9 VDD mp15  l=0.13u w=0.48u m=1
M28 VDD N_2 N_7 VDD mp15  l=0.13u w=0.4u m=1
M29 VDD N_9 N_11 VDD mp15  l=0.13u w=0.31u m=1
M30 N_12 N_2 N_44 VDD mp15  l=0.13u w=0.17u m=1
M31 N_12 N_7 N_11 VDD mp15  l=0.13u w=0.57u m=1
M32 N_44 N_21 VDD VDD mp15  l=0.13u w=0.17u m=1
M33 N_12 SN VDD VDD mp15  l=0.13u w=0.35u m=1
M34 Q N_21 VDD VDD mp15  l=0.13u w=0.69u m=1
M35 QN N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 N_21 N_12 VDD VDD mp15  l=0.13u w=0.39u m=1
.ends sdpfb1
* SPICE INPUT		Tue Jul 31 20:29:41 2018	sdpfb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdpfb2
.subckt sdpfb2 Q GND QN VDD SN CKN SI D SE
M1 GND N_14 Q GND mn15  l=0.13u w=0.46u m=1
M2 GND N_14 Q GND mn15  l=0.13u w=0.46u m=1
M3 GND SN N_5 GND mn15  l=0.13u w=0.46u m=1
M4 N_5 SN GND GND mn15  l=0.13u w=0.46u m=1
M5 N_28 D GND GND mn15  l=0.13u w=0.37u m=1
M6 N_28 N_9 N_11 GND mn15  l=0.13u w=0.37u m=1
M7 N_29 SE N_11 GND mn15  l=0.13u w=0.28u m=1
M8 GND SE N_9 GND mn15  l=0.13u w=0.24u m=1
M9 N_29 SI GND GND mn15  l=0.13u w=0.28u m=1
M10 N_8 CKN GND GND mn15  l=0.13u w=0.27u m=1
M11 GND N_22 QN GND mn15  l=0.13u w=0.46u m=1
M12 GND N_22 QN GND mn15  l=0.13u w=0.46u m=1
M13 GND N_22 N_14 GND mn15  l=0.13u w=0.37u m=1
M14 N_11 N_16 N_18 GND mn15  l=0.13u w=0.3u m=1
M15 N_30 N_21 GND GND mn15  l=0.13u w=0.17u m=1
M16 GND N_8 N_16 GND mn15  l=0.13u w=0.22u m=1
M17 N_30 N_8 N_18 GND mn15  l=0.13u w=0.17u m=1
M18 N_31 N_14 N_5 GND mn15  l=0.13u w=0.17u m=1
M19 N_22 N_8 N_21 GND mn15  l=0.13u w=0.41u m=1
M20 N_22 N_8 N_21 GND mn15  l=0.13u w=0.41u m=1
M21 N_22 N_16 N_31 GND mn15  l=0.13u w=0.17u m=1
M22 N_5 N_18 N_21 GND mn15  l=0.13u w=0.27u m=1
M23 N_21 N_18 N_5 GND mn15  l=0.13u w=0.22u m=1
M24 N_5 N_18 N_21 GND mn15  l=0.13u w=0.2u m=1
M25 N_48 D VDD VDD mp15  l=0.13u w=0.53u m=1
M26 N_11 SE N_48 VDD mp15  l=0.13u w=0.53u m=1
M27 N_9 SE VDD VDD mp15  l=0.13u w=0.37u m=1
M28 N_49 N_9 N_11 VDD mp15  l=0.13u w=0.42u m=1
M29 N_49 SI VDD VDD mp15  l=0.13u w=0.42u m=1
M30 VDD CKN N_8 VDD mp15  l=0.13u w=0.67u m=1
M31 Q N_14 VDD VDD mp15  l=0.13u w=0.69u m=1
M32 VDD N_14 Q VDD mp15  l=0.13u w=0.69u m=1
M33 N_50 N_14 VDD VDD mp15  l=0.13u w=0.17u m=1
M34 N_22 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M35 N_22 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M36 N_50 N_8 N_22 VDD mp15  l=0.13u w=0.17u m=1
M37 N_51 N_16 N_18 VDD mp15  l=0.13u w=0.17u m=1
M38 N_51 N_21 VDD VDD mp15  l=0.13u w=0.17u m=1
M39 N_16 N_8 VDD VDD mp15  l=0.13u w=0.55u m=1
M40 N_11 N_8 N_18 VDD mp15  l=0.13u w=0.53u m=1
M41 VDD N_22 QN VDD mp15  l=0.13u w=0.69u m=1
M42 VDD N_22 QN VDD mp15  l=0.13u w=0.69u m=1
M43 N_14 N_22 VDD VDD mp15  l=0.13u w=0.55u m=1
M44 VDD N_18 N_21 VDD mp15  l=0.13u w=0.32u m=1
M45 VDD N_18 N_21 VDD mp15  l=0.13u w=0.32u m=1
M46 N_21 N_16 N_22 VDD mp15  l=0.13u w=0.56u m=1
M47 N_22 N_16 N_21 VDD mp15  l=0.13u w=0.44u m=1
.ends sdpfb2
* SPICE INPUT		Tue Jul 31 20:29:54 2018	sdprb0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb0
.subckt sdprb0 GND QN Q SN CK SI D SE VDD
M1 N_22 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_22 N_4 N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_23 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.17u m=1
M5 N_23 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 QN N_17 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_9 N_17 GND GND mn15  l=0.13u w=0.18u m=1
M9 N_6 N_2 N_12 GND mn15  l=0.13u w=0.26u m=1
M10 N_24 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_24 N_10 N_12 GND mn15  l=0.13u w=0.17u m=1
M12 GND N_2 N_10 GND mn15  l=0.13u w=0.17u m=1
M13 N_15 N_12 N_14 GND mn15  l=0.13u w=0.16u m=1
M14 N_14 N_12 N_15 GND mn15  l=0.13u w=0.15u m=1
M15 N_15 N_10 N_17 GND mn15  l=0.13u w=0.3u m=1
M16 N_17 N_2 N_25 GND mn15  l=0.13u w=0.17u m=1
M17 N_25 N_9 N_14 GND mn15  l=0.13u w=0.17u m=1
M18 N_14 SN GND GND mn15  l=0.13u w=0.31u m=1
M19 Q N_9 GND GND mn15  l=0.13u w=0.26u m=1
M20 N_42 D VDD VDD mp15  l=0.13u w=0.37u m=1
M21 N_43 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M22 N_6 SE N_42 VDD mp15  l=0.13u w=0.37u m=1
M23 N_4 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M24 N_43 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M25 N_2 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M26 N_44 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M27 N_6 N_10 N_12 VDD mp15  l=0.13u w=0.37u m=1
M28 VDD N_2 N_10 VDD mp15  l=0.13u w=0.42u m=1
M29 N_44 N_2 N_12 VDD mp15  l=0.13u w=0.17u m=1
M30 N_15 N_12 VDD VDD mp15  l=0.13u w=0.2u m=1
M31 VDD N_12 N_15 VDD mp15  l=0.13u w=0.19u m=1
M32 N_17 N_10 N_45 VDD mp15  l=0.13u w=0.17u m=1
M33 N_45 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M34 N_17 N_2 N_15 VDD mp15  l=0.13u w=0.39u m=1
M35 N_17 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M36 VDD N_9 Q VDD mp15  l=0.13u w=0.4u m=1
M37 QN N_17 VDD VDD mp15  l=0.13u w=0.4u m=1
M38 N_9 N_17 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends sdprb0
* SPICE INPUT		Tue Jul 31 20:30:07 2018	sdprb1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb1
.subckt sdprb1 VDD Q QN D SI CK SE SN GND
M1 N_40 N_13 N_37 GND mn15  l=0.13u w=0.17u m=1
M2 N_3 N_21 N_37 GND mn15  l=0.13u w=0.19u m=1
M3 N_37 N_21 N_3 GND mn15  l=0.13u w=0.17u m=1
M4 N_3 N_19 N_6 GND mn15  l=0.13u w=0.36u m=1
M5 N_6 N_15 N_40 GND mn15  l=0.13u w=0.17u m=1
M6 N_37 SN GND GND mn15  l=0.13u w=0.2u m=1
M7 N_37 SN GND GND mn15  l=0.13u w=0.18u m=1
M8 Q N_13 GND GND mn15  l=0.13u w=0.46u m=1
M9 GND CK N_15 GND mn15  l=0.13u w=0.2u m=1
M10 N_41 N_16 N_18 GND mn15  l=0.13u w=0.24u m=1
M11 N_41 D GND GND mn15  l=0.13u w=0.24u m=1
M12 N_42 SI GND GND mn15  l=0.13u w=0.18u m=1
M13 N_42 SE N_18 GND mn15  l=0.13u w=0.18u m=1
M14 GND SE N_16 GND mn15  l=0.13u w=0.17u m=1
M15 QN N_6 GND GND mn15  l=0.13u w=0.46u m=1
M16 N_13 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M17 N_43 N_3 GND GND mn15  l=0.13u w=0.17u m=1
M18 N_43 N_19 N_21 GND mn15  l=0.13u w=0.17u m=1
M19 N_21 N_15 N_18 GND mn15  l=0.13u w=0.24u m=1
M20 GND N_15 N_19 GND mn15  l=0.13u w=0.17u m=1
M21 N_3 N_21 VDD VDD mp15  l=0.13u w=0.21u m=1
M22 VDD N_21 N_3 VDD mp15  l=0.13u w=0.2u m=1
M23 N_23 N_13 VDD VDD mp15  l=0.13u w=0.17u m=1
M24 N_6 N_19 N_23 VDD mp15  l=0.13u w=0.17u m=1
M25 N_6 N_15 N_3 VDD mp15  l=0.13u w=0.5u m=1
M26 N_6 SN VDD VDD mp15  l=0.13u w=0.45u m=1
M27 Q N_13 VDD VDD mp15  l=0.13u w=0.35u m=1
M28 Q N_13 VDD VDD mp15  l=0.13u w=0.35u m=1
M29 QN N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M30 N_13 N_6 VDD VDD mp15  l=0.13u w=0.42u m=1
M31 N_15 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M32 N_25 N_16 N_18 VDD mp15  l=0.13u w=0.28u m=1
M33 N_24 D VDD VDD mp15  l=0.13u w=0.37u m=1
M34 N_25 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M35 N_18 SE N_24 VDD mp15  l=0.13u w=0.37u m=1
M36 VDD SE N_16 VDD mp15  l=0.13u w=0.24u m=1
M37 N_26 N_3 VDD VDD mp15  l=0.13u w=0.17u m=1
M38 N_18 N_19 N_21 VDD mp15  l=0.13u w=0.37u m=1
M39 VDD N_15 N_19 VDD mp15  l=0.13u w=0.42u m=1
M40 N_26 N_15 N_21 VDD mp15  l=0.13u w=0.17u m=1
.ends sdprb1
* SPICE INPUT		Tue Jul 31 20:30:20 2018	sdprb2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprb2
.subckt sdprb2 GND Q QN SN VDD CK SI D SE
M1 N_25 D GND GND mn15  l=0.13u w=0.33u m=1
M2 N_25 N_3 N_5 GND mn15  l=0.13u w=0.33u m=1
M3 N_26 SE N_5 GND mn15  l=0.13u w=0.24u m=1
M4 GND SE N_3 GND mn15  l=0.13u w=0.24u m=1
M5 N_26 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.23u m=1
M7 N_27 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M8 N_10 N_2 N_5 GND mn15  l=0.13u w=0.28u m=1
M9 GND N_2 N_7 GND mn15  l=0.13u w=0.17u m=1
M10 N_27 N_7 N_10 GND mn15  l=0.13u w=0.17u m=1
M11 N_12 N_10 N_11 GND mn15  l=0.13u w=0.24u m=1
M12 N_11 N_10 N_12 GND mn15  l=0.13u w=0.22u m=1
M13 N_15 N_2 N_28 GND mn15  l=0.13u w=0.17u m=1
M14 N_15 N_7 N_12 GND mn15  l=0.13u w=0.36u m=1
M15 N_28 N_23 N_11 GND mn15  l=0.13u w=0.17u m=1
M16 N_11 SN GND GND mn15  l=0.13u w=0.47u m=1
M17 N_11 SN GND GND mn15  l=0.13u w=0.47u m=1
M18 GND N_23 Q GND mn15  l=0.13u w=0.46u m=1
M19 GND N_23 Q GND mn15  l=0.13u w=0.46u m=1
M20 GND N_15 QN GND mn15  l=0.13u w=0.46u m=1
M21 GND N_15 QN GND mn15  l=0.13u w=0.46u m=1
M22 GND N_15 N_23 GND mn15  l=0.13u w=0.37u m=1
M23 N_45 D VDD VDD mp15  l=0.13u w=0.5u m=1
M24 N_5 SE N_45 VDD mp15  l=0.13u w=0.5u m=1
M25 N_3 SE VDD VDD mp15  l=0.13u w=0.37u m=1
M26 N_46 N_3 N_5 VDD mp15  l=0.13u w=0.37u m=1
M27 N_46 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M28 N_2 CK VDD VDD mp15  l=0.13u w=0.57u m=1
M29 N_47 N_12 VDD VDD mp15  l=0.13u w=0.17u m=1
M30 VDD N_2 N_7 VDD mp15  l=0.13u w=0.42u m=1
M31 N_47 N_2 N_10 VDD mp15  l=0.13u w=0.17u m=1
M32 N_5 N_7 N_10 VDD mp15  l=0.13u w=0.42u m=1
M33 N_12 N_10 VDD VDD mp15  l=0.13u w=0.32u m=1
M34 N_12 N_10 VDD VDD mp15  l=0.13u w=0.31u m=1
M35 N_48 N_23 VDD VDD mp15  l=0.13u w=0.17u m=1
M36 N_15 N_2 N_12 VDD mp15  l=0.13u w=0.56u m=1
M37 N_15 N_7 N_48 VDD mp15  l=0.13u w=0.17u m=1
M38 N_15 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M39 N_15 SN VDD VDD mp15  l=0.13u w=0.28u m=1
M40 Q N_23 VDD VDD mp15  l=0.13u w=0.69u m=1
M41 VDD N_23 Q VDD mp15  l=0.13u w=0.69u m=1
M42 VDD N_15 QN VDD mp15  l=0.13u w=0.69u m=1
M43 VDD N_15 QN VDD mp15  l=0.13u w=0.69u m=1
M44 N_23 N_15 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends sdprb2
* SPICE INPUT		Tue Jul 31 20:30:32 2018	sdprq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq0
.subckt sdprq0 GND Q VDD SN CK SI D SE
M1 N_20 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_20 N_4 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M4 N_21 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M5 N_21 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.18u m=1
M7 Q N_10 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_9 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_22 N_6 GND GND mn15  l=0.13u w=0.17u m=1
M10 N_23 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_24 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M12 GND N_18 N_10 GND mn15  l=0.13u w=0.18u m=1
M13 N_15 N_13 GND GND mn15  l=0.13u w=0.22u m=1
M14 N_10 N_11 N_15 GND mn15  l=0.13u w=0.22u m=1
M15 N_23 N_11 N_13 GND mn15  l=0.13u w=0.17u m=1
M16 GND N_2 N_11 GND mn15  l=0.13u w=0.17u m=1
M17 N_24 N_2 N_10 GND mn15  l=0.13u w=0.17u m=1
M18 N_22 N_2 N_13 GND mn15  l=0.13u w=0.17u m=1
M19 GND SN N_18 GND mn15  l=0.13u w=0.18u m=1
M20 Q N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_9 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_95 D VDD VDD mp15  l=0.13u w=0.28u m=1
M23 N_96 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M24 N_95 SE N_6 VDD mp15  l=0.13u w=0.28u m=1
M25 N_4 SE VDD VDD mp15  l=0.13u w=0.26u m=1
M26 N_96 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M27 N_2 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M28 N_98 N_6 VDD VDD mp15  l=0.13u w=0.36u m=1
M29 N_98 N_11 N_13 VDD mp15  l=0.13u w=0.36u m=1
M30 N_97 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M31 N_13 N_2 N_97 VDD mp15  l=0.13u w=0.17u m=1
M32 N_11 N_2 VDD VDD mp15  l=0.13u w=0.42u m=1
M33 N_99 N_9 N_32 VDD mp15  l=0.13u w=0.17u m=1
M34 N_32 N_18 VDD VDD mp15  l=0.13u w=0.57u m=1
M35 N_15 N_13 N_32 VDD mp15  l=0.13u w=0.2u m=1
M36 N_32 N_13 N_15 VDD mp15  l=0.13u w=0.2u m=1
M37 N_10 N_2 N_15 VDD mp15  l=0.13u w=0.42u m=1
M38 N_99 N_11 N_10 VDD mp15  l=0.13u w=0.17u m=1
M39 VDD SN N_18 VDD mp15  l=0.13u w=0.26u m=1
.ends sdprq0
* SPICE INPUT		Tue Jul 31 20:30:45 2018	sdprq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq1
.subckt sdprq1 GND Q VDD SN CK SI D SE
M1 N_20 D GND GND mn15  l=0.13u w=0.28u m=1
M2 N_20 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M3 GND SE N_4 GND mn15  l=0.13u w=0.18u m=1
M4 N_21 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M5 N_21 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 N_22 N_6 GND GND mn15  l=0.13u w=0.35u m=1
M8 N_23 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_12 N_10 GND GND mn15  l=0.13u w=0.27u m=1
M10 N_7 N_8 N_12 GND mn15  l=0.13u w=0.35u m=1
M11 N_23 N_8 N_10 GND mn15  l=0.13u w=0.17u m=1
M12 N_22 N_2 N_10 GND mn15  l=0.13u w=0.35u m=1
M13 N_24 N_2 N_7 GND mn15  l=0.13u w=0.17u m=1
M14 GND N_2 N_8 GND mn15  l=0.13u w=0.2u m=1
M15 N_24 N_19 GND GND mn15  l=0.13u w=0.17u m=1
M16 GND N_15 N_7 GND mn15  l=0.13u w=0.28u m=1
M17 GND SN N_15 GND mn15  l=0.13u w=0.18u m=1
M18 Q N_7 GND GND mn15  l=0.13u w=0.46u m=1
M19 N_19 N_7 GND GND mn15  l=0.13u w=0.17u m=1
M20 N_100 D VDD VDD mp15  l=0.13u w=0.42u m=1
M21 N_101 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M22 N_100 SE N_6 VDD mp15  l=0.13u w=0.42u m=1
M23 N_4 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M24 N_101 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M25 N_2 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M26 N_103 N_6 VDD VDD mp15  l=0.13u w=0.53u m=1
M27 N_103 N_8 N_10 VDD mp15  l=0.13u w=0.53u m=1
M28 N_102 N_12 VDD VDD mp15  l=0.13u w=0.17u m=1
M29 N_10 N_2 N_102 VDD mp15  l=0.13u w=0.17u m=1
M30 N_8 N_2 VDD VDD mp15  l=0.13u w=0.51u m=1
M31 N_12 N_10 N_32 VDD mp15  l=0.13u w=0.32u m=1
M32 N_12 N_10 N_32 VDD mp15  l=0.13u w=0.32u m=1
M33 N_7 N_2 N_12 VDD mp15  l=0.13u w=0.54u m=1
M34 N_104 N_8 N_7 VDD mp15  l=0.13u w=0.17u m=1
M35 N_32 N_19 N_104 VDD mp15  l=0.13u w=0.17u m=1
M36 N_32 N_15 VDD VDD mp15  l=0.13u w=0.69u m=1
M37 VDD SN N_15 VDD mp15  l=0.13u w=0.28u m=1
M38 Q N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M39 N_19 N_7 VDD VDD mp15  l=0.13u w=0.17u m=1
.ends sdprq1
* SPICE INPUT		Tue Jul 31 20:30:58 2018	sdprq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprq2
.subckt sdprq2 GND Q VDD SN CK SI D SE
M1 Q N_7 GND GND mn15  l=0.13u w=0.46u m=1
M2 Q N_7 GND GND mn15  l=0.13u w=0.46u m=1
M3 GND N_7 N_4 GND mn15  l=0.13u w=0.17u m=1
M4 GND SN N_2 GND mn15  l=0.13u w=0.24u m=1
M5 GND N_2 N_7 GND mn15  l=0.13u w=0.36u m=1
M6 N_12 N_10 N_22 GND mn15  l=0.13u w=0.17u m=1
M7 N_23 N_18 N_12 GND mn15  l=0.13u w=0.37u m=1
M8 GND N_18 N_10 GND mn15  l=0.13u w=0.2u m=1
M9 N_23 N_21 GND GND mn15  l=0.13u w=0.37u m=1
M10 N_22 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_7 N_10 N_15 GND mn15  l=0.13u w=0.37u m=1
M12 N_7 N_18 N_24 GND mn15  l=0.13u w=0.17u m=1
M13 N_24 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M14 N_15 N_12 GND GND mn15  l=0.13u w=0.27u m=1
M15 N_18 CK GND GND mn15  l=0.13u w=0.28u m=1
M16 N_26 SI GND GND mn15  l=0.13u w=0.24u m=1
M17 N_26 SE N_21 GND mn15  l=0.13u w=0.24u m=1
M18 GND SE N_19 GND mn15  l=0.13u w=0.18u m=1
M19 N_25 N_19 N_21 GND mn15  l=0.13u w=0.24u m=1
M20 N_25 D GND GND mn15  l=0.13u w=0.24u m=1
M21 N_18 CK VDD VDD mp15  l=0.13u w=0.7u m=1
M22 N_46 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M23 N_46 N_19 N_21 VDD mp15  l=0.13u w=0.37u m=1
M24 N_21 SE N_45 VDD mp15  l=0.13u w=0.37u m=1
M25 N_19 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M26 N_45 D VDD VDD mp15  l=0.13u w=0.37u m=1
M27 Q N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M28 Q N_7 VDD VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_7 N_4 VDD mp15  l=0.13u w=0.17u m=1
M30 N_2 SN VDD VDD mp15  l=0.13u w=0.34u m=1
M31 N_10 N_18 VDD VDD mp15  l=0.13u w=0.51u m=1
M32 N_12 N_18 N_47 VDD mp15  l=0.13u w=0.17u m=1
M33 N_48 N_21 VDD VDD mp15  l=0.13u w=0.53u m=1
M34 N_48 N_10 N_12 VDD mp15  l=0.13u w=0.53u m=1
M35 N_47 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M36 N_7 N_18 N_15 VDD mp15  l=0.13u w=0.57u m=1
M37 N_34 N_2 VDD VDD mp15  l=0.13u w=0.68u m=1
M38 VDD N_2 N_34 VDD mp15  l=0.13u w=0.39u m=1
M39 N_34 N_4 N_49 VDD mp15  l=0.13u w=0.17u m=1
M40 N_15 N_12 N_34 VDD mp15  l=0.13u w=0.32u m=1
M41 N_15 N_12 N_34 VDD mp15  l=0.13u w=0.32u m=1
M42 N_15 N_12 N_34 VDD mp15  l=0.13u w=0.32u m=1
M43 N_49 N_10 N_7 VDD mp15  l=0.13u w=0.17u m=1
.ends sdprq2
* SPICE INPUT		Tue Jul 31 20:31:11 2018	sdprqm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdprqm
.subckt sdprqm GND Q VDD SN CK SI D SE
M1 N_20 D GND GND mn15  l=0.13u w=0.18u m=1
M2 N_20 N_4 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 N_21 SE N_6 GND mn15  l=0.13u w=0.18u m=1
M4 GND SE N_4 GND mn15  l=0.13u w=0.17u m=1
M5 N_21 SI GND GND mn15  l=0.13u w=0.18u m=1
M6 GND CK N_2 GND mn15  l=0.13u w=0.2u m=1
M7 Q N_10 GND GND mn15  l=0.13u w=0.36u m=1
M8 N_9 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M9 N_22 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M10 N_23 N_15 GND GND mn15  l=0.13u w=0.17u m=1
M11 N_24 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M12 GND N_18 N_10 GND mn15  l=0.13u w=0.24u m=1
M13 N_15 N_13 GND GND mn15  l=0.13u w=0.27u m=1
M14 N_10 N_11 N_15 GND mn15  l=0.13u w=0.28u m=1
M15 N_23 N_11 N_13 GND mn15  l=0.13u w=0.17u m=1
M16 N_22 N_2 N_13 GND mn15  l=0.13u w=0.28u m=1
M17 N_24 N_2 N_10 GND mn15  l=0.13u w=0.17u m=1
M18 GND N_2 N_11 GND mn15  l=0.13u w=0.17u m=1
M19 GND SN N_18 GND mn15  l=0.13u w=0.17u m=1
M20 Q N_10 VDD VDD mp15  l=0.13u w=0.55u m=1
M21 N_9 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M22 N_100 D VDD VDD mp15  l=0.13u w=0.28u m=1
M23 N_101 N_4 N_6 VDD mp15  l=0.13u w=0.28u m=1
M24 N_100 SE N_6 VDD mp15  l=0.13u w=0.28u m=1
M25 VDD SE N_4 VDD mp15  l=0.13u w=0.24u m=1
M26 N_101 SI VDD VDD mp15  l=0.13u w=0.28u m=1
M27 N_2 CK VDD VDD mp15  l=0.13u w=0.46u m=1
M28 N_103 N_6 VDD VDD mp15  l=0.13u w=0.42u m=1
M29 N_103 N_11 N_13 VDD mp15  l=0.13u w=0.42u m=1
M30 N_102 N_15 VDD VDD mp15  l=0.13u w=0.17u m=1
M31 N_11 N_2 VDD VDD mp15  l=0.13u w=0.42u m=1
M32 N_13 N_2 N_102 VDD mp15  l=0.13u w=0.17u m=1
M33 N_104 N_9 N_32 VDD mp15  l=0.13u w=0.17u m=1
M34 N_32 N_18 VDD VDD mp15  l=0.13u w=0.61u m=1
M35 N_15 N_13 N_32 VDD mp15  l=0.13u w=0.305u m=1
M36 N_32 N_13 N_15 VDD mp15  l=0.13u w=0.305u m=1
M37 N_10 N_2 N_15 VDD mp15  l=0.13u w=0.42u m=1
M38 N_104 N_11 N_10 VDD mp15  l=0.13u w=0.17u m=1
M39 VDD SN N_18 VDD mp15  l=0.13u w=0.24u m=1
.ends sdprqm
* SPICE INPUT		Tue Jul 31 20:31:24 2018	sdscrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdscrq0
.subckt sdscrq0 GND Q VDD CK SE SI RN D
M1 Q N_15 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_4 N_15 GND GND mn15  l=0.13u w=0.18u m=1
M3 N_18 D GND GND mn15  l=0.13u w=0.26u m=1
M4 N_8 RN N_18 GND mn15  l=0.13u w=0.26u m=1
M5 N_19 SE N_9 GND mn15  l=0.13u w=0.24u m=1
M6 N_9 N_5 N_8 GND mn15  l=0.13u w=0.28u m=1
M7 N_19 SI GND GND mn15  l=0.13u w=0.24u m=1
M8 GND SE N_5 GND mn15  l=0.13u w=0.18u m=1
M9 N_22 N_4 GND GND mn15  l=0.13u w=0.17u m=1
M10 N_16 N_10 N_15 GND mn15  l=0.13u w=0.28u m=1
M11 N_22 N_11 N_15 GND mn15  l=0.13u w=0.17u m=1
M12 GND N_11 N_10 GND mn15  l=0.13u w=0.17u m=1
M13 GND CK N_11 GND mn15  l=0.13u w=0.17u m=1
M14 N_20 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M15 N_13 N_11 N_20 GND mn15  l=0.13u w=0.28u m=1
M16 N_21 N_10 N_13 GND mn15  l=0.13u w=0.17u m=1
M17 N_21 N_16 GND GND mn15  l=0.13u w=0.17u m=1
M18 N_16 N_13 GND GND mn15  l=0.13u w=0.28u m=1
M19 VDD D N_8 VDD mp15  l=0.13u w=0.35u m=1
M20 N_8 RN VDD VDD mp15  l=0.13u w=0.35u m=1
M21 N_38 N_5 N_9 VDD mp15  l=0.13u w=0.37u m=1
M22 N_38 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M23 N_9 SE N_8 VDD mp15  l=0.13u w=0.42u m=1
M24 N_5 SE VDD VDD mp15  l=0.13u w=0.28u m=1
M25 N_41 N_4 VDD VDD mp15  l=0.13u w=0.17u m=1
M26 N_10 N_11 VDD VDD mp15  l=0.13u w=0.42u m=1
M27 N_15 N_11 N_16 VDD mp15  l=0.13u w=0.42u m=1
M28 N_41 N_10 N_15 VDD mp15  l=0.13u w=0.17u m=1
M29 VDD CK N_11 VDD mp15  l=0.13u w=0.42u m=1
M30 N_39 N_9 VDD VDD mp15  l=0.13u w=0.42u m=1
M31 N_13 N_10 N_39 VDD mp15  l=0.13u w=0.42u m=1
M32 N_40 N_11 N_13 VDD mp15  l=0.13u w=0.17u m=1
M33 VDD N_16 N_40 VDD mp15  l=0.13u w=0.17u m=1
M34 N_16 N_13 VDD VDD mp15  l=0.13u w=0.42u m=1
M35 Q N_15 VDD VDD mp15  l=0.13u w=0.4u m=1
M36 N_4 N_15 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends sdscrq0
* SPICE INPUT		Tue Jul 31 20:31:38 2018	sdscrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdscrq1
.subckt sdscrq1 GND Q VDD CK SE SI RN D
M1 N_18 D GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 RN N_18 GND mn15  l=0.13u w=0.26u m=1
M3 N_19 SE N_6 GND mn15  l=0.13u w=0.24u m=1
M4 N_6 N_2 N_5 GND mn15  l=0.13u w=0.28u m=1
M5 N_19 SI GND GND mn15  l=0.13u w=0.24u m=1
M6 GND SE N_2 GND mn15  l=0.13u w=0.18u m=1
M7 Q N_17 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_9 N_17 GND GND mn15  l=0.13u w=0.28u m=1
M9 N_22 N_12 N_17 GND mn15  l=0.13u w=0.17u m=1
M10 GND N_12 N_10 GND mn15  l=0.13u w=0.2u m=1
M11 GND CK N_12 GND mn15  l=0.13u w=0.2u m=1
M12 N_20 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M13 N_20 N_12 N_14 GND mn15  l=0.13u w=0.28u m=1
M14 N_21 N_10 N_14 GND mn15  l=0.13u w=0.17u m=1
M15 GND N_16 N_21 GND mn15  l=0.13u w=0.17u m=1
M16 N_16 N_14 GND GND mn15  l=0.13u w=0.36u m=1
M17 N_22 N_9 GND GND mn15  l=0.13u w=0.17u m=1
M18 N_17 N_10 N_16 GND mn15  l=0.13u w=0.36u m=1
M19 N_5 D VDD VDD mp15  l=0.13u w=0.35u m=1
M20 N_5 RN VDD VDD mp15  l=0.13u w=0.35u m=1
M21 N_91 N_2 N_6 VDD mp15  l=0.13u w=0.37u m=1
M22 N_91 SI VDD VDD mp15  l=0.13u w=0.37u m=1
M23 N_6 SE N_5 VDD mp15  l=0.13u w=0.42u m=1
M24 VDD SE N_2 VDD mp15  l=0.13u w=0.28u m=1
M25 N_17 N_12 N_16 VDD mp15  l=0.13u w=0.52u m=1
M26 N_10 N_12 VDD VDD mp15  l=0.13u w=0.51u m=1
M27 N_94 N_10 N_17 VDD mp15  l=0.13u w=0.17u m=1
M28 N_12 CK VDD VDD mp15  l=0.13u w=0.51u m=1
M29 N_92 N_6 VDD VDD mp15  l=0.13u w=0.42u m=1
M30 N_92 N_10 N_14 VDD mp15  l=0.13u w=0.42u m=1
M31 N_93 N_12 N_14 VDD mp15  l=0.13u w=0.17u m=1
M32 VDD N_16 N_93 VDD mp15  l=0.13u w=0.17u m=1
M33 N_16 N_14 VDD VDD mp15  l=0.13u w=0.52u m=1
M34 N_94 N_9 VDD VDD mp15  l=0.13u w=0.17u m=1
M35 Q N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M36 N_9 N_17 VDD VDD mp15  l=0.13u w=0.35u m=1
.ends sdscrq1
* SPICE INPUT		Tue Jul 31 20:31:51 2018	sdscrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=sdscrq2
.subckt sdscrq2 GND Q VDD CK SI SE RN D
M1 GND D N_20 GND mn15  l=0.13u w=0.46u m=1
M2 N_2 RN N_20 GND mn15  l=0.13u w=0.46u m=1
M3 N_2 N_4 N_6 GND mn15  l=0.13u w=0.41u m=1
M4 N_21 SI GND GND mn15  l=0.13u w=0.28u m=1
M5 N_21 SE N_6 GND mn15  l=0.13u w=0.28u m=1
M6 GND SE N_4 GND mn15  l=0.13u w=0.24u m=1
M7 GND N_18 Q GND mn15  l=0.13u w=0.46u m=1
M8 GND N_18 Q GND mn15  l=0.13u w=0.46u m=1
M9 GND N_18 N_10 GND mn15  l=0.13u w=0.37u m=1
M10 GND CK N_13 GND mn15  l=0.13u w=0.28u m=1
M11 N_22 N_6 GND GND mn15  l=0.13u w=0.41u m=1
M12 N_22 N_13 N_15 GND mn15  l=0.13u w=0.41u m=1
M13 N_23 N_12 N_15 GND mn15  l=0.13u w=0.17u m=1
M14 GND N_17 N_23 GND mn15  l=0.13u w=0.17u m=1
M15 N_17 N_15 GND GND mn15  l=0.13u w=0.41u m=1
M16 N_18 N_12 N_17 GND mn15  l=0.13u w=0.41u m=1
M17 N_24 N_10 GND GND mn15  l=0.13u w=0.17u m=1
M18 N_24 N_13 N_18 GND mn15  l=0.13u w=0.17u m=1
M19 GND N_13 N_12 GND mn15  l=0.13u w=0.22u m=1
M20 VDD D N_2 VDD mp15  l=0.13u w=0.61u m=1
M21 N_2 RN VDD VDD mp15  l=0.13u w=0.61u m=1
M22 N_6 SE N_2 VDD mp15  l=0.13u w=0.63u m=1
M23 N_98 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M24 N_98 SI VDD VDD mp15  l=0.13u w=0.4u m=1
M25 VDD SE N_4 VDD mp15  l=0.13u w=0.37u m=1
M26 N_13 CK VDD VDD mp15  l=0.13u w=0.67u m=1
M27 N_99 N_6 VDD VDD mp15  l=0.13u w=0.62u m=1
M28 N_100 N_13 N_15 VDD mp15  l=0.13u w=0.17u m=1
M29 N_99 N_12 N_15 VDD mp15  l=0.13u w=0.62u m=1
M30 N_100 N_17 VDD VDD mp15  l=0.13u w=0.17u m=1
M31 N_17 N_15 VDD VDD mp15  l=0.13u w=0.32u m=1
M32 N_17 N_15 VDD VDD mp15  l=0.13u w=0.31u m=1
M33 N_101 N_12 N_18 VDD mp15  l=0.13u w=0.17u m=1
M34 N_101 N_10 VDD VDD mp15  l=0.13u w=0.17u m=1
M35 N_18 N_13 N_17 VDD mp15  l=0.13u w=0.63u m=1
M36 VDD N_13 N_12 VDD mp15  l=0.13u w=0.55u m=1
M37 VDD N_18 Q VDD mp15  l=0.13u w=0.69u m=1
M38 VDD N_18 Q VDD mp15  l=0.13u w=0.69u m=1
M39 N_10 N_18 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends sdscrq2
* SPICE INPUT		Tue Jul 31 20:32:05 2018	senrq0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=senrq0
.subckt senrq0 GND Q D E SE VDD CK SI
M1 N_5 N_14 N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_22 N_6 N_4 GND mn15  l=0.13u w=0.17u m=1
M3 N_22 N_2 GND GND mn15  l=0.13u w=0.17u m=1
M4 GND N_4 N_2 GND mn15  l=0.13u w=0.18u m=1
M5 Q N_4 GND GND mn15  l=0.13u w=0.26u m=1
M6 GND CK N_6 GND mn15  l=0.13u w=0.17u m=1
M7 GND E N_11 GND mn15  l=0.13u w=0.18u m=1
M8 N_23 D GND GND mn15  l=0.13u w=0.18u m=1
M9 N_23 E N_13 GND mn15  l=0.13u w=0.18u m=1
M10 N_24 N_11 N_13 GND mn15  l=0.13u w=0.18u m=1
M11 N_24 N_2 GND GND mn15  l=0.13u w=0.18u m=1
M12 GND SE N_9 GND mn15  l=0.13u w=0.18u m=1
M13 N_25 SE N_17 GND mn15  l=0.13u w=0.24u m=1
M14 N_17 N_9 N_13 GND mn15  l=0.13u w=0.28u m=1
M15 N_25 SI GND GND mn15  l=0.13u w=0.24u m=1
M16 N_26 N_17 GND GND mn15  l=0.13u w=0.28u m=1
M17 N_19 N_6 N_26 GND mn15  l=0.13u w=0.28u m=1
M18 GND N_5 N_27 GND mn15  l=0.13u w=0.17u m=1
M19 N_5 N_19 GND GND mn15  l=0.13u w=0.14u m=1
M20 N_5 N_19 GND GND mn15  l=0.13u w=0.14u m=1
M21 N_27 N_14 N_19 GND mn15  l=0.13u w=0.17u m=1
M22 GND N_6 N_14 GND mn15  l=0.13u w=0.17u m=1
M23 N_42 N_14 N_4 VDD mp15  l=0.13u w=0.17u m=1
M24 N_42 N_2 VDD VDD mp15  l=0.13u w=0.17u m=1
M25 N_4 N_6 N_5 VDD mp15  l=0.13u w=0.42u m=1
M26 VDD N_4 N_2 VDD mp15  l=0.13u w=0.26u m=1
M27 Q N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M28 N_6 CK VDD VDD mp15  l=0.13u w=0.42u m=1
M29 N_13 SE N_17 VDD mp15  l=0.13u w=0.42u m=1
M30 N_43 N_9 N_17 VDD mp15  l=0.13u w=0.37u m=1
M31 VDD SI N_43 VDD mp15  l=0.13u w=0.37u m=1
M32 N_44 N_17 VDD VDD mp15  l=0.13u w=0.42u m=1
M33 N_45 N_6 N_19 VDD mp15  l=0.13u w=0.17u m=1
M34 VDD N_5 N_45 VDD mp15  l=0.13u w=0.17u m=1
M35 N_5 N_19 VDD VDD mp15  l=0.13u w=0.21u m=1
M36 N_5 N_19 VDD VDD mp15  l=0.13u w=0.21u m=1
M37 N_44 N_14 N_19 VDD mp15  l=0.13u w=0.42u m=1
M38 N_14 N_6 VDD VDD mp15  l=0.13u w=0.42u m=1
M39 VDD E N_11 VDD mp15  l=0.13u w=0.26u m=1
M40 N_46 D VDD VDD mp15  l=0.13u w=0.28u m=1
M41 N_13 N_11 N_46 VDD mp15  l=0.13u w=0.28u m=1
M42 N_47 E N_13 VDD mp15  l=0.13u w=0.28u m=1
M43 N_47 N_2 VDD VDD mp15  l=0.13u w=0.28u m=1
M44 VDD SE N_9 VDD mp15  l=0.13u w=0.28u m=1
.ends senrq0
* SPICE INPUT		Tue Jul 31 20:32:20 2018	senrq1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=senrq1
.subckt senrq1 GND Q SE VDD CK SI E D
M1 GND E N_4 GND mn15  l=0.13u w=0.17u m=1
M2 N_22 D GND GND mn15  l=0.13u w=0.28u m=1
M3 N_6 E N_22 GND mn15  l=0.13u w=0.28u m=1
M4 N_23 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_23 N_16 GND GND mn15  l=0.13u w=0.28u m=1
M6 GND SE N_2 GND mn15  l=0.13u w=0.18u m=1
M7 N_24 SE N_10 GND mn15  l=0.13u w=0.24u m=1
M8 N_10 N_2 N_6 GND mn15  l=0.13u w=0.28u m=1
M9 N_24 SI GND GND mn15  l=0.13u w=0.24u m=1
M10 N_25 N_10 GND GND mn15  l=0.13u w=0.28u m=1
M11 N_12 N_19 N_25 GND mn15  l=0.13u w=0.28u m=1
M12 GND N_14 N_26 GND mn15  l=0.13u w=0.17u m=1
M13 N_14 N_12 GND GND mn15  l=0.13u w=0.19u m=1
M14 N_14 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M15 N_26 N_7 N_12 GND mn15  l=0.13u w=0.17u m=1
M16 GND N_19 N_7 GND mn15  l=0.13u w=0.2u m=1
M17 N_14 N_7 N_17 GND mn15  l=0.13u w=0.36u m=1
M18 N_27 N_19 N_17 GND mn15  l=0.13u w=0.17u m=1
M19 N_27 N_16 GND GND mn15  l=0.13u w=0.17u m=1
M20 N_16 N_17 GND GND mn15  l=0.13u w=0.28u m=1
M21 Q N_17 GND GND mn15  l=0.13u w=0.46u m=1
M22 GND CK N_19 GND mn15  l=0.13u w=0.2u m=1
M23 VDD E N_4 VDD mp15  l=0.13u w=0.24u m=1
M24 N_48 D VDD VDD mp15  l=0.13u w=0.42u m=1
M25 N_6 N_4 N_48 VDD mp15  l=0.13u w=0.42u m=1
M26 N_49 E N_6 VDD mp15  l=0.13u w=0.42u m=1
M27 N_49 N_16 VDD VDD mp15  l=0.13u w=0.42u m=1
M28 VDD SE N_2 VDD mp15  l=0.13u w=0.28u m=1
M29 N_6 SE N_10 VDD mp15  l=0.13u w=0.42u m=1
M30 N_50 N_2 N_10 VDD mp15  l=0.13u w=0.37u m=1
M31 VDD SI N_50 VDD mp15  l=0.13u w=0.37u m=1
M32 N_51 N_10 VDD VDD mp15  l=0.13u w=0.42u m=1
M33 N_52 N_19 N_12 VDD mp15  l=0.13u w=0.17u m=1
M34 VDD N_14 N_52 VDD mp15  l=0.13u w=0.17u m=1
M35 N_14 N_12 VDD VDD mp15  l=0.13u w=0.26u m=1
M36 N_14 N_12 VDD VDD mp15  l=0.13u w=0.26u m=1
M37 N_51 N_7 N_12 VDD mp15  l=0.13u w=0.42u m=1
M38 N_7 N_19 VDD VDD mp15  l=0.13u w=0.51u m=1
M39 N_53 N_7 N_17 VDD mp15  l=0.13u w=0.17u m=1
M40 N_53 N_16 VDD VDD mp15  l=0.13u w=0.17u m=1
M41 N_17 N_19 N_14 VDD mp15  l=0.13u w=0.52u m=1
M42 VDD N_17 N_16 VDD mp15  l=0.13u w=0.35u m=1
M43 Q N_17 VDD VDD mp15  l=0.13u w=0.69u m=1
M44 N_19 CK VDD VDD mp15  l=0.13u w=0.51u m=1
.ends senrq1
* SPICE INPUT		Tue Jul 31 20:32:33 2018	senrq2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=senrq2
.subckt senrq2 VDD Q GND CK SI SE E D
M1 GND E N_4 GND mn15  l=0.13u w=0.24u m=1
M2 N_44 D GND GND mn15  l=0.13u w=0.28u m=1
M3 N_6 E N_44 GND mn15  l=0.13u w=0.28u m=1
M4 N_45 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_45 N_21 GND GND mn15  l=0.13u w=0.28u m=1
M6 GND SE N_2 GND mn15  l=0.13u w=0.24u m=1
M7 N_9 N_2 N_6 GND mn15  l=0.13u w=0.41u m=1
M8 N_46 SE N_9 GND mn15  l=0.13u w=0.28u m=1
M9 N_46 SI GND GND mn15  l=0.13u w=0.28u m=1
M10 N_47 N_9 GND GND mn15  l=0.13u w=0.41u m=1
M11 N_12 N_19 N_47 GND mn15  l=0.13u w=0.41u m=1
M12 GND N_14 N_48 GND mn15  l=0.13u w=0.17u m=1
M13 N_14 N_12 GND GND mn15  l=0.13u w=0.25u m=1
M14 N_14 N_12 GND GND mn15  l=0.13u w=0.17u m=1
M15 N_48 N_8 N_12 GND mn15  l=0.13u w=0.17u m=1
M16 GND N_19 N_8 GND mn15  l=0.13u w=0.23u m=1
M17 Q N_16 GND GND mn15  l=0.13u w=0.46u m=1
M18 Q N_16 GND GND mn15  l=0.13u w=0.46u m=1
M19 GND N_16 N_21 GND mn15  l=0.13u w=0.37u m=1
M20 N_19 CK GND GND mn15  l=0.13u w=0.28u m=1
M21 N_14 N_8 N_16 GND mn15  l=0.13u w=0.41u m=1
M22 N_16 N_19 N_49 GND mn15  l=0.13u w=0.17u m=1
M23 N_49 N_21 GND GND mn15  l=0.13u w=0.17u m=1
M24 VDD E N_4 VDD mp15  l=0.13u w=0.37u m=1
M25 N_23 D VDD VDD mp15  l=0.13u w=0.42u m=1
M26 N_6 N_4 N_23 VDD mp15  l=0.13u w=0.42u m=1
M27 N_24 E N_6 VDD mp15  l=0.13u w=0.42u m=1
M28 N_24 N_21 VDD VDD mp15  l=0.13u w=0.42u m=1
M29 VDD SE N_2 VDD mp15  l=0.13u w=0.37u m=1
M30 N_6 SE N_9 VDD mp15  l=0.13u w=0.63u m=1
M31 N_25 N_2 N_9 VDD mp15  l=0.13u w=0.42u m=1
M32 VDD SI N_25 VDD mp15  l=0.13u w=0.42u m=1
M33 N_26 N_9 VDD VDD mp15  l=0.13u w=0.62u m=1
M34 N_27 N_19 N_12 VDD mp15  l=0.13u w=0.17u m=1
M35 VDD N_14 N_27 VDD mp15  l=0.13u w=0.17u m=1
M36 N_14 N_12 VDD VDD mp15  l=0.13u w=0.305u m=1
M37 N_14 N_12 VDD VDD mp15  l=0.13u w=0.325u m=1
M38 N_26 N_8 N_12 VDD mp15  l=0.13u w=0.62u m=1
M39 N_8 N_19 VDD VDD mp15  l=0.13u w=0.55u m=1
M40 N_14 N_19 N_16 VDD mp15  l=0.13u w=0.62u m=1
M41 N_28 N_8 N_16 VDD mp15  l=0.13u w=0.17u m=1
M42 N_28 N_21 VDD VDD mp15  l=0.13u w=0.17u m=1
M43 Q N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M44 Q N_16 VDD VDD mp15  l=0.13u w=0.69u m=1
M45 N_21 N_16 VDD VDD mp15  l=0.13u w=0.55u m=1
M46 N_19 CK VDD VDD mp15  l=0.13u w=0.69u m=1
.ends senrq2
* SPICE INPUT		Tue Jul 31 20:32:47 2018	tiehi
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tiehi
.subckt tiehi VDD GND Y
M1 N_5 N_5 GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends tiehi
* SPICE INPUT		Tue Jul 31 20:33:00 2018	tielo
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tielo
.subckt tielo Y VDD GND
M1 Y N_5 GND GND mn15  l=0.13u w=0.26u m=1
M2 N_5 N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
.ends tielo
* SPICE INPUT		Tue Jul 31 20:33:14 2018	tlatncad0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad0
.subckt tlatncad0 VDD ECK GND CK E
M1 GND N_6 N_3 GND mn15  l=0.13u w=0.26u m=1
M2 N_50 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_50 N_5 N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_49 N_10 N_6 GND mn15  l=0.13u w=0.18u m=1
M5 GND N_10 N_5 GND mn15  l=0.13u w=0.18u m=1
M6 N_49 E GND GND mn15  l=0.13u w=0.18u m=1
M7 N_10 CK GND GND mn15  l=0.13u w=0.23u m=1
M8 N_51 CK N_11 GND mn15  l=0.13u w=0.26u m=1
M9 N_51 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M10 ECK N_11 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_3 N_6 VDD VDD mp15  l=0.13u w=0.38u m=1
M12 N_13 N_3 VDD VDD mp15  l=0.13u w=0.26u m=1
M13 N_12 N_5 N_6 VDD mp15  l=0.13u w=0.27u m=1
M14 N_5 N_10 VDD VDD mp15  l=0.13u w=0.46u m=1
M15 N_13 N_10 N_6 VDD mp15  l=0.13u w=0.26u m=1
M16 N_12 E VDD VDD mp15  l=0.13u w=0.27u m=1
M17 N_10 CK VDD VDD mp15  l=0.13u w=0.58u m=1
M18 N_11 CK VDD VDD mp15  l=0.13u w=0.31u m=1
M19 N_11 N_3 VDD VDD mp15  l=0.13u w=0.31u m=1
M20 ECK N_11 VDD VDD mp15  l=0.13u w=0.65u m=1
.ends tlatncad0
* SPICE INPUT		Tue Jul 31 20:33:27 2018	tlatncad1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad1
.subckt tlatncad1 VDD ECK GND CK E
M1 N_49 E GND GND mn15  l=0.13u w=0.18u m=1
M2 N_49 N_10 N_6 GND mn15  l=0.13u w=0.18u m=1
M3 GND N_10 N_5 GND mn15  l=0.13u w=0.18u m=1
M4 N_50 N_5 N_6 GND mn15  l=0.13u w=0.26u m=1
M5 N_50 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M6 GND N_6 N_3 GND mn15  l=0.13u w=0.26u m=1
M7 N_10 CK GND GND mn15  l=0.13u w=0.23u m=1
M8 N_51 CK N_11 GND mn15  l=0.13u w=0.26u m=1
M9 N_51 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M10 ECK N_11 GND GND mn15  l=0.13u w=0.27u m=1
M11 N_12 E VDD VDD mp15  l=0.13u w=0.27u m=1
M12 N_5 N_10 VDD VDD mp15  l=0.13u w=0.46u m=1
M13 N_13 N_10 N_6 VDD mp15  l=0.13u w=0.26u m=1
M14 N_12 N_5 N_6 VDD mp15  l=0.13u w=0.27u m=1
M15 N_13 N_3 VDD VDD mp15  l=0.13u w=0.26u m=1
M16 N_3 N_6 VDD VDD mp15  l=0.13u w=0.38u m=1
M17 N_10 CK VDD VDD mp15  l=0.13u w=0.58u m=1
M18 N_11 CK VDD VDD mp15  l=0.13u w=0.31u m=1
M19 N_11 N_3 VDD VDD mp15  l=0.13u w=0.31u m=1
M20 ECK N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends tlatncad1
* SPICE INPUT		Tue Jul 31 20:33:41 2018	tlatncad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad2
.subckt tlatncad2 ECK GND VDD CK E
M1 GND N_4 ECK GND mn15  l=0.13u w=0.275u m=1
M2 GND N_4 ECK GND mn15  l=0.13u w=0.275u m=1
M3 N_13 N_7 GND GND mn15  l=0.13u w=0.46u m=1
M4 N_13 CK N_4 GND mn15  l=0.13u w=0.46u m=1
M5 GND N_12 N_8 GND mn15  l=0.13u w=0.19u m=1
M6 N_14 N_12 N_10 GND mn15  l=0.13u w=0.25u m=1
M7 N_15 N_8 N_10 GND mn15  l=0.13u w=0.26u m=1
M8 N_7 N_10 GND GND mn15  l=0.13u w=0.26u m=1
M9 N_15 N_7 GND GND mn15  l=0.13u w=0.26u m=1
M10 N_14 E GND GND mn15  l=0.13u w=0.25u m=1
M11 N_12 CK GND GND mn15  l=0.13u w=0.23u m=1
M12 VDD N_4 ECK VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_4 ECK VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_7 N_4 VDD mp15  l=0.13u w=0.57u m=1
M15 N_4 CK VDD VDD mp15  l=0.13u w=0.57u m=1
M16 N_12 CK VDD VDD mp15  l=0.13u w=0.58u m=1
M17 N_8 N_12 VDD VDD mp15  l=0.13u w=0.48u m=1
M18 N_57 N_8 N_10 VDD mp15  l=0.13u w=0.38u m=1
M19 N_7 N_10 VDD VDD mp15  l=0.13u w=0.4u m=1
M20 N_58 N_7 VDD VDD mp15  l=0.13u w=0.26u m=1
M21 N_58 N_12 N_10 VDD mp15  l=0.13u w=0.26u m=1
M22 N_57 E VDD VDD mp15  l=0.13u w=0.38u m=1
.ends tlatncad2
* SPICE INPUT		Tue Jul 31 20:33:54 2018	tlatncad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatncad4
.subckt tlatncad4 ECK VDD GND CK E
M1 N_25 CK N_6 GND mn15  l=0.13u w=0.38u m=1
M2 GND N_13 N_24 GND mn15  l=0.13u w=0.38u m=1
M3 N_25 N_13 GND GND mn15  l=0.13u w=0.38u m=1
M4 N_6 CK N_24 GND mn15  l=0.13u w=0.38u m=1
M5 ECK N_6 GND GND mn15  l=0.13u w=0.265u m=1
M6 GND N_6 ECK GND mn15  l=0.13u w=0.265u m=1
M7 GND N_6 ECK GND mn15  l=0.13u w=0.265u m=1
M8 GND N_6 ECK GND mn15  l=0.13u w=0.265u m=1
M9 GND CK N_5 GND mn15  l=0.13u w=0.27u m=1
M10 N_27 N_13 GND GND mn15  l=0.13u w=0.26u m=1
M11 GND N_5 N_15 GND mn15  l=0.13u w=0.23u m=1
M12 N_16 N_5 N_26 GND mn15  l=0.13u w=0.26u m=1
M13 GND N_16 N_13 GND mn15  l=0.13u w=0.46u m=1
M14 N_26 E GND GND mn15  l=0.13u w=0.26u m=1
M15 N_27 N_15 N_16 GND mn15  l=0.13u w=0.26u m=1
M16 N_5 CK VDD VDD mp15  l=0.13u w=0.69u m=1
M17 N_6 CK VDD VDD mp15  l=0.13u w=0.49u m=1
M18 VDD N_13 N_6 VDD mp15  l=0.13u w=0.49u m=1
M19 N_6 N_13 VDD VDD mp15  l=0.13u w=0.49u m=1
M20 VDD CK N_6 VDD mp15  l=0.13u w=0.49u m=1
M21 VDD N_6 ECK VDD mp15  l=0.13u w=0.69u m=1
M22 VDD N_6 ECK VDD mp15  l=0.13u w=0.69u m=1
M23 VDD N_6 ECK VDD mp15  l=0.13u w=0.69u m=1
M24 ECK N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_18 N_13 VDD VDD mp15  l=0.13u w=0.26u m=1
M26 N_15 N_5 VDD VDD mp15  l=0.13u w=0.57u m=1
M27 N_13 N_16 VDD VDD mp15  l=0.13u w=0.58u m=1
M28 N_17 E VDD VDD mp15  l=0.13u w=0.48u m=1
M29 N_17 N_15 N_16 VDD mp15  l=0.13u w=0.48u m=1
M30 N_18 N_5 N_16 VDD mp15  l=0.13u w=0.26u m=1
.ends tlatncad4
* SPICE INPUT		Tue Jul 31 20:34:07 2018	tlatnfcad0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatnfcad0
.subckt tlatnfcad0 VDD ECK GND CKN E
M1 GND CKN N_2 GND mn15  l=0.13u w=0.23u m=1
M2 N_11 CKN GND GND mn15  l=0.13u w=0.17u m=1
M3 N_11 N_8 GND GND mn15  l=0.13u w=0.17u m=1
M4 ECK N_11 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_5 N_8 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_22 N_7 N_8 GND mn15  l=0.13u w=0.39u m=1
M7 GND N_2 N_7 GND mn15  l=0.13u w=0.19u m=1
M8 N_22 E GND GND mn15  l=0.13u w=0.39u m=1
M9 N_23 N_2 N_8 GND mn15  l=0.13u w=0.26u m=1
M10 N_23 N_5 GND GND mn15  l=0.13u w=0.26u m=1
M11 VDD CKN N_2 VDD mp15  l=0.13u w=0.57u m=1
M12 N_5 N_8 VDD VDD mp15  l=0.13u w=0.26u m=1
M13 N_7 N_2 VDD VDD mp15  l=0.13u w=0.48u m=1
M14 N_12 E VDD VDD mp15  l=0.13u w=0.58u m=1
M15 N_12 N_2 N_8 VDD mp15  l=0.13u w=0.58u m=1
M16 N_13 N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
M17 N_13 N_7 N_8 VDD mp15  l=0.13u w=0.26u m=1
M18 N_14 CKN N_11 VDD mp15  l=0.13u w=0.69u m=1
M19 N_14 N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 ECK N_11 VDD VDD mp15  l=0.13u w=0.63u m=1
.ends tlatnfcad0
* SPICE INPUT		Tue Jul 31 20:34:20 2018	tlatnfcad1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatnfcad1
.subckt tlatnfcad1 VDD ECK GND CKN E
M1 GND CKN N_2 GND mn15  l=0.13u w=0.23u m=1
M2 N_11 CKN GND GND mn15  l=0.13u w=0.18u m=1
M3 N_11 N_8 GND GND mn15  l=0.13u w=0.18u m=1
M4 ECK N_11 GND GND mn15  l=0.13u w=0.27u m=1
M5 N_5 N_8 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_22 N_7 N_8 GND mn15  l=0.13u w=0.39u m=1
M7 GND N_2 N_7 GND mn15  l=0.13u w=0.19u m=1
M8 N_22 E GND GND mn15  l=0.13u w=0.39u m=1
M9 N_23 N_2 N_8 GND mn15  l=0.13u w=0.26u m=1
M10 N_23 N_5 GND GND mn15  l=0.13u w=0.26u m=1
M11 VDD CKN N_2 VDD mp15  l=0.13u w=0.55u m=1
M12 N_5 N_8 VDD VDD mp15  l=0.13u w=0.26u m=1
M13 N_7 N_2 VDD VDD mp15  l=0.13u w=0.48u m=1
M14 N_12 E VDD VDD mp15  l=0.13u w=0.58u m=1
M15 N_12 N_2 N_8 VDD mp15  l=0.13u w=0.58u m=1
M16 N_13 N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
M17 N_13 N_7 N_8 VDD mp15  l=0.13u w=0.26u m=1
M18 N_14 CKN N_11 VDD mp15  l=0.13u w=0.69u m=1
M19 N_14 N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 ECK N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends tlatnfcad1
* SPICE INPUT		Tue Jul 31 20:34:33 2018	tlatnfcad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatnfcad2
.subckt tlatnfcad2 VDD ECK GND CKN E
M1 N_10 CKN GND GND mn15  l=0.13u w=0.26u m=1
M2 N_11 CKN GND GND mn15  l=0.13u w=0.27u m=1
M3 N_11 N_6 GND GND mn15  l=0.13u w=0.27u m=1
M4 GND N_11 ECK GND mn15  l=0.13u w=0.275u m=1
M5 GND N_11 ECK GND mn15  l=0.13u w=0.275u m=1
M6 GND N_10 N_5 GND mn15  l=0.13u w=0.19u m=1
M7 N_26 E GND GND mn15  l=0.13u w=0.41u m=1
M8 N_26 N_5 N_6 GND mn15  l=0.13u w=0.41u m=1
M9 N_3 N_6 GND GND mn15  l=0.13u w=0.26u m=1
M10 N_27 N_10 N_6 GND mn15  l=0.13u w=0.26u m=1
M11 N_27 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_5 N_10 VDD VDD mp15  l=0.13u w=0.48u m=1
M13 N_13 E VDD VDD mp15  l=0.13u w=0.62u m=1
M14 N_14 N_5 N_6 VDD mp15  l=0.13u w=0.26u m=1
M15 N_3 N_6 VDD VDD mp15  l=0.13u w=0.26u m=1
M16 N_13 N_10 N_6 VDD mp15  l=0.13u w=0.62u m=1
M17 N_14 N_3 VDD VDD mp15  l=0.13u w=0.26u m=1
M18 N_10 CKN VDD VDD mp15  l=0.13u w=0.59u m=1
M19 VDD N_6 N_16 VDD mp15  l=0.13u w=0.54u m=1
M20 N_16 CKN N_11 VDD mp15  l=0.13u w=0.54u m=1
M21 N_11 CKN N_15 VDD mp15  l=0.13u w=0.54u m=1
M22 N_15 N_6 VDD VDD mp15  l=0.13u w=0.54u m=1
M23 VDD N_11 ECK VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_11 ECK VDD mp15  l=0.13u w=0.69u m=1
.ends tlatnfcad2
* SPICE INPUT		Tue Jul 31 20:34:46 2018	tlatnfcad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatnfcad4
.subckt tlatnfcad4 ECK GND VDD CKN E
M1 ECK N_6 GND GND mn15  l=0.13u w=0.265u m=1
M2 ECK N_6 GND GND mn15  l=0.13u w=0.265u m=1
M3 GND N_6 ECK GND mn15  l=0.13u w=0.26u m=1
M4 GND N_6 ECK GND mn15  l=0.13u w=0.26u m=1
M5 N_6 N_13 GND GND mn15  l=0.13u w=0.39u m=1
M6 N_6 CKN GND GND mn15  l=0.13u w=0.39u m=1
M7 GND N_14 N_11 GND mn15  l=0.13u w=0.23u m=1
M8 N_16 E GND GND mn15  l=0.13u w=0.41u m=1
M9 N_16 N_11 N_13 GND mn15  l=0.13u w=0.41u m=1
M10 N_17 N_14 N_13 GND mn15  l=0.13u w=0.26u m=1
M11 N_17 N_10 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_10 N_13 GND GND mn15  l=0.13u w=0.26u m=1
M13 GND CKN N_14 GND mn15  l=0.13u w=0.26u m=1
M14 N_11 N_14 VDD VDD mp15  l=0.13u w=0.58u m=1
M15 N_30 E VDD VDD mp15  l=0.13u w=0.62u m=1
M16 N_31 N_11 N_13 VDD mp15  l=0.13u w=0.26u m=1
M17 N_30 N_14 N_13 VDD mp15  l=0.13u w=0.62u m=1
M18 N_31 N_10 VDD VDD mp15  l=0.13u w=0.26u m=1
M19 N_10 N_13 VDD VDD mp15  l=0.13u w=0.26u m=1
M20 VDD CKN N_14 VDD mp15  l=0.13u w=0.62u m=1
M21 N_33 N_13 VDD VDD mp15  l=0.13u w=0.52u m=1
M22 N_34 CKN N_6 VDD mp15  l=0.13u w=0.52u m=1
M23 N_6 CKN N_33 VDD mp15  l=0.13u w=0.52u m=1
M24 VDD N_13 N_32 VDD mp15  l=0.13u w=0.51u m=1
M25 N_34 N_13 VDD VDD mp15  l=0.13u w=0.52u m=1
M26 N_6 CKN N_32 VDD mp15  l=0.13u w=0.51u m=1
M27 VDD N_6 ECK VDD mp15  l=0.13u w=0.69u m=1
M28 VDD N_6 ECK VDD mp15  l=0.13u w=0.69u m=1
M29 VDD N_6 ECK VDD mp15  l=0.13u w=0.69u m=1
M30 ECK N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends tlatnfcad4
* SPICE INPUT		Tue Jul 31 20:34:59 2018	tlatnftscad0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatnftscad0
.subckt tlatnftscad0 VDD ECK GND E SE CKN
M1 N_4 CKN GND GND mn15  l=0.13u w=0.19u m=1
M2 GND N_4 N_3 GND mn15  l=0.13u w=0.19u m=1
M3 GND SE N_9 GND mn15  l=0.13u w=0.19u m=1
M4 N_9 E GND GND mn15  l=0.13u w=0.19u m=1
M5 N_8 N_3 N_9 GND mn15  l=0.13u w=0.31u m=1
M6 N_52 N_6 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_6 N_8 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_52 N_4 N_8 GND mn15  l=0.13u w=0.26u m=1
M9 ECK N_4 N_53 GND mn15  l=0.13u w=0.26u m=1
M10 GND N_6 N_53 GND mn15  l=0.13u w=0.26u m=1
M11 N_4 CKN VDD VDD mp15  l=0.13u w=0.48u m=1
M12 N_3 N_4 VDD VDD mp15  l=0.13u w=0.48u m=1
M13 N_13 SE VDD VDD mp15  l=0.13u w=0.48u m=1
M14 N_9 E N_13 VDD mp15  l=0.13u w=0.48u m=1
M15 N_9 N_4 N_8 VDD mp15  l=0.13u w=0.48u m=1
M16 N_14 N_3 N_8 VDD mp15  l=0.13u w=0.26u m=1
M17 N_14 N_6 VDD VDD mp15  l=0.13u w=0.26u m=1
M18 N_6 N_8 VDD VDD mp15  l=0.13u w=0.38u m=1
M19 ECK N_4 VDD VDD mp15  l=0.13u w=0.325u m=1
M20 ECK N_6 VDD VDD mp15  l=0.13u w=0.325u m=1
.ends tlatnftscad0
* SPICE INPUT		Tue Jul 31 20:35:12 2018	tlatnftscad1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatnftscad1
.subckt tlatnftscad1 VDD ECK GND E SE CKN
M1 GND N_4 N_3 GND mn15  l=0.13u w=0.19u m=1
M2 N_4 CKN GND GND mn15  l=0.13u w=0.23u m=1
M3 ECK N_4 N_53 GND mn15  l=0.13u w=0.46u m=1
M4 GND N_6 N_53 GND mn15  l=0.13u w=0.46u m=1
M5 GND SE N_8 GND mn15  l=0.13u w=0.23u m=1
M6 N_8 E GND GND mn15  l=0.13u w=0.23u m=1
M7 N_6 N_9 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_54 N_6 GND GND mn15  l=0.13u w=0.26u m=1
M9 N_54 N_4 N_9 GND mn15  l=0.13u w=0.26u m=1
M10 N_9 N_3 N_8 GND mn15  l=0.13u w=0.39u m=1
M11 N_3 N_4 VDD VDD mp15  l=0.13u w=0.48u m=1
M12 N_4 CKN VDD VDD mp15  l=0.13u w=0.6u m=1
M13 N_6 N_9 VDD VDD mp15  l=0.13u w=0.38u m=1
M14 N_14 N_6 VDD VDD mp15  l=0.13u w=0.26u m=1
M15 N_14 N_3 N_9 VDD mp15  l=0.13u w=0.26u m=1
M16 N_9 N_4 N_8 VDD mp15  l=0.13u w=0.57u m=1
M17 N_13 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M18 N_13 E N_8 VDD mp15  l=0.13u w=0.58u m=1
M19 VDD N_4 ECK VDD mp15  l=0.13u w=0.57u m=1
M20 VDD N_6 ECK VDD mp15  l=0.13u w=0.53u m=1
.ends tlatnftscad1
* SPICE INPUT		Tue Jul 31 20:35:26 2018	tlatnftscad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatnftscad2
.subckt tlatnftscad2 GND ECK VDD E SE CKN
M1 N_4 CKN GND GND mn15  l=0.13u w=0.27u m=1
M2 GND N_4 N_2 GND mn15  l=0.13u w=0.23u m=1
M3 GND SE N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 E GND GND mn15  l=0.13u w=0.26u m=1
M5 N_16 N_4 ECK GND mn15  l=0.13u w=0.46u m=1
M6 N_16 N_12 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_12 N_15 GND mn15  l=0.13u w=0.46u m=1
M8 ECK N_4 N_15 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 N_13 GND GND mn15  l=0.13u w=0.35u m=1
M10 N_6 N_2 N_13 GND mn15  l=0.13u w=0.35u m=1
M11 N_17 N_12 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_17 N_4 N_13 GND mn15  l=0.13u w=0.26u m=1
M13 N_4 CKN VDD VDD mp15  l=0.13u w=0.69u m=1
M14 N_2 N_4 VDD VDD mp15  l=0.13u w=0.58u m=1
M15 N_28 SE VDD VDD mp15  l=0.13u w=0.61u m=1
M16 N_12 N_13 VDD VDD mp15  l=0.13u w=0.52u m=1
M17 N_29 N_2 N_13 VDD mp15  l=0.13u w=0.26u m=1
M18 N_28 E N_6 VDD mp15  l=0.13u w=0.61u m=1
M19 N_29 N_12 VDD VDD mp15  l=0.13u w=0.26u m=1
M20 N_13 N_4 N_6 VDD mp15  l=0.13u w=0.53u m=1
M21 ECK N_4 VDD VDD mp15  l=0.13u w=0.56u m=1
M22 VDD N_12 ECK VDD mp15  l=0.13u w=0.57u m=1
M23 ECK N_12 VDD VDD mp15  l=0.13u w=0.57u m=1
M24 VDD N_4 ECK VDD mp15  l=0.13u w=0.57u m=1
.ends tlatnftscad2
* SPICE INPUT		Tue Jul 31 20:35:39 2018	tlatnftscad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatnftscad4
.subckt tlatnftscad4 VDD ECK GND SE E CKN
M1 N_12 N_2 GND GND mn15  l=0.13u w=0.3u m=1
M2 N_12 N_9 GND GND mn15  l=0.13u w=0.305u m=1
M3 N_12 N_9 GND GND mn15  l=0.13u w=0.3u m=1
M4 N_12 N_2 GND GND mn15  l=0.13u w=0.305u m=1
M5 N_12 N_2 GND GND mn15  l=0.13u w=0.305u m=1
M6 N_12 N_9 GND GND mn15  l=0.13u w=0.305u m=1
M7 GND N_12 ECK GND mn15  l=0.13u w=0.265u m=1
M8 GND N_12 ECK GND mn15  l=0.13u w=0.265u m=1
M9 ECK N_12 GND GND mn15  l=0.13u w=0.265u m=1
M10 GND N_12 ECK GND mn15  l=0.13u w=0.265u m=1
M11 N_4 CKN GND GND mn15  l=0.13u w=0.27u m=1
M12 N_2 N_4 GND GND mn15  l=0.13u w=0.27u m=1
M13 GND SE N_8 GND mn15  l=0.13u w=0.26u m=1
M14 N_8 E GND GND mn15  l=0.13u w=0.26u m=1
M15 N_9 N_2 N_8 GND mn15  l=0.13u w=0.32u m=1
M16 N_33 N_4 N_9 GND mn15  l=0.13u w=0.26u m=1
M17 N_33 N_5 GND GND mn15  l=0.13u w=0.26u m=1
M18 N_5 N_9 GND GND mn15  l=0.13u w=0.26u m=1
M19 N_4 CKN VDD VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_4 N_2 VDD mp15  l=0.13u w=0.69u m=1
M21 N_18 SE VDD VDD mp15  l=0.13u w=0.62u m=1
M22 N_18 E N_8 VDD mp15  l=0.13u w=0.62u m=1
M23 N_19 N_2 N_9 VDD mp15  l=0.13u w=0.26u m=1
M24 N_9 N_4 N_8 VDD mp15  l=0.13u w=0.53u m=1
M25 N_19 N_5 VDD VDD mp15  l=0.13u w=0.26u m=1
M26 VDD N_9 N_5 VDD mp15  l=0.13u w=0.26u m=1
M27 N_20 N_2 N_12 VDD mp15  l=0.13u w=0.61u m=1
M28 N_21 N_9 VDD VDD mp15  l=0.13u w=0.61u m=1
M29 N_20 N_9 VDD VDD mp15  l=0.13u w=0.61u m=1
M30 N_22 N_2 N_12 VDD mp15  l=0.13u w=0.61u m=1
M31 N_12 N_2 N_21 VDD mp15  l=0.13u w=0.61u m=1
M32 N_22 N_9 VDD VDD mp15  l=0.13u w=0.61u m=1
M33 VDD N_12 ECK VDD mp15  l=0.13u w=0.69u m=1
M34 VDD N_12 ECK VDD mp15  l=0.13u w=0.69u m=1
M35 VDD N_12 ECK VDD mp15  l=0.13u w=0.69u m=1
M36 ECK N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends tlatnftscad4
* SPICE INPUT		Tue Jul 31 20:35:52 2018	tlatntscad0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad0
.subckt tlatntscad0 VDD ECK GND E SE CK
M1 N_8 E GND GND mn15  l=0.13u w=0.19u m=1
M2 GND SE N_8 GND mn15  l=0.13u w=0.19u m=1
M3 N_8 N_4 N_9 GND mn15  l=0.13u w=0.32u m=1
M4 N_55 N_6 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_6 N_9 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_55 N_3 N_9 GND mn15  l=0.13u w=0.26u m=1
M7 GND N_4 N_3 GND mn15  l=0.13u w=0.19u m=1
M8 N_4 CK GND GND mn15  l=0.13u w=0.23u m=1
M9 GND N_9 ECK GND mn15  l=0.13u w=0.26u m=1
M10 ECK N_4 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_3 N_4 VDD VDD mp15  l=0.13u w=0.48u m=1
M12 N_4 CK VDD VDD mp15  l=0.13u w=0.58u m=1
M13 N_13 N_4 N_9 VDD mp15  l=0.13u w=0.26u m=1
M14 N_12 E N_8 VDD mp15  l=0.13u w=0.48u m=1
M15 N_13 N_6 VDD VDD mp15  l=0.13u w=0.26u m=1
M16 N_12 SE VDD VDD mp15  l=0.13u w=0.48u m=1
M17 N_6 N_9 VDD VDD mp15  l=0.13u w=0.26u m=1
M18 N_9 N_3 N_8 VDD mp15  l=0.13u w=0.48u m=1
M19 VDD N_9 N_14 VDD mp15  l=0.13u w=0.69u m=1
M20 ECK N_4 N_14 VDD mp15  l=0.13u w=0.69u m=1
.ends tlatntscad0
* SPICE INPUT		Tue Jul 31 20:36:05 2018	tlatntscad1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad1
.subckt tlatntscad1 GND ECK VDD E SE CK
M1 N_15 N_12 GND GND mn15  l=0.13u w=0.26u m=1
M2 ECK N_4 GND GND mn15  l=0.13u w=0.27u m=1
M3 N_15 N_5 N_4 GND mn15  l=0.13u w=0.26u m=1
M4 N_7 CK GND GND mn15  l=0.13u w=0.19u m=1
M5 GND N_7 N_5 GND mn15  l=0.13u w=0.23u m=1
M6 GND SE N_9 GND mn15  l=0.13u w=0.23u m=1
M7 N_9 E GND GND mn15  l=0.13u w=0.23u m=1
M8 N_16 N_5 N_14 GND mn15  l=0.13u w=0.26u m=1
M9 N_14 N_7 N_9 GND mn15  l=0.13u w=0.35u m=1
M10 N_16 N_12 GND GND mn15  l=0.13u w=0.26u m=1
M11 N_12 N_14 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_7 CK VDD VDD mp15  l=0.13u w=0.48u m=1
M13 VDD N_7 N_5 VDD mp15  l=0.13u w=0.58u m=1
M14 N_57 SE VDD VDD mp15  l=0.13u w=0.58u m=1
M15 N_14 N_5 N_9 VDD mp15  l=0.13u w=0.52u m=1
M16 N_57 E N_9 VDD mp15  l=0.13u w=0.58u m=1
M17 N_58 N_7 N_14 VDD mp15  l=0.13u w=0.26u m=1
M18 N_58 N_12 VDD VDD mp15  l=0.13u w=0.26u m=1
M19 VDD N_14 N_12 VDD mp15  l=0.13u w=0.38u m=1
M20 N_4 N_12 VDD VDD mp15  l=0.13u w=0.325u m=1
M21 ECK N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M22 N_4 N_5 VDD VDD mp15  l=0.13u w=0.325u m=1
.ends tlatntscad1
* SPICE INPUT		Tue Jul 31 20:36:18 2018	tlatntscad2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad2
.subckt tlatntscad2 GND ECK VDD E SE CK
M1 GND N_5 N_2 GND mn15  l=0.13u w=0.34u m=1
M2 N_16 N_2 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_16 N_7 N_5 GND mn15  l=0.13u w=0.26u m=1
M4 N_5 N_8 N_4 GND mn15  l=0.13u w=0.27u m=1
M5 N_8 CK GND GND mn15  l=0.13u w=0.21u m=1
M6 N_7 N_8 GND GND mn15  l=0.13u w=0.26u m=1
M7 GND N_11 ECK GND mn15  l=0.13u w=0.275u m=1
M8 GND N_11 ECK GND mn15  l=0.13u w=0.275u m=1
M9 N_17 N_2 GND GND mn15  l=0.13u w=0.43u m=1
M10 N_17 N_7 N_11 GND mn15  l=0.13u w=0.43u m=1
M11 GND SE N_4 GND mn15  l=0.13u w=0.26u m=1
M12 N_4 E GND GND mn15  l=0.13u w=0.26u m=1
M13 N_61 SE VDD VDD mp15  l=0.13u w=0.61u m=1
M14 N_61 E N_4 VDD mp15  l=0.13u w=0.61u m=1
M15 N_2 N_5 VDD VDD mp15  l=0.13u w=0.53u m=1
M16 N_62 N_2 VDD VDD mp15  l=0.13u w=0.26u m=1
M17 N_5 N_7 N_4 VDD mp15  l=0.13u w=0.53u m=1
M18 N_62 N_8 N_5 VDD mp15  l=0.13u w=0.26u m=1
M19 VDD N_11 ECK VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_11 ECK VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_2 N_11 VDD mp15  l=0.13u w=0.53u m=1
M22 N_11 N_7 VDD VDD mp15  l=0.13u w=0.53u m=1
M23 N_8 CK VDD VDD mp15  l=0.13u w=0.53u m=1
M24 N_7 N_8 VDD VDD mp15  l=0.13u w=0.63u m=1
.ends tlatntscad2
* SPICE INPUT		Tue Jul 31 20:36:31 2018	tlatntscad4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=tlatntscad4
.subckt tlatntscad4 GND ECK VDD E SE CK
M1 N_4 CK GND GND mn15  l=0.13u w=0.26u m=1
M2 N_3 N_4 GND GND mn15  l=0.13u w=0.27u m=1
M3 GND SE N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_6 E GND GND mn15  l=0.13u w=0.26u m=1
M5 N_11 N_4 N_6 GND mn15  l=0.13u w=0.35u m=1
M6 N_19 N_9 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_9 N_11 GND GND mn15  l=0.13u w=0.35u m=1
M8 N_19 N_3 N_11 GND mn15  l=0.13u w=0.26u m=1
M9 N_20 N_9 GND GND mn15  l=0.13u w=0.46u m=1
M10 N_21 N_3 N_15 GND mn15  l=0.13u w=0.46u m=1
M11 N_15 N_3 N_20 GND mn15  l=0.13u w=0.46u m=1
M12 N_21 N_9 GND GND mn15  l=0.13u w=0.46u m=1
M13 ECK N_15 GND GND mn15  l=0.13u w=0.265u m=1
M14 ECK N_15 GND GND mn15  l=0.13u w=0.265u m=1
M15 GND N_15 ECK GND mn15  l=0.13u w=0.26u m=1
M16 GND N_15 ECK GND mn15  l=0.13u w=0.26u m=1
M17 N_4 CK VDD VDD mp15  l=0.13u w=0.63u m=1
M18 N_3 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_82 SE VDD VDD mp15  l=0.13u w=0.61u m=1
M20 N_82 E N_6 VDD mp15  l=0.13u w=0.61u m=1
M21 N_83 N_4 N_11 VDD mp15  l=0.13u w=0.26u m=1
M22 N_83 N_9 VDD VDD mp15  l=0.13u w=0.26u m=1
M23 VDD N_11 N_9 VDD mp15  l=0.13u w=0.35u m=1
M24 N_9 N_11 VDD VDD mp15  l=0.13u w=0.35u m=1
M25 N_11 N_3 N_6 VDD mp15  l=0.13u w=0.52u m=1
M26 N_15 N_9 VDD VDD mp15  l=0.13u w=0.57u m=1
M27 N_15 N_3 VDD VDD mp15  l=0.13u w=0.57u m=1
M28 VDD N_3 N_15 VDD mp15  l=0.13u w=0.57u m=1
M29 VDD N_9 N_15 VDD mp15  l=0.13u w=0.57u m=1
M30 VDD N_15 ECK VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_15 ECK VDD mp15  l=0.13u w=0.69u m=1
M32 VDD N_15 ECK VDD mp15  l=0.13u w=0.69u m=1
M33 ECK N_15 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends tlatntscad4
* SPICE INPUT		Tue Jul 31 20:36:45 2018	xn02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d0
.subckt xn02d0 GND Y VDD B A
M1 N_7 B GND GND mn15  l=0.13u w=0.3u m=1
M2 N_8 N_7 GND GND mn15  l=0.13u w=0.23u m=1
M3 N_7 A N_6 GND mn15  l=0.13u w=0.26u m=1
M4 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M5 Y N_6 GND GND mn15  l=0.13u w=0.26u m=1
M6 N_8 N_5 N_6 GND mn15  l=0.13u w=0.23u m=1
M7 N_7 B VDD VDD mp15  l=0.13u w=0.45u m=1
M8 N_14 N_7 VDD VDD mp15  l=0.13u w=0.33u m=1
M9 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M10 N_6 A N_14 VDD mp15  l=0.13u w=0.33u m=1
M11 Y N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M12 N_7 N_5 N_6 VDD mp15  l=0.13u w=0.26u m=1
.ends xn02d0
* SPICE INPUT		Tue Jul 31 20:36:59 2018	xn02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d1
.subckt xn02d1 GND Y VDD B A
M1 N_8 N_7 GND GND mn15  l=0.13u w=0.3u m=1
M2 N_8 N_4 N_6 GND mn15  l=0.13u w=0.3u m=1
M3 N_7 A N_6 GND mn15  l=0.13u w=0.3u m=1
M4 GND A N_4 GND mn15  l=0.13u w=0.26u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.33u m=1
M6 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M7 N_32 N_7 VDD VDD mp15  l=0.13u w=0.45u m=1
M8 N_7 N_4 N_6 VDD mp15  l=0.13u w=0.3u m=1
M9 N_6 A N_32 VDD mp15  l=0.13u w=0.45u m=1
M10 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
M11 N_7 B VDD VDD mp15  l=0.13u w=0.5u m=1
M12 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends xn02d1
* SPICE INPUT		Tue Jul 31 20:37:12 2018	xn02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d2
.subckt xn02d2 GND Y VDD A B
M1 GND B N_2 GND mn15  l=0.13u w=0.41u m=1
M2 N_10 N_2 GND GND mn15  l=0.13u w=0.41u m=1
M3 N_10 N_8 N_3 GND mn15  l=0.13u w=0.41u m=1
M4 N_3 A N_2 GND mn15  l=0.13u w=0.39u m=1
M5 GND A N_8 GND mn15  l=0.13u w=0.26u m=1
M6 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M7 GND N_3 Y GND mn15  l=0.13u w=0.46u m=1
M8 VDD B N_2 VDD mp15  l=0.13u w=0.63u m=1
M9 N_16 N_2 VDD VDD mp15  l=0.13u w=0.63u m=1
M10 N_2 N_8 N_3 VDD mp15  l=0.13u w=0.31u m=1
M11 N_16 A N_3 VDD mp15  l=0.13u w=0.63u m=1
M12 VDD A N_8 VDD mp15  l=0.13u w=0.4u m=1
M13 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
M14 VDD N_3 Y VDD mp15  l=0.13u w=0.69u m=1
.ends xn02d2
* SPICE INPUT		Tue Jul 31 20:37:25 2018	xn02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02d4
.subckt xn02d4 Y GND VDD B A
M1 N_4 A N_2 GND mn15  l=0.13u w=0.37u m=1
M2 N_4 A N_2 GND mn15  l=0.13u w=0.37u m=1
M3 GND A N_8 GND mn15  l=0.13u w=0.19u m=1
M4 N_8 A GND GND mn15  l=0.13u w=0.19u m=1
M5 N_10 N_8 N_2 GND mn15  l=0.13u w=0.53u m=1
M6 N_2 N_8 N_10 GND mn15  l=0.13u w=0.27u m=1
M7 N_10 N_4 GND GND mn15  l=0.13u w=0.35u m=1
M8 GND N_4 N_10 GND mn15  l=0.13u w=0.45u m=1
M9 GND B N_4 GND mn15  l=0.13u w=0.42u m=1
M10 N_4 B GND GND mn15  l=0.13u w=0.42u m=1
M11 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M14 GND N_2 Y GND mn15  l=0.13u w=0.46u m=1
M15 N_4 N_8 N_2 VDD mp15  l=0.13u w=0.46u m=1
M16 N_4 N_8 N_2 VDD mp15  l=0.13u w=0.46u m=1
M17 N_8 A VDD VDD mp15  l=0.13u w=0.6u m=1
M18 N_2 A N_20 VDD mp15  l=0.13u w=0.62u m=1
M19 N_2 A N_20 VDD mp15  l=0.13u w=0.62u m=1
M20 N_20 N_4 VDD VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_4 N_20 VDD mp15  l=0.13u w=0.55u m=1
M22 N_4 B VDD VDD mp15  l=0.13u w=0.63u m=1
M23 N_4 B VDD VDD mp15  l=0.13u w=0.63u m=1
M24 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M25 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M26 VDD N_2 Y VDD mp15  l=0.13u w=0.69u m=1
M27 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends xn02d4
* SPICE INPUT		Tue Jul 31 20:37:39 2018	xn02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn02dm
.subckt xn02dm GND Y VDD B A
M1 N_8 N_7 GND GND mn15  l=0.13u w=0.23u m=1
M2 N_7 A N_6 GND mn15  l=0.13u w=0.26u m=1
M3 N_5 A GND GND mn15  l=0.13u w=0.26u m=1
M4 N_7 B GND GND mn15  l=0.13u w=0.3u m=1
M5 Y N_6 GND GND mn15  l=0.13u w=0.36u m=1
M6 N_8 N_5 N_6 GND mn15  l=0.13u w=0.23u m=1
M7 N_14 N_7 VDD VDD mp15  l=0.13u w=0.33u m=1
M8 N_5 A VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_6 A N_14 VDD mp15  l=0.13u w=0.33u m=1
M10 N_7 B VDD VDD mp15  l=0.13u w=0.45u m=1
M11 Y N_6 VDD VDD mp15  l=0.13u w=0.55u m=1
M12 N_7 N_5 N_6 VDD mp15  l=0.13u w=0.26u m=1
.ends xn02dm
* SPICE INPUT		Tue Jul 31 20:37:52 2018	xn03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d0
.subckt xn03d0 GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_13 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_13 A N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_11 GND GND mn15  l=0.13u w=0.26u m=1
M8 N_12 C GND GND mn15  l=0.13u w=0.28u m=1
M9 N_14 N_12 GND GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 N_11 GND mn15  l=0.13u w=0.28u m=1
M11 N_12 N_3 N_11 GND mn15  l=0.13u w=0.28u m=1
M12 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M13 N_23 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_7 A N_6 VDD mp15  l=0.13u w=0.28u m=1
M15 N_23 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_3 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 Y N_11 VDD VDD mp15  l=0.13u w=0.4u m=1
M19 N_12 C VDD VDD mp15  l=0.13u w=0.4u m=1
M20 N_12 N_6 N_11 VDD mp15  l=0.13u w=0.28u m=1
M21 N_24 N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 N_24 N_3 N_11 VDD mp15  l=0.13u w=0.4u m=1
.ends xn03d0
* SPICE INPUT		Tue Jul 31 20:38:05 2018	xn03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d1
.subckt xn03d1 GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_13 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_13 A N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_11 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_12 C GND GND mn15  l=0.13u w=0.28u m=1
M9 N_14 N_12 GND GND mn15  l=0.13u w=0.3u m=1
M10 N_14 N_6 N_11 GND mn15  l=0.13u w=0.3u m=1
M11 N_12 N_3 N_11 GND mn15  l=0.13u w=0.28u m=1
M12 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M13 N_23 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_7 A N_6 VDD mp15  l=0.13u w=0.28u m=1
M15 N_23 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_3 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 Y N_11 VDD VDD mp15  l=0.13u w=0.69u m=1
M19 N_12 C VDD VDD mp15  l=0.13u w=0.42u m=1
M20 N_12 N_6 N_11 VDD mp15  l=0.13u w=0.28u m=1
M21 N_24 N_12 VDD VDD mp15  l=0.13u w=0.45u m=1
M22 N_24 N_3 N_11 VDD mp15  l=0.13u w=0.45u m=1
.ends xn03d1
* SPICE INPUT		Tue Jul 31 20:38:18 2018	xn03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d2
.subckt xn03d2 GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_14 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_14 A N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M7 N_15 N_12 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_15 N_6 N_11 GND mn15  l=0.13u w=0.46u m=1
M9 N_12 N_3 N_11 GND mn15  l=0.13u w=0.45u m=1
M10 GND C N_12 GND mn15  l=0.13u w=0.42u m=1
M11 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M12 GND N_11 Y GND mn15  l=0.13u w=0.46u m=1
M13 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M14 N_60 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M15 N_7 A N_6 VDD mp15  l=0.13u w=0.36u m=1
M16 N_60 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M17 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_3 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M19 N_61 N_12 VDD VDD mp15  l=0.13u w=0.69u m=1
M20 N_61 N_3 N_11 VDD mp15  l=0.13u w=0.69u m=1
M21 N_12 N_6 N_11 VDD mp15  l=0.13u w=0.57u m=1
M22 N_12 C VDD VDD mp15  l=0.13u w=0.62u m=1
M23 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
M24 VDD N_11 Y VDD mp15  l=0.13u w=0.69u m=1
.ends xn03d2
* SPICE INPUT		Tue Jul 31 20:38:31 2018	xn03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03d4
.subckt xn03d4 GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_18 N_7 GND GND mn15  l=0.13u w=0.38u m=1
M3 N_18 A N_6 GND mn15  l=0.13u w=0.38u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.38u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.33u m=1
M7 N_10 N_6 N_19 GND mn15  l=0.13u w=0.32u m=1
M8 N_10 N_6 N_20 GND mn15  l=0.13u w=0.32u m=1
M9 GND N_14 N_20 GND mn15  l=0.13u w=0.44u m=1
M10 N_19 N_14 GND GND mn15  l=0.13u w=0.2u m=1
M11 N_14 N_3 N_10 GND mn15  l=0.13u w=0.5u m=1
M12 GND C N_14 GND mn15  l=0.13u w=0.46u m=1
M13 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M14 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M15 Y N_10 GND GND mn15  l=0.13u w=0.46u m=1
M16 GND N_10 Y GND mn15  l=0.13u w=0.46u m=1
M17 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M18 N_79 N_7 VDD VDD mp15  l=0.13u w=0.57u m=1
M19 N_79 N_4 N_6 VDD mp15  l=0.13u w=0.57u m=1
M20 N_7 A N_6 VDD mp15  l=0.13u w=0.38u m=1
M21 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M22 N_3 N_6 VDD VDD mp15  l=0.13u w=0.52u m=1
M23 N_81 N_3 N_10 VDD mp15  l=0.13u w=0.425u m=1
M24 N_10 N_3 N_80 VDD mp15  l=0.13u w=0.425u m=1
M25 N_80 N_14 VDD VDD mp15  l=0.13u w=0.53u m=1
M26 N_81 N_14 VDD VDD mp15  l=0.13u w=0.32u m=1
M27 N_14 N_6 N_10 VDD mp15  l=0.13u w=0.5u m=1
M28 N_14 C VDD VDD mp15  l=0.13u w=0.66u m=1
M29 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M30 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M31 VDD N_10 Y VDD mp15  l=0.13u w=0.69u m=1
M32 Y N_10 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends xn03d4
* SPICE INPUT		Tue Jul 31 20:38:44 2018	xn03dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xn03dm
.subckt xn03dm GND Y VDD C B A
M1 GND A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_13 N_7 GND GND mn15  l=0.13u w=0.28u m=1
M3 N_13 A N_6 GND mn15  l=0.13u w=0.28u m=1
M4 N_7 N_4 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_7 B GND GND mn15  l=0.13u w=0.28u m=1
M6 N_3 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M7 Y N_11 GND GND mn15  l=0.13u w=0.36u m=1
M8 N_12 C GND GND mn15  l=0.13u w=0.28u m=1
M9 N_14 N_12 GND GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 N_11 GND mn15  l=0.13u w=0.28u m=1
M11 N_12 N_3 N_11 GND mn15  l=0.13u w=0.28u m=1
M12 VDD A N_4 VDD mp15  l=0.13u w=0.4u m=1
M13 N_23 N_7 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_7 A N_6 VDD mp15  l=0.13u w=0.28u m=1
M15 N_23 N_4 N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 N_7 B VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_3 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 Y N_11 VDD VDD mp15  l=0.13u w=0.55u m=1
M19 N_12 C VDD VDD mp15  l=0.13u w=0.4u m=1
M20 N_12 N_6 N_11 VDD mp15  l=0.13u w=0.28u m=1
M21 N_24 N_12 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 N_24 N_3 N_11 VDD mp15  l=0.13u w=0.4u m=1
.ends xn03dm
* SPICE INPUT		Tue Jul 31 20:38:58 2018	xr02d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d0
.subckt xr02d0 GND Y A VDD B
M1 GND B N_3 GND mn15  l=0.13u w=0.28u m=1
M2 N_9 N_3 GND GND mn15  l=0.13u w=0.26u m=1
M3 N_3 N_8 N_2 GND mn15  l=0.13u w=0.26u m=1
M4 N_9 A N_2 GND mn15  l=0.13u w=0.26u m=1
M5 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M6 Y N_2 GND GND mn15  l=0.13u w=0.26u m=1
M7 N_3 B VDD VDD mp15  l=0.13u w=0.42u m=1
M8 N_15 N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_15 N_8 N_2 VDD mp15  l=0.13u w=0.4u m=1
M10 N_2 A N_3 VDD mp15  l=0.13u w=0.26u m=1
M11 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M12 Y N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr02d0
* SPICE INPUT		Tue Jul 31 20:39:12 2018	xr02d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d1
.subckt xr02d1 GND Y A VDD B
M1 GND B N_3 GND mn15  l=0.13u w=0.32u m=1
M2 N_9 N_3 GND GND mn15  l=0.13u w=0.32u m=1
M3 N_3 N_8 N_2 GND mn15  l=0.13u w=0.28u m=1
M4 N_9 A N_2 GND mn15  l=0.13u w=0.32u m=1
M5 Y N_2 GND GND mn15  l=0.13u w=0.46u m=1
M6 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M7 VDD B N_3 VDD mp15  l=0.13u w=0.52u m=1
M8 N_34 N_3 VDD VDD mp15  l=0.13u w=0.52u m=1
M9 N_34 N_8 N_2 VDD mp15  l=0.13u w=0.52u m=1
M10 N_2 A N_3 VDD mp15  l=0.13u w=0.42u m=1
M11 Y N_2 VDD VDD mp15  l=0.13u w=0.69u m=1
M12 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr02d1
* SPICE INPUT		Tue Jul 31 20:39:24 2018	xr02d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d2
.subckt xr02d2 Y GND VDD A B
M1 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M2 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M3 GND A N_4 GND mn15  l=0.13u w=0.26u m=1
M4 GND B N_7 GND mn15  l=0.13u w=0.41u m=1
M5 N_10 N_7 GND GND mn15  l=0.13u w=0.39u m=1
M6 N_7 N_4 N_6 GND mn15  l=0.13u w=0.32u m=1
M7 N_10 A N_6 GND mn15  l=0.13u w=0.39u m=1
M8 N_7 B VDD VDD mp15  l=0.13u w=0.63u m=1
M9 N_38 N_7 VDD VDD mp15  l=0.13u w=0.54u m=1
M10 N_38 N_4 N_6 VDD mp15  l=0.13u w=0.54u m=1
M11 N_6 A N_7 VDD mp15  l=0.13u w=0.46u m=1
M12 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M13 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M14 N_4 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr02d2
* SPICE INPUT		Tue Jul 31 20:39:37 2018	xr02d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02d4
.subckt xr02d4 GND Y VDD A B
M1 N_5 B GND GND mn15  l=0.13u w=0.42u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.42u m=1
M3 N_17 N_5 GND GND mn15  l=0.13u w=0.51u m=1
M4 N_18 N_5 GND GND mn15  l=0.13u w=0.27u m=1
M5 N_17 A N_6 GND mn15  l=0.13u w=0.51u m=1
M6 N_18 A N_6 GND mn15  l=0.13u w=0.27u m=1
M7 N_6 N_13 N_5 GND mn15  l=0.13u w=0.26u m=1
M8 N_5 N_13 N_6 GND mn15  l=0.13u w=0.26u m=1
M9 N_5 N_13 N_6 GND mn15  l=0.13u w=0.24u m=1
M10 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M11 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M12 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M13 GND N_6 Y GND mn15  l=0.13u w=0.46u m=1
M14 GND A N_13 GND mn15  l=0.13u w=0.41u m=1
M15 VDD B N_5 VDD mp15  l=0.13u w=0.66u m=1
M16 VDD B N_5 VDD mp15  l=0.13u w=0.59u m=1
M17 VDD N_5 N_23 VDD mp15  l=0.13u w=0.59u m=1
M18 VDD N_5 N_23 VDD mp15  l=0.13u w=0.59u m=1
M19 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M20 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M21 VDD N_6 Y VDD mp15  l=0.13u w=0.69u m=1
M22 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M23 N_13 A VDD VDD mp15  l=0.13u w=0.61u m=1
M24 N_23 N_13 N_6 VDD mp15  l=0.13u w=0.59u m=1
M25 N_23 N_13 N_6 VDD mp15  l=0.13u w=0.59u m=1
M26 N_6 A N_5 VDD mp15  l=0.13u w=0.52u m=1
M27 N_6 A N_5 VDD mp15  l=0.13u w=0.42u m=1
.ends xr02d4
* SPICE INPUT		Tue Jul 31 20:39:49 2018	xr02dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr02dm
.subckt xr02dm VDD Y GND A B
M1 N_8 A GND GND mn15  l=0.13u w=0.26u m=1
M2 Y N_3 GND GND mn15  l=0.13u w=0.36u m=1
M3 GND B N_2 GND mn15  l=0.13u w=0.28u m=1
M4 N_14 N_2 GND GND mn15  l=0.13u w=0.26u m=1
M5 N_3 N_8 N_2 GND mn15  l=0.13u w=0.3u m=1
M6 N_14 A N_3 GND mn15  l=0.13u w=0.26u m=1
M7 N_2 B VDD VDD mp15  l=0.13u w=0.42u m=1
M8 N_9 N_2 VDD VDD mp15  l=0.13u w=0.4u m=1
M9 N_9 N_8 N_3 VDD mp15  l=0.13u w=0.4u m=1
M10 N_3 A N_2 VDD mp15  l=0.13u w=0.3u m=1
M11 N_8 A VDD VDD mp15  l=0.13u w=0.4u m=1
M12 Y N_3 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends xr02dm
* SPICE INPUT		Tue Jul 31 20:40:02 2018	xr03d0
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d0
.subckt xr03d0 GND Y VDD B A C
M1 N_3 A GND GND mn15  l=0.13u w=0.28u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.28u m=1
M3 N_15 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_15 N_3 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_5 A N_6 GND mn15  l=0.13u w=0.28u m=1
M6 GND C N_9 GND mn15  l=0.13u w=0.28u m=1
M7 N_16 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_9 N_14 N_8 GND mn15  l=0.13u w=0.28u m=1
M9 N_16 N_6 N_8 GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M11 Y N_8 GND GND mn15  l=0.13u w=0.26u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_58 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.28u m=1
M15 N_58 A N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 VDD C N_9 VDD mp15  l=0.13u w=0.4u m=1
M17 N_59 N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_59 N_14 N_8 VDD mp15  l=0.13u w=0.4u m=1
M19 N_9 N_6 N_8 VDD mp15  l=0.13u w=0.28u m=1
M20 N_3 A VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_14 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 Y N_8 VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr03d0
* SPICE INPUT		Tue Jul 31 20:40:15 2018	xr03d1
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d1
.subckt xr03d1 GND Y VDD B A C
M1 N_3 A GND GND mn15  l=0.13u w=0.28u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.28u m=1
M3 N_15 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_15 N_3 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_5 A N_6 GND mn15  l=0.13u w=0.28u m=1
M6 GND C N_9 GND mn15  l=0.13u w=0.28u m=1
M7 N_16 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_9 N_14 N_8 GND mn15  l=0.13u w=0.28u m=1
M9 N_16 N_6 N_8 GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M11 Y N_8 GND GND mn15  l=0.13u w=0.46u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_60 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.28u m=1
M15 N_60 A N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 VDD C N_9 VDD mp15  l=0.13u w=0.4u m=1
M17 N_61 N_9 VDD VDD mp15  l=0.13u w=0.42u m=1
M18 N_61 N_14 N_8 VDD mp15  l=0.13u w=0.42u m=1
M19 N_9 N_6 N_8 VDD mp15  l=0.13u w=0.28u m=1
M20 N_3 A VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_14 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 Y N_8 VDD VDD mp15  l=0.13u w=0.69u m=1
.ends xr03d1
* SPICE INPUT		Tue Jul 31 20:40:28 2018	xr03d2
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d2
.subckt xr03d2 VDD Y GND B A C
M1 N_3 A N_4 GND mn15  l=0.13u w=0.28u m=1
M2 N_23 N_11 N_4 GND mn15  l=0.13u w=0.28u m=1
M3 N_23 N_3 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_3 B GND GND mn15  l=0.13u w=0.28u m=1
M5 GND N_4 N_13 GND mn15  l=0.13u w=0.28u m=1
M6 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M7 Y N_6 GND GND mn15  l=0.13u w=0.46u m=1
M8 N_11 A GND GND mn15  l=0.13u w=0.28u m=1
M9 GND C N_7 GND mn15  l=0.13u w=0.42u m=1
M10 N_24 N_7 GND GND mn15  l=0.13u w=0.45u m=1
M11 N_7 N_13 N_6 GND mn15  l=0.13u w=0.21u m=1
M12 N_6 N_13 N_7 GND mn15  l=0.13u w=0.2u m=1
M13 N_24 N_4 N_6 GND mn15  l=0.13u w=0.45u m=1
M14 N_15 A N_4 VDD mp15  l=0.13u w=0.4u m=1
M15 N_3 N_11 N_4 VDD mp15  l=0.13u w=0.33u m=1
M16 N_15 N_3 VDD VDD mp15  l=0.13u w=0.4u m=1
M17 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M18 VDD C N_7 VDD mp15  l=0.13u w=0.62u m=1
M19 N_16 N_7 VDD VDD mp15  l=0.13u w=0.67u m=1
M20 N_16 N_13 N_6 VDD mp15  l=0.13u w=0.67u m=1
M21 N_7 N_4 N_6 VDD mp15  l=0.13u w=0.56u m=1
M22 N_13 N_4 VDD VDD mp15  l=0.13u w=0.4u m=1
M23 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_6 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 N_11 A VDD VDD mp15  l=0.13u w=0.4u m=1
.ends xr03d2
* SPICE INPUT		Tue Jul 31 20:40:41 2018	xr03d4
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03d4
.subckt xr03d4 VDD Y C A B GND
M1 N_3 B GND GND mn15  l=0.13u w=0.28u m=1
M2 N_80 N_3 GND GND mn15  l=0.13u w=0.38u m=1
M3 N_80 N_7 N_5 GND mn15  l=0.13u w=0.38u m=1
M4 N_3 A N_5 GND mn15  l=0.13u w=0.36u m=1
M5 N_7 A GND GND mn15  l=0.13u w=0.28u m=1
M6 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M7 GND N_13 Y GND mn15  l=0.13u w=0.46u m=1
M8 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M9 Y N_13 GND GND mn15  l=0.13u w=0.46u m=1
M10 GND N_5 N_9 GND mn15  l=0.13u w=0.34u m=1
M11 N_14 N_9 N_13 GND mn15  l=0.13u w=0.23u m=1
M12 N_13 N_9 N_14 GND mn15  l=0.13u w=0.23u m=1
M13 N_82 N_5 N_13 GND mn15  l=0.13u w=0.43u m=1
M14 N_13 N_5 N_81 GND mn15  l=0.13u w=0.23u m=1
M15 N_81 N_14 GND GND mn15  l=0.13u w=0.23u m=1
M16 N_82 N_14 GND GND mn15  l=0.13u w=0.43u m=1
M17 N_14 C GND GND mn15  l=0.13u w=0.46u m=1
M18 N_3 B VDD VDD mp15  l=0.13u w=0.4u m=1
M19 N_19 N_3 VDD VDD mp15  l=0.13u w=0.58u m=1
M20 N_5 N_7 N_3 VDD mp15  l=0.13u w=0.33u m=1
M21 N_19 A N_5 VDD mp15  l=0.13u w=0.58u m=1
M22 N_7 A VDD VDD mp15  l=0.13u w=0.4u m=1
M23 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M24 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M25 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M26 Y N_13 VDD VDD mp15  l=0.13u w=0.69u m=1
M27 N_9 N_5 VDD VDD mp15  l=0.13u w=0.52u m=1
M28 N_14 N_5 N_13 VDD mp15  l=0.13u w=0.46u m=1
M29 VDD N_14 N_20 VDD mp15  l=0.13u w=0.31u m=1
M30 N_21 N_14 VDD VDD mp15  l=0.13u w=0.62u m=1
M31 N_14 C VDD VDD mp15  l=0.13u w=0.66u m=1
M32 N_21 N_9 N_13 VDD mp15  l=0.13u w=0.62u m=1
M33 N_13 N_9 N_20 VDD mp15  l=0.13u w=0.31u m=1
.ends xr03d4
* SPICE INPUT		Tue Jul 31 20:40:54 2018	xr03dm
* EV_NETLIST Version AMD.64 Release B-2008.09.SP5.HF4.26013 2015/05/03
*
*The following line needed for Star-CR:
*CRU_OPT (KEEP_ELEMENTS "^[CR]D")
*
*The following line needed for CDL:
*.BIPOLAR

* Hierarchy Level 0

* Top of hierarchy  cell=xr03dm
.subckt xr03dm GND Y VDD B A C
M1 N_3 A GND GND mn15  l=0.13u w=0.28u m=1
M2 N_5 B GND GND mn15  l=0.13u w=0.28u m=1
M3 N_15 N_5 GND GND mn15  l=0.13u w=0.28u m=1
M4 N_15 N_3 N_6 GND mn15  l=0.13u w=0.28u m=1
M5 N_5 A N_6 GND mn15  l=0.13u w=0.3u m=1
M6 GND C N_9 GND mn15  l=0.13u w=0.28u m=1
M7 N_16 N_9 GND GND mn15  l=0.13u w=0.28u m=1
M8 N_9 N_14 N_8 GND mn15  l=0.13u w=0.28u m=1
M9 N_16 N_6 N_8 GND mn15  l=0.13u w=0.28u m=1
M10 N_14 N_6 GND GND mn15  l=0.13u w=0.28u m=1
M11 Y N_8 GND GND mn15  l=0.13u w=0.36u m=1
M12 N_5 B VDD VDD mp15  l=0.13u w=0.4u m=1
M13 N_58 N_5 VDD VDD mp15  l=0.13u w=0.4u m=1
M14 N_6 N_3 N_5 VDD mp15  l=0.13u w=0.3u m=1
M15 N_58 A N_6 VDD mp15  l=0.13u w=0.4u m=1
M16 VDD C N_9 VDD mp15  l=0.13u w=0.4u m=1
M17 N_59 N_9 VDD VDD mp15  l=0.13u w=0.4u m=1
M18 N_59 N_14 N_8 VDD mp15  l=0.13u w=0.4u m=1
M19 N_9 N_6 N_8 VDD mp15  l=0.13u w=0.28u m=1
M20 N_3 A VDD VDD mp15  l=0.13u w=0.4u m=1
M21 N_14 N_6 VDD VDD mp15  l=0.13u w=0.4u m=1
M22 Y N_8 VDD VDD mp15  l=0.13u w=0.55u m=1
.ends xr03dm
